* File: sky130_fd_sc_hvl__xnor2_1.pex.spice
* Created: Wed Sep  2 09:10:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__XNOR2_1%VNB 5 7 11 25
r33 7 25 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=0.057
+ $X2=2.64 $Y2=0.058
r34 7 11 0.00134943 $w=5.28e-06 $l=5.7e-08 $layer=MET1_cond $X=2.64 $Y=0.057
+ $X2=2.64 $Y2=0
r35 5 11 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r36 5 11 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__XNOR2_1%VPB 4 6 14 21
r42 10 21 0.00134943 $w=5.28e-06 $l=5.7e-08 $layer=MET1_cond $X=2.64 $Y=4.07
+ $X2=2.64 $Y2=4.013
r43 10 14 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=4.07
+ $X2=5.04 $Y2=4.07
r44 9 14 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=5.04
+ $Y2=4.07
r45 9 10 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r46 6 21 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=4.012
+ $X2=2.64 $Y2=4.013
r47 4 14 33.0909 $w=1.7e-07 $l=5.08232e-06 $layer=licon1_NTAP_notbjt $count=5
+ $X=0 $Y=3.985 $X2=5.04 $Y2=4.07
r48 4 9 33.0909 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=5
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__XNOR2_1%B 3 7 9 12 13 17 18 19 20 26 32
c68 12 0 1.35104e-19 $X=0.74 $Y=1.89
r69 29 32 115.031 $w=5e-07 $l=1.075e-06 $layer=POLY_cond $X=3.155 $Y=1.89
+ $X2=3.155 $Y2=2.965
r70 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.89 $X2=3.09 $Y2=1.89
r71 26 29 104.866 $w=5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.155 $Y=0.91
+ $X2=3.155 $Y2=1.89
r72 20 30 1.71028 $w=2.14e-07 $l=3e-08 $layer=LI1_cond $X=3.12 $Y=1.962 $X2=3.09
+ $Y2=1.962
r73 19 30 25.6542 $w=2.14e-07 $l=4.5e-07 $layer=LI1_cond $X=2.64 $Y=1.962
+ $X2=3.09 $Y2=1.962
r74 18 19 27.3645 $w=2.14e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.962
+ $X2=2.64 $Y2=1.962
r75 17 18 27.3645 $w=2.14e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.962
+ $X2=2.16 $Y2=1.962
r76 13 36 19.4394 $w=5.55e-07 $l=1.95e-07 $layer=POLY_cond $X=0.832 $Y=1.89
+ $X2=0.832 $Y2=2.085
r77 13 35 46.4319 $w=5.55e-07 $l=4.75e-07 $layer=POLY_cond $X=0.832 $Y=1.89
+ $X2=0.832 $Y2=1.415
r78 12 15 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.74 $Y=1.89
+ $X2=0.74 $Y2=2.015
r79 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.74
+ $Y=1.89 $X2=0.74 $Y2=1.89
r80 10 15 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=2.015
+ $X2=0.74 $Y2=2.015
r81 9 17 7.10644 $w=2.14e-07 $l=1.38996e-07 $layer=LI1_cond $X=1.565 $Y=2.015
+ $X2=1.68 $Y2=1.962
r82 9 10 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.565 $Y=2.015
+ $X2=0.905 $Y2=2.015
r83 7 36 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.86 $Y=2.965 $X2=0.86
+ $Y2=2.085
r84 3 35 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.86 $Y=0.91 $X2=0.86
+ $Y2=1.415
.ends

.subckt PM_SKY130_FD_SC_HVL__XNOR2_1%A 3 7 11 15 17 18 26 28
c47 7 0 1.35104e-19 $X=1.64 $Y=2.965
c48 3 0 1.58691e-19 $X=1.57 $Y=0.91
r49 27 28 8.56047 $w=5e-07 $l=8e-08 $layer=POLY_cond $X=2.365 $Y=1.665 $X2=2.445
+ $Y2=1.665
r50 25 27 50.2928 $w=5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.895 $Y=1.665
+ $X2=2.365 $Y2=1.665
r51 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.895
+ $Y=1.665 $X2=1.895 $Y2=1.665
r52 23 25 27.2865 $w=5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.64 $Y=1.665
+ $X2=1.895 $Y2=1.665
r53 21 23 7.49041 $w=5e-07 $l=7e-08 $layer=POLY_cond $X=1.57 $Y=1.665 $X2=1.64
+ $Y2=1.665
r54 18 26 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.895 $Y2=1.665
r55 17 18 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.665
+ $X2=1.68 $Y2=1.665
r56 13 28 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.445 $Y=1.915
+ $X2=2.445 $Y2=1.665
r57 13 15 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.445 $Y=1.915
+ $X2=2.445 $Y2=2.965
r58 9 27 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.365 $Y=1.415
+ $X2=2.365 $Y2=1.665
r59 9 11 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.365 $Y=1.415
+ $X2=2.365 $Y2=0.91
r60 5 23 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.64 $Y=1.915 $X2=1.64
+ $Y2=1.665
r61 5 7 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=1.64 $Y=1.915 $X2=1.64
+ $Y2=2.965
r62 1 21 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.57 $Y=1.415 $X2=1.57
+ $Y2=1.665
r63 1 3 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.57 $Y=1.415 $X2=1.57
+ $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HVL__XNOR2_1%A_30_107# 1 2 9 11 13 16 19 20 21 22 24 26
+ 28 30 33 37 46
c88 33 0 1.58691e-19 $X=2.325 $Y=1.315
r89 45 46 2.05781 $w=6.5e-07 $l=2.5e-08 $layer=POLY_cond $X=4.5 $Y=1.76
+ $X2=4.525 $Y2=1.76
r90 41 45 56.3839 $w=6.5e-07 $l=6.85e-07 $layer=POLY_cond $X=3.815 $Y=1.76
+ $X2=4.5 $Y2=1.76
r91 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.815
+ $Y=1.62 $X2=3.815 $Y2=1.62
r92 37 40 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.815 $Y=1.54 $X2=3.815
+ $Y2=1.62
r93 33 35 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.325 $Y=1.315
+ $X2=2.325 $Y2=1.54
r94 29 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=1.54
+ $X2=2.325 $Y2=1.54
r95 28 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.65 $Y=1.54
+ $X2=3.815 $Y2=1.54
r96 28 29 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.65 $Y=1.54
+ $X2=2.41 $Y2=1.54
r97 24 32 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=2.45 $X2=1.25
+ $Y2=2.365
r98 24 26 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=1.25 $Y=2.45
+ $X2=1.25 $Y2=3.59
r99 23 30 3.3199 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.44 $Y=1.315
+ $X2=0.275 $Y2=1.315
r100 22 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=1.315
+ $X2=2.325 $Y2=1.315
r101 22 23 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=2.24 $Y=1.315
+ $X2=0.44 $Y2=1.315
r102 20 32 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=2.365
+ $X2=1.25 $Y2=2.365
r103 20 21 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.165 $Y=2.365
+ $X2=0.36 $Y2=2.365
r104 19 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.235 $Y=2.28
+ $X2=0.36 $Y2=2.365
r105 18 30 3.24686 $w=2.9e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.235 $Y=1.4
+ $X2=0.275 $Y2=1.315
r106 18 19 40.566 $w=2.48e-07 $l=8.8e-07 $layer=LI1_cond $X=0.235 $Y=1.4
+ $X2=0.235 $Y2=2.28
r107 14 30 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.275 $Y=1.23
+ $X2=0.275 $Y2=1.315
r108 14 16 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=0.275 $Y=1.23
+ $X2=0.275 $Y2=0.68
r109 11 46 8.99251 $w=5e-07 $l=3.25e-07 $layer=POLY_cond $X=4.525 $Y=1.435
+ $X2=4.525 $Y2=1.76
r110 11 13 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.525 $Y=1.435
+ $X2=4.525 $Y2=0.95
r111 7 45 8.99251 $w=5e-07 $l=3.25e-07 $layer=POLY_cond $X=4.5 $Y=2.085 $X2=4.5
+ $Y2=1.76
r112 7 9 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=4.5 $Y=2.085 $X2=4.5
+ $Y2=2.965
r113 2 32 300 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=2.215 $X2=1.25 $Y2=2.445
r114 2 26 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=2.215 $X2=1.25 $Y2=3.59
r115 1 16 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.535 $X2=0.275 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__XNOR2_1%VPWR 1 2 3 10 13 30 34 39
r44 37 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.94 $Y=3.59
+ $X2=4.94 $Y2=3.59
r45 34 37 25.3406 $w=5.88e-07 $l=1.25e-06 $layer=LI1_cond $X=4.76 $Y=2.34
+ $X2=4.76 $Y2=3.59
r46 31 39 0.453008 $w=3.7e-07 $l=1.18e-06 $layer=MET1_cond $X=3.76 $Y=3.63
+ $X2=4.94 $Y2=3.63
r47 30 31 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.76 $Y=3.59
+ $X2=3.76 $Y2=3.59
r48 27 30 14.5058 $w=1.453e-06 $l=1.73e-06 $layer=LI1_cond $X=2.03 $Y=3.027
+ $X2=3.76 $Y2=3.027
r49 23 27 3.6055 $w=1.453e-06 $l=4.3e-07 $layer=LI1_cond $X=1.6 $Y=3.027
+ $X2=2.03 $Y2=3.027
r50 23 24 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.6 $Y=3.59
+ $X2=1.6 $Y2=3.59
r51 20 24 0.268734 $w=3.7e-07 $l=7e-07 $layer=MET1_cond $X=0.9 $Y=3.63 $X2=1.6
+ $Y2=3.63
r52 17 20 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.18 $Y=3.63
+ $X2=0.9 $Y2=3.63
r53 16 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.9 $Y=3.59 $X2=0.9
+ $Y2=3.59
r54 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.18 $Y=3.59
+ $X2=0.18 $Y2=3.59
r55 13 16 11.9274 $w=8.93e-07 $l=8.75e-07 $layer=LI1_cond $X=0.537 $Y=2.715
+ $X2=0.537 $Y2=3.59
r56 10 31 0.429974 $w=3.7e-07 $l=1.12e-06 $layer=MET1_cond $X=2.64 $Y=3.63
+ $X2=3.76 $Y2=3.63
r57 10 24 0.399262 $w=3.7e-07 $l=1.04e-06 $layer=MET1_cond $X=2.64 $Y=3.63
+ $X2=1.6 $Y2=3.63
r58 3 37 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=4.75
+ $Y=2.215 $X2=4.89 $Y2=3.59
r59 3 34 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.75
+ $Y=2.215 $X2=4.89 $Y2=2.34
r60 2 27 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.89
+ $Y=2.215 $X2=2.03 $Y2=3.59
r61 2 27 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=1.89
+ $Y=2.215 $X2=2.03 $Y2=2.385
r62 1 16 400 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=2.215 $X2=0.47 $Y2=3.59
r63 1 13 400 $w=1.7e-07 $l=5.67891e-07 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=2.215 $X2=0.47 $Y2=2.715
.ends

.subckt PM_SKY130_FD_SC_HVL__XNOR2_1%Y 1 2 9 13 14 15 21
r25 19 28 0.594378 $w=4.05e-07 $l=2.65e-07 $layer=LI1_cond $X=4.952 $Y=1.545
+ $X2=4.952 $Y2=1.81
r26 15 28 2.71111 $w=3.96e-07 $l=8.8e-08 $layer=LI1_cond $X=5.04 $Y=1.81
+ $X2=4.952 $Y2=1.81
r27 14 19 7.11385 $w=4.03e-07 $l=2.5e-07 $layer=LI1_cond $X=4.952 $Y=1.295
+ $X2=4.952 $Y2=1.545
r28 14 21 16.931 $w=4.03e-07 $l=5.95e-07 $layer=LI1_cond $X=4.952 $Y=1.295
+ $X2=4.952 $Y2=0.7
r29 13 28 12.0768 $w=3.96e-07 $l=3.92e-07 $layer=LI1_cond $X=4.56 $Y=1.81
+ $X2=4.952 $Y2=1.81
r30 9 11 57.6222 $w=2.48e-07 $l=1.25e-06 $layer=LI1_cond $X=4.15 $Y=2.34
+ $X2=4.15 $Y2=3.59
r31 7 13 12.6313 $w=3.96e-07 $l=5.2607e-07 $layer=LI1_cond $X=4.15 $Y=2.075
+ $X2=4.56 $Y2=1.81
r32 7 9 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=4.15 $Y=2.075
+ $X2=4.15 $Y2=2.34
r33 2 11 300 $w=1.7e-07 $l=1.69115e-06 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=2.215 $X2=4.11 $Y2=3.59
r34 2 9 300 $w=1.7e-07 $l=7.64951e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=2.215 $X2=4.11 $Y2=2.34
r35 1 21 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.775
+ $Y=0.575 $X2=4.915 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__XNOR2_1%VGND 1 2 7 16 20 21
r35 20 24 5.19053 $w=5.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.365 $Y=0.48
+ $X2=3.365 $Y2=0.71
r36 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.545 $Y=0.48
+ $X2=3.545 $Y2=0.48
r37 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.325 $Y=0.48
+ $X2=2.325 $Y2=0.48
r38 14 16 6.37326 $w=6.83e-07 $l=3.65e-07 $layer=LI1_cond $X=1.96 $Y=0.707
+ $X2=2.325 $Y2=0.707
r39 11 17 0.552824 $w=3.7e-07 $l=1.44e-06 $layer=MET1_cond $X=0.885 $Y=0.44
+ $X2=2.325 $Y2=0.44
r40 10 14 18.7706 $w=6.83e-07 $l=1.075e-06 $layer=LI1_cond $X=0.885 $Y=0.707
+ $X2=1.96 $Y2=0.707
r41 10 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.885 $Y=0.48
+ $X2=0.885 $Y2=0.48
r42 7 21 0.347434 $w=3.7e-07 $l=9.05e-07 $layer=MET1_cond $X=2.64 $Y=0.44
+ $X2=3.545 $Y2=0.44
r43 7 17 0.12093 $w=3.7e-07 $l=3.15e-07 $layer=MET1_cond $X=2.64 $Y=0.44
+ $X2=2.325 $Y2=0.44
r44 2 24 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=3.405
+ $Y=0.535 $X2=3.545 $Y2=0.71
r45 1 14 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.535 $X2=1.96 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HVL__XNOR2_1%A_523_107# 1 2 9 11 12 15
r31 13 15 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=4.135 $Y=1.105
+ $X2=4.135 $Y2=0.7
r32 11 13 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.97 $Y=1.195
+ $X2=4.135 $Y2=1.105
r33 11 12 64.697 $w=1.78e-07 $l=1.05e-06 $layer=LI1_cond $X=3.97 $Y=1.195
+ $X2=2.92 $Y2=1.195
r34 7 12 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.755 $Y=1.105
+ $X2=2.92 $Y2=1.195
r35 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.755 $Y=1.105
+ $X2=2.755 $Y2=0.66
r36 2 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=3.99
+ $Y=0.575 $X2=4.135 $Y2=0.7
r37 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.615
+ $Y=0.535 $X2=2.755 $Y2=0.66
.ends

