# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__o22a_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__o22a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 1.775000 2.150000 2.055000 ;
        RECT 1.980000 1.400000 2.775000 1.570000 ;
        RECT 1.980000 1.570000 2.150000 1.775000 ;
        RECT 2.605000 1.230000 4.880000 1.400000 ;
        RECT 3.035000 1.210000 3.710000 1.230000 ;
        RECT 4.550000 1.400000 4.880000 2.015000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.580000 4.195000 1.910000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.330000 1.750000 2.755000 2.120000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.955000 1.580000 3.250000 2.120000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.495000 0.380000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 5.280000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 5.280000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 5.280000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 5.280000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.985000 5.280000 4.155000 ;
      RECT 0.560000  0.365000 1.450000 1.245000 ;
      RECT 0.560000  2.650000 3.250000 3.755000 ;
      RECT 0.585000  1.425000 1.800000 1.595000 ;
      RECT 0.585000  1.595000 0.915000 2.300000 ;
      RECT 0.585000  2.300000 3.680000 2.470000 ;
      RECT 1.630000  1.050000 2.425000 1.220000 ;
      RECT 1.630000  1.220000 1.800000 1.425000 ;
      RECT 1.745000  0.265000 3.680000 0.435000 ;
      RECT 1.745000  0.435000 2.075000 0.870000 ;
      RECT 2.255000  0.880000 2.855000 1.050000 ;
      RECT 2.525000  0.615000 2.855000 0.880000 ;
      RECT 3.350000  0.435000 3.680000 1.030000 ;
      RECT 3.430000  2.175000 3.680000 2.300000 ;
      RECT 3.430000  2.470000 3.680000 3.755000 ;
      RECT 3.860000  2.195000 5.170000 3.735000 ;
      RECT 3.890000  0.365000 5.190000 1.050000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.560000  0.395000 0.730000 0.565000 ;
      RECT 0.560000  3.505000 0.730000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.920000  0.395000 1.090000 0.565000 ;
      RECT 0.920000  3.505000 1.090000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.280000  0.395000 1.450000 0.565000 ;
      RECT 1.280000  3.505000 1.450000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.640000  3.505000 1.810000 3.675000 ;
      RECT 2.000000  3.505000 2.170000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.360000  3.505000 2.530000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.720000  3.505000 2.890000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.080000  3.505000 3.250000 3.675000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.890000  3.505000 4.060000 3.675000 ;
      RECT 3.915000  0.395000 4.085000 0.565000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.250000  3.505000 4.420000 3.675000 ;
      RECT 4.275000  0.395000 4.445000 0.565000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.610000  3.505000 4.780000 3.675000 ;
      RECT 4.635000  0.395000 4.805000 0.565000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 4.970000  3.505000 5.140000 3.675000 ;
      RECT 4.995000  0.395000 5.165000 0.565000 ;
  END
END sky130_fd_sc_hvl__o22a_1
