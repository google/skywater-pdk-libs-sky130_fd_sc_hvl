* File: sky130_fd_sc_hvl__lsbuflv2hv_1.pex.spice
* Created: Wed Sep  2 09:07:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%VNB 9 11 12 23 35 42 49
r90 29 49 2.92572 $w=2.3e-07 $l=4.56e-06 $layer=MET1_cond $X=0.24 $Y=8.14
+ $X2=4.8 $Y2=8.14
r91 17 42 2.92572 $w=2.3e-07 $l=4.56e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.8
+ $Y2=0
r92 12 35 3.23369 $w=2.3e-07 $l=5.04e-06 $layer=MET1_cond $X=5.28 $Y=8.14
+ $X2=10.32 $Y2=8.14
r93 12 49 0.30797 $w=2.3e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=8.14 $X2=4.8
+ $Y2=8.14
r94 11 23 3.23369 $w=2.3e-07 $l=5.04e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=10.32
+ $Y2=0
r95 11 42 0.30797 $w=2.3e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=0 $X2=4.8
+ $Y2=0
r96 9 35 0.845455 $w=1.7e-07 $l=1.87e-06 $layer=mcon $count=11 $X=10.32 $Y=8.14
+ $X2=10.32 $Y2=8.14
r97 9 29 0.845455 $w=1.7e-07 $l=1.87e-06 $layer=mcon $count=11 $X=0.24 $Y=8.14
+ $X2=0.24 $Y2=8.14
r98 9 23 0.845455 $w=1.7e-07 $l=1.87e-06 $layer=mcon $count=11 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r99 9 17 0.845455 $w=1.7e-07 $l=1.87e-06 $layer=mcon $count=11 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%VPB 7 8 11 14 25 26 32
c69 26 0 1.93214e-19 $X=10.32 $Y=4.07
r70 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=4.07
+ $X2=10.32 $Y2=4.07
r71 21 26 1.53985 $w=2.3e-07 $l=2.4e-06 $layer=MET1_cond $X=7.92 $Y=4.07
+ $X2=10.32 $Y2=4.07
r72 20 25 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=7.92 $Y=4.07
+ $X2=10.32 $Y2=4.07
r73 20 21 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=4.07
+ $X2=7.92 $Y2=4.07
r74 15 32 2.92572 $w=2.3e-07 $l=4.56e-06 $layer=MET1_cond $X=0.24 $Y=4.07
+ $X2=4.8 $Y2=4.07
r75 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r76 11 21 1.69384 $w=2.3e-07 $l=2.64e-06 $layer=MET1_cond $X=5.28 $Y=4.07
+ $X2=7.92 $Y2=4.07
r77 11 32 0.30797 $w=2.3e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=4.07 $X2=4.8
+ $Y2=4.07
r78 8 25 60.6667 $w=1.7e-07 $l=2.64716e-06 $layer=licon1_NTAP_notbjt $count=3
+ $X=7.715 $Y=3.985 $X2=10.32 $Y2=4.07
r79 8 20 60.6667 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=3
+ $X=7.715 $Y=3.985 $X2=7.92 $Y2=4.07
r80 7 14 182 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=1 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%LVPWR 1 7 11 13 19 27
c55 13 0 1.70062e-19 $X=0.07 $Y=3.02
r56 20 27 0.433611 $w=2.85e-07 $l=8.7e-07 $layer=MET1_cond $X=3.93 $Y=3.162
+ $X2=4.8 $Y2=3.162
r57 19 22 4.74802 $w=7.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.73 $Y=3.19
+ $X2=3.73 $Y2=3.485
r58 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.93 $Y=3.19
+ $X2=3.93 $Y2=3.19
r59 17 20 0.179425 $w=2.85e-07 $l=3.6e-07 $layer=MET1_cond $X=3.57 $Y=3.162
+ $X2=3.93 $Y2=3.162
r60 16 19 0.885224 $w=7.58e-07 $l=5.5e-08 $layer=LI1_cond $X=3.73 $Y=3.135
+ $X2=3.73 $Y2=3.19
r61 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.57 $Y=3.135
+ $X2=3.57 $Y2=3.135
r62 13 27 0.239234 $w=2.85e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=3.162
+ $X2=4.8 $Y2=3.162
r63 9 16 6.31558 $w=7.58e-07 $l=1.87617e-07 $layer=LI1_cond $X=3.57 $Y=3.075
+ $X2=3.73 $Y2=3.135
r64 9 11 31.7989 $w=2.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.57 $Y=3.075
+ $X2=3.57 $Y2=2.33
r65 7 22 45.5 $w=1.7e-07 $l=7.69756e-07 $layer=licon1_NTAP_notbjt $count=4
+ $X=3.265 $Y=3.305 $X2=3.95 $Y2=3.485
r66 1 11 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=3.43
+ $Y=2.195 $X2=3.57 $Y2=2.33
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A 1 3 5 8 10 11 12 16
r32 16 19 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.66 $Y=1.695
+ $X2=2.66 $Y2=1.87
r33 11 12 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.65 $Y=1.665
+ $X2=2.65 $Y2=2.035
r34 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.66
+ $Y=1.695 $X2=2.66 $Y2=1.695
r35 6 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=2.035
+ $X2=3.355 $Y2=1.87
r36 6 8 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.355 $Y=2.035
+ $X2=3.355 $Y2=2.615
r37 3 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.705
+ $X2=3.355 $Y2=1.87
r38 3 5 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.355 $Y=1.705
+ $X2=3.355 $Y2=1.175
r39 2 19 2.83073 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.825 $Y=1.87
+ $X2=2.66 $Y2=1.87
r40 1 10 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.28 $Y=1.87
+ $X2=3.355 $Y2=1.87
r41 1 2 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=3.28 $Y=1.87
+ $X2=2.825 $Y2=1.87
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_404_1133# 1 2 7 9 10 12 13 15 16 18
+ 21 23 25 26 28 39 42 43 50 55 58 59 62 63
c103 43 0 1.93214e-19 $X=3.03 $Y=4.65
c104 26 0 1.48222e-19 $X=5.39 $Y=5.995
r105 61 62 8.79496 $w=3.78e-07 $l=2.9e-07 $layer=LI1_cond $X=3.075 $Y=2.765
+ $X2=3.075 $Y2=3.055
r106 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.145
+ $Y=1.87 $X2=4.145 $Y2=1.87
r107 56 63 1.88208 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=3.265 $Y=1.87
+ $X2=3.12 $Y2=1.87
r108 56 58 40.566 $w=2.48e-07 $l=8.8e-07 $layer=LI1_cond $X=3.265 $Y=1.87
+ $X2=4.145 $Y2=1.87
r109 55 61 17.2866 $w=2.88e-07 $l=4.35e-07 $layer=LI1_cond $X=3.12 $Y=2.33
+ $X2=3.12 $Y2=2.765
r110 52 63 4.55795 $w=2.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.12 $Y=1.995
+ $X2=3.12 $Y2=1.87
r111 52 55 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=3.12 $Y=1.995
+ $X2=3.12 $Y2=2.33
r112 48 63 4.55795 $w=2.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.12 $Y=1.745
+ $X2=3.12 $Y2=1.87
r113 48 50 33.5798 $w=2.88e-07 $l=8.45e-07 $layer=LI1_cond $X=3.12 $Y=1.745
+ $X2=3.12 $Y2=0.9
r114 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.03
+ $Y=5.33 $X2=3.03 $Y2=5.33
r115 43 46 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=3.03 $Y=4.65
+ $X2=3.03 $Y2=5.33
r116 42 45 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=3.03 $Y=4.65
+ $X2=3.03 $Y2=5.33
r117 42 62 63.3844 $w=2.88e-07 $l=1.595e-06 $layer=LI1_cond $X=3.03 $Y=4.65
+ $X2=3.03 $Y2=3.055
r118 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.03
+ $Y=4.65 $X2=3.03 $Y2=4.65
r119 38 59 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=3.86 $Y=1.87
+ $X2=4.145 $Y2=1.87
r120 38 39 5.03009 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.86 $Y=1.87
+ $X2=3.75 $Y2=1.87
r121 32 46 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=3.03 $Y=5.665
+ $X2=3.03 $Y2=5.33
r122 31 32 2.83073 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.03 $Y=5.83
+ $X2=3.03 $Y2=5.665
r123 26 28 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.39 $Y=5.995 $X2=5.39
+ $Y2=6.855
r124 23 26 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=4.61 $Y=5.83
+ $X2=5.39 $Y2=5.83
r125 23 25 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.61 $Y=5.995 $X2=4.61
+ $Y2=6.855
r126 19 39 37.0704 $w=1.5e-07 $l=1.81659e-07 $layer=POLY_cond $X=3.785 $Y=2.035
+ $X2=3.75 $Y2=1.87
r127 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.785 $Y=2.035
+ $X2=3.785 $Y2=2.615
r128 16 39 37.0704 $w=1.5e-07 $l=1.81659e-07 $layer=POLY_cond $X=3.785 $Y=1.705
+ $X2=3.75 $Y2=1.87
r129 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.785 $Y=1.705
+ $X2=3.785 $Y2=1.175
r130 13 23 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=3.83 $Y=5.83
+ $X2=4.61 $Y2=5.83
r131 13 15 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.83 $Y=5.995 $X2=3.83
+ $Y2=6.855
r132 10 13 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=3.05 $Y=5.83
+ $X2=3.83 $Y2=5.83
r133 10 31 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.05 $Y=5.83 $X2=3.03
+ $Y2=5.83
r134 10 12 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.05 $Y=5.995 $X2=3.05
+ $Y2=6.855
r135 7 31 132.895 $w=3.3e-07 $l=7.6e-07 $layer=POLY_cond $X=2.27 $Y=5.83
+ $X2=3.03 $Y2=5.83
r136 7 9 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.27 $Y=5.995 $X2=2.27
+ $Y2=6.855
r137 2 55 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=2.195 $X2=3.14 $Y2=2.33
r138 1 50 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=2.985
+ $Y=0.755 $X2=3.14 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_1197_107# 1 2 3 4 15 19 20 21 26 28
+ 31 35 36 39 48 50 54
r76 48 54 29.1379 $w=8.85e-07 $l=5.35e-07 $layer=POLY_cond $X=7.53 $Y=3.56
+ $X2=7.53 $Y2=3.025
r77 48 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.67
+ $Y=3.56 $X2=7.67 $Y2=3.56
r78 47 50 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=7.33 $Y=3.6 $X2=7.67
+ $Y2=3.6
r79 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.33
+ $Y=3.56 $X2=7.33 $Y2=3.56
r80 43 44 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=7.33 $Y=2.31
+ $X2=7.685 $Y2=2.31
r81 39 42 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=9.245 $Y=0.68
+ $X2=9.245 $Y2=1.89
r82 37 42 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=9.245 $Y=2.145
+ $X2=9.245 $Y2=1.89
r83 36 44 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.85 $Y=2.31
+ $X2=7.685 $Y2=2.31
r84 35 37 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=9.08 $Y=2.31
+ $X2=9.245 $Y2=2.145
r85 35 36 42.9547 $w=3.28e-07 $l=1.23e-06 $layer=LI1_cond $X=9.08 $Y=2.31
+ $X2=7.85 $Y2=2.31
r86 31 34 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=7.685 $Y=0.68
+ $X2=7.685 $Y2=1.89
r87 29 44 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.685 $Y=2.145
+ $X2=7.685 $Y2=2.31
r88 29 34 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.685 $Y=2.145
+ $X2=7.685 $Y2=1.89
r89 27 47 2.01087 $w=3.3e-07 $l=2.05e-07 $layer=LI1_cond $X=7.33 $Y=3.805
+ $X2=7.33 $Y2=3.6
r90 27 28 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=7.33 $Y=3.805
+ $X2=7.33 $Y2=4.47
r91 26 47 2.01087 $w=3.3e-07 $l=2.05e-07 $layer=LI1_cond $X=7.33 $Y=3.395
+ $X2=7.33 $Y2=3.6
r92 25 43 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.33 $Y=2.475
+ $X2=7.33 $Y2=2.31
r93 25 26 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=7.33 $Y=2.475
+ $X2=7.33 $Y2=3.395
r94 21 28 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=7.165 $Y=4.635
+ $X2=7.33 $Y2=4.47
r95 21 23 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=7.165 $Y=4.635
+ $X2=6.85 $Y2=4.635
r96 19 43 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.165 $Y=2.31
+ $X2=7.33 $Y2=2.31
r97 19 20 30.5572 $w=3.28e-07 $l=8.75e-07 $layer=LI1_cond $X=7.165 $Y=2.31
+ $X2=6.29 $Y2=2.31
r98 15 18 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=6.125 $Y=0.68
+ $X2=6.125 $Y2=1.89
r99 13 20 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=6.125 $Y=2.145
+ $X2=6.29 $Y2=2.31
r100 13 18 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.125 $Y=2.145
+ $X2=6.125 $Y2=1.89
r101 4 23 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=6.665
+ $Y=4.425 $X2=6.85 $Y2=4.635
r102 3 42 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=9.105
+ $Y=0.535 $X2=9.245 $Y2=1.89
r103 3 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.105
+ $Y=0.535 $X2=9.245 $Y2=0.68
r104 2 34 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=7.545
+ $Y=0.535 $X2=7.685 $Y2=1.89
r105 2 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.545
+ $Y=0.535 $X2=7.685 $Y2=0.68
r106 1 18 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=5.985
+ $Y=0.535 $X2=6.125 $Y2=1.89
r107 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.985
+ $Y=0.535 $X2=6.125 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_772_151# 1 2 7 9 10 12 13 15 16 18
+ 19 21 24 29 30 35 40 44 46
r78 44 45 23.6688 $w=3.17e-07 $l=6.15e-07 $layer=LI1_cond $X=4.03 $Y=2.31
+ $X2=4.645 $Y2=2.31
r79 43 44 1.15457 $w=3.17e-07 $l=3e-08 $layer=LI1_cond $X=4 $Y=2.31 $X2=4.03
+ $Y2=2.31
r80 38 40 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=4.03 $Y=1.41
+ $X2=4.645 $Y2=1.41
r81 36 46 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.625 $Y=2.31
+ $X2=5.485 $Y2=2.31
r82 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.625
+ $Y=2.31 $X2=5.625 $Y2=2.31
r83 33 46 94.4251 $w=3.3e-07 $l=5.4e-07 $layer=POLY_cond $X=4.945 $Y=2.31
+ $X2=5.485 $Y2=2.31
r84 32 35 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.945 $Y=2.31
+ $X2=5.625 $Y2=2.31
r85 32 33 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.945
+ $Y=2.31 $X2=4.945 $Y2=2.31
r86 30 45 6.1 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.81 $Y=2.31 $X2=4.645
+ $Y2=2.31
r87 30 32 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=4.81 $Y=2.31
+ $X2=4.945 $Y2=2.31
r88 29 45 0.469914 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=2.145
+ $X2=4.645 $Y2=2.31
r89 28 40 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=1.575
+ $X2=4.645 $Y2=1.41
r90 28 29 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=4.645 $Y=1.575
+ $X2=4.645 $Y2=2.145
r91 22 38 1.09485 $w=3.1e-07 $l=1.65e-07 $layer=LI1_cond $X=4.03 $Y=1.245
+ $X2=4.03 $Y2=1.41
r92 22 24 12.8256 $w=3.08e-07 $l=3.45e-07 $layer=LI1_cond $X=4.03 $Y=1.245
+ $X2=4.03 $Y2=0.9
r93 19 21 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.855 $Y=2.145
+ $X2=8.855 $Y2=1.285
r94 16 19 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=8.075 $Y=2.31
+ $X2=8.855 $Y2=2.31
r95 16 18 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.075 $Y=2.145
+ $X2=8.075 $Y2=1.285
r96 13 16 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=7.295 $Y=2.31
+ $X2=8.075 $Y2=2.31
r97 13 15 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.295 $Y=2.145
+ $X2=7.295 $Y2=1.285
r98 10 13 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=6.515 $Y=2.31
+ $X2=7.295 $Y2=2.31
r99 10 12 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.515 $Y=2.145
+ $X2=6.515 $Y2=1.285
r100 7 10 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=5.735 $Y=2.31
+ $X2=6.515 $Y2=2.31
r101 7 36 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=5.735 $Y=2.31
+ $X2=5.625 $Y2=2.31
r102 7 9 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.735 $Y=2.145 $X2=5.735
+ $Y2=1.285
r103 2 43 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=3.86
+ $Y=2.195 $X2=4 $Y2=2.33
r104 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.86
+ $Y=0.755 $X2=4 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_504_1221# 1 2 3 4 13 15 17 18 20 22
+ 24 30 34 35 38 42 46 51 52 53 56 60 61 65 68 73 75 76
c103 56 0 9.32604e-20 $X=6.89 $Y=2.96
c104 51 0 1.70062e-19 $X=6.35 $Y=5.665
c105 46 0 1.48222e-19 $X=5.78 $Y=6.25
r106 71 73 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.35 $Y=3.3
+ $X2=6.83 $Y2=3.3
r107 69 70 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=5.78 $Y=5.83
+ $X2=6.35 $Y2=5.83
r108 66 76 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.825 $Y=6.39
+ $X2=7.825 $Y2=6.225
r109 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.825
+ $Y=6.39 $X2=7.825 $Y2=6.39
r110 63 75 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.825 $Y=5.995
+ $X2=7.825 $Y2=5.83
r111 63 65 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=7.825 $Y=5.995
+ $X2=7.825 $Y2=6.39
r112 61 76 149.506 $w=3.3e-07 $l=8.55e-07 $layer=POLY_cond $X=7.825 $Y=5.37
+ $X2=7.825 $Y2=6.225
r113 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.825
+ $Y=5.37 $X2=7.825 $Y2=5.37
r114 58 75 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.825 $Y=5.665
+ $X2=7.825 $Y2=5.83
r115 58 60 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.825 $Y=5.665
+ $X2=7.825 $Y2=5.37
r116 54 73 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.83 $Y=3.135
+ $X2=6.83 $Y2=3.3
r117 54 56 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=6.83 $Y=3.135
+ $X2=6.83 $Y2=2.96
r118 53 70 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.515 $Y=5.83
+ $X2=6.35 $Y2=5.83
r119 52 75 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.66 $Y=5.83
+ $X2=7.825 $Y2=5.83
r120 52 53 39.9863 $w=3.28e-07 $l=1.145e-06 $layer=LI1_cond $X=7.66 $Y=5.83
+ $X2=6.515 $Y2=5.83
r121 51 70 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.35 $Y=5.665
+ $X2=6.35 $Y2=5.83
r122 50 71 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.35 $Y=3.465
+ $X2=6.35 $Y2=3.3
r123 50 51 76.8295 $w=3.28e-07 $l=2.2e-06 $layer=LI1_cond $X=6.35 $Y=3.465
+ $X2=6.35 $Y2=5.665
r124 46 48 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=5.78 $Y=6.25
+ $X2=5.78 $Y2=7.46
r125 44 69 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.78 $Y=5.995
+ $X2=5.78 $Y2=5.83
r126 44 46 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.78 $Y=5.995
+ $X2=5.78 $Y2=6.25
r127 43 68 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.385 $Y=5.83
+ $X2=4.22 $Y2=5.83
r128 42 69 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.615 $Y=5.83
+ $X2=5.78 $Y2=5.83
r129 42 43 42.9547 $w=3.28e-07 $l=1.23e-06 $layer=LI1_cond $X=5.615 $Y=5.83
+ $X2=4.385 $Y2=5.83
r130 38 40 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=4.22 $Y=6.25
+ $X2=4.22 $Y2=7.46
r131 36 68 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.22 $Y=5.995
+ $X2=4.22 $Y2=5.83
r132 36 38 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.22 $Y=5.995
+ $X2=4.22 $Y2=6.25
r133 34 68 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.055 $Y=5.83
+ $X2=4.22 $Y2=5.83
r134 34 35 42.9547 $w=3.28e-07 $l=1.23e-06 $layer=LI1_cond $X=4.055 $Y=5.83
+ $X2=2.825 $Y2=5.83
r135 30 32 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=2.66 $Y=6.25
+ $X2=2.66 $Y2=7.46
r136 28 35 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=2.66 $Y=5.995
+ $X2=2.825 $Y2=5.83
r137 28 30 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.66 $Y=5.995
+ $X2=2.66 $Y2=6.25
r138 25 61 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=7.825 $Y=4.975
+ $X2=7.825 $Y2=5.37
r139 24 25 19.6718 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.825 $Y=4.635
+ $X2=7.825 $Y2=4.975
r140 22 24 26.3581 $w=6.8e-07 $l=3.35e-07 $layer=POLY_cond $X=7.49 $Y=4.635
+ $X2=7.825 $Y2=4.635
r141 18 27 56.8991 $w=5e-07 $l=5.85e-07 $layer=POLY_cond $X=9.07 $Y=6.975
+ $X2=9.07 $Y2=6.39
r142 18 20 24.582 $w=5e-07 $l=2.55e-07 $layer=POLY_cond $X=9.07 $Y=6.975
+ $X2=9.07 $Y2=7.23
r143 15 27 56.8991 $w=5e-07 $l=5.85e-07 $layer=POLY_cond $X=9.07 $Y=5.805
+ $X2=9.07 $Y2=6.39
r144 15 17 60.732 $w=5e-07 $l=6.3e-07 $layer=POLY_cond $X=9.07 $Y=5.805 $X2=9.07
+ $Y2=5.175
r145 14 66 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.99 $Y=6.39
+ $X2=7.825 $Y2=6.39
r146 13 27 10.2987 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=8.82 $Y=6.39
+ $X2=9.07 $Y2=6.39
r147 13 14 145.135 $w=3.3e-07 $l=8.3e-07 $layer=POLY_cond $X=8.82 $Y=6.39
+ $X2=7.99 $Y2=6.39
r148 4 56 300 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=2 $X=6.665
+ $Y=2.815 $X2=6.89 $Y2=2.96
r149 3 48 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=5.64
+ $Y=6.105 $X2=5.78 $Y2=7.46
r150 3 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.64
+ $Y=6.105 $X2=5.78 $Y2=6.25
r151 2 40 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=4.08
+ $Y=6.105 $X2=4.22 $Y2=7.46
r152 2 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.08
+ $Y=6.105 $X2=4.22 $Y2=6.25
r153 1 32 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=2.52
+ $Y=6.105 $X2=2.66 $Y2=7.46
r154 1 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.52
+ $Y=6.105 $X2=2.66 $Y2=6.25
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_1711_885# 1 2 9 13 17 23 27 28 30
r48 28 33 16.3371 $w=6.95e-07 $l=1.65e-07 $layer=POLY_cond $X=9.797 $Y=6.39
+ $X2=9.797 $Y2=6.555
r49 28 32 16.3371 $w=6.95e-07 $l=1.65e-07 $layer=POLY_cond $X=9.797 $Y=6.39
+ $X2=9.797 $Y2=6.225
r50 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.955
+ $Y=6.39 $X2=9.955 $Y2=6.39
r51 25 30 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.845 $Y=6.39
+ $X2=8.68 $Y2=6.39
r52 25 27 38.764 $w=3.28e-07 $l=1.11e-06 $layer=LI1_cond $X=8.845 $Y=6.39
+ $X2=9.955 $Y2=6.39
r53 21 30 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.68 $Y=6.555
+ $X2=8.68 $Y2=6.39
r54 21 23 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.68 $Y=6.555
+ $X2=8.68 $Y2=7
r55 17 20 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=8.68 $Y=4.57
+ $X2=8.68 $Y2=5.78
r56 15 30 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.68 $Y=6.225
+ $X2=8.68 $Y2=6.39
r57 15 20 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.68 $Y=6.225
+ $X2=8.68 $Y2=5.78
r58 13 33 72.229 $w=5e-07 $l=6.75e-07 $layer=POLY_cond $X=9.895 $Y=7.23
+ $X2=9.895 $Y2=6.555
r59 9 32 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=9.895 $Y=5.175
+ $X2=9.895 $Y2=6.225
r60 2 20 300 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_PDIFF $count=2 $X=8.555
+ $Y=4.425 $X2=8.68 $Y2=5.78
r61 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=8.555
+ $Y=4.425 $X2=8.68 $Y2=4.57
r62 1 23 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=8.555
+ $Y=6.855 $X2=8.68 $Y2=7
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%VPWR 1 2 3 10 11 15 21 25 28 32 37 43
c66 25 0 9.32604e-20 $X=8.48 $Y=3.56
r67 31 34 24.327 $w=5.88e-07 $l=1.2e-06 $layer=LI1_cond $X=9.505 $Y=4.58
+ $X2=9.505 $Y2=5.78
r68 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.685 $Y=4.58
+ $X2=9.685 $Y2=4.58
r69 28 31 0.202725 $w=5.88e-07 $l=1e-08 $layer=LI1_cond $X=9.505 $Y=4.57
+ $X2=9.505 $Y2=4.58
r70 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.48 $Y=3.56
+ $X2=8.48 $Y2=3.56
r71 21 24 12.1635 $w=5.88e-07 $l=6e-07 $layer=LI1_cond $X=8.3 $Y=2.96 $X2=8.3
+ $Y2=3.56
r72 18 32 0.558582 $w=3.7e-07 $l=1.455e-06 $layer=MET1_cond $X=8.23 $Y=4.51
+ $X2=9.685 $Y2=4.51
r73 15 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.23 $Y=4.58
+ $X2=8.23 $Y2=4.58
r74 11 18 1.13252 $w=3.7e-07 $l=2.95e-06 $layer=MET1_cond $X=5.28 $Y=4.51
+ $X2=8.23 $Y2=4.51
r75 11 43 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=4.51
+ $X2=4.8 $Y2=4.51
r76 10 25 1.2285 $w=3.7e-07 $l=3.2e-06 $layer=MET1_cond $X=5.28 $Y=3.63 $X2=8.48
+ $Y2=3.63
r77 10 37 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=3.63
+ $X2=4.8 $Y2=3.63
r78 3 34 300 $w=1.7e-07 $l=1.44454e-06 $layer=licon1_PDIFF $count=2 $X=9.32
+ $Y=4.425 $X2=9.505 $Y2=5.78
r79 3 28 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=9.32
+ $Y=4.425 $X2=9.505 $Y2=4.57
r80 2 21 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.03
+ $Y=2.815 $X2=8.17 $Y2=2.96
r81 1 15 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.99
+ $Y=4.425 $X2=8.13 $Y2=4.635
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%X 1 2 7 8 9 10 11 21 31 45
r17 35 45 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=10.285 $Y=6.89
+ $X2=10.285 $Y2=6.845
r18 31 41 2.40092 $w=2.38e-07 $l=5e-08 $layer=LI1_cond $X=10.33 $Y=6.105
+ $X2=10.33 $Y2=6.055
r19 11 45 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=10.285 $Y=6.825
+ $X2=10.285 $Y2=6.845
r20 11 43 4.36998 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=10.285 $Y=6.825
+ $X2=10.285 $Y2=6.725
r21 11 38 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=10.285 $Y=6.91
+ $X2=10.285 $Y2=7
r22 11 35 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=10.285 $Y=6.91
+ $X2=10.285 $Y2=6.89
r23 10 43 12.0046 $w=2.38e-07 $l=2.5e-07 $layer=LI1_cond $X=10.33 $Y=6.475
+ $X2=10.33 $Y2=6.725
r24 9 41 1.50633 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=10.285 $Y=6.037
+ $X2=10.285 $Y2=6.055
r25 9 19 5.13361 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=10.285 $Y=6.037
+ $X2=10.285 $Y2=5.89
r26 9 10 16.9505 $w=2.38e-07 $l=3.53e-07 $layer=LI1_cond $X=10.33 $Y=6.122
+ $X2=10.33 $Y2=6.475
r27 9 31 0.816314 $w=2.38e-07 $l=1.7e-08 $layer=LI1_cond $X=10.33 $Y=6.122
+ $X2=10.33 $Y2=6.105
r28 8 19 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=10.285 $Y=5.735
+ $X2=10.285 $Y2=5.89
r29 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.285 $Y=5.365
+ $X2=10.285 $Y2=5.735
r30 7 21 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=10.285 $Y=5.365
+ $X2=10.285 $Y2=4.57
r31 2 8 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=10.145
+ $Y=4.425 $X2=10.285 $Y2=5.78
r32 2 21 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=10.145
+ $Y=4.425 $X2=10.285 $Y2=4.57
r33 1 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.145
+ $Y=6.855 $X2=10.285 $Y2=7
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%VGND 1 2 3 4 5 6 7 8 25 26 29 31 33 34
+ 35 39 43 45 46 50 57 63 72 76 84 92 100 101 108 112 115 122 132
r129 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.57 $Y=0.51
+ $X2=3.57 $Y2=0.51
r130 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.685 $Y=7.63
+ $X2=9.685 $Y2=7.63
r131 108 111 12.7717 $w=5.88e-07 $l=6.3e-07 $layer=LI1_cond $X=9.505 $Y=7
+ $X2=9.505 $Y2=7.63
r132 103 105 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=8.465 $Y=0.68
+ $X2=8.465 $Y2=1.89
r133 100 103 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=8.465 $Y=0.51
+ $X2=8.465 $Y2=0.68
r134 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.645 $Y=0.51
+ $X2=8.645 $Y2=0.51
r135 95 97 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=6.905 $Y=0.68
+ $X2=6.905 $Y2=1.89
r136 93 101 0.598892 $w=3.7e-07 $l=1.56e-06 $layer=MET1_cond $X=7.085 $Y=0.44
+ $X2=8.645 $Y2=0.44
r137 92 95 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=6.905 $Y=0.51
+ $X2=6.905 $Y2=0.68
r138 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.085 $Y=0.51
+ $X2=7.085 $Y2=0.51
r139 87 89 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=5.345 $Y=0.68
+ $X2=5.345 $Y2=1.89
r140 85 93 0.598892 $w=3.7e-07 $l=1.56e-06 $layer=MET1_cond $X=5.525 $Y=0.44
+ $X2=7.085 $Y2=0.44
r141 84 87 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=5.345 $Y=0.51
+ $X2=5.345 $Y2=0.68
r142 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.525 $Y=0.51
+ $X2=5.525 $Y2=0.51
r143 82 132 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=5.18 $Y=7.7
+ $X2=4.7 $Y2=7.7
r144 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.18 $Y=7.63
+ $X2=5.18 $Y2=7.63
r145 79 81 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=5 $Y=7.46 $X2=5
+ $Y2=7.63
r146 76 79 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=5 $Y=6.25 $X2=5
+ $Y2=7.46
r147 73 122 0.333998 $w=3.7e-07 $l=8.7e-07 $layer=MET1_cond $X=3.93 $Y=0.44
+ $X2=4.8 $Y2=0.44
r148 73 116 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=3.93 $Y=0.44
+ $X2=3.57 $Y2=0.44
r149 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.93 $Y=0.45
+ $X2=3.93 $Y2=0.45
r150 70 115 5.89082 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=3.705 $Y=0.45
+ $X2=3.57 $Y2=0.45
r151 70 72 11.2739 $w=2.28e-07 $l=2.25e-07 $layer=LI1_cond $X=3.705 $Y=0.45
+ $X2=3.93 $Y2=0.45
r152 69 132 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=3.62 $Y=7.7
+ $X2=4.7 $Y2=7.7
r153 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.62 $Y=7.63
+ $X2=3.62 $Y2=7.63
r154 66 68 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=3.44 $Y=7.46
+ $X2=3.44 $Y2=7.63
r155 63 66 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=3.44 $Y=6.25
+ $X2=3.44 $Y2=7.46
r156 60 116 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=3.21 $Y=0.44
+ $X2=3.57 $Y2=0.44
r157 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.21 $Y=0.45
+ $X2=3.21 $Y2=0.45
r158 57 115 5.89082 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=3.435 $Y=0.45
+ $X2=3.57 $Y2=0.45
r159 57 59 11.2739 $w=2.28e-07 $l=2.25e-07 $layer=LI1_cond $X=3.435 $Y=0.45
+ $X2=3.21 $Y2=0.45
r160 56 69 0.598892 $w=3.7e-07 $l=1.56e-06 $layer=MET1_cond $X=2.06 $Y=7.7
+ $X2=3.62 $Y2=7.7
r161 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.06 $Y=7.63
+ $X2=2.06 $Y2=7.63
r162 53 55 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=1.88 $Y=7.46
+ $X2=1.88 $Y2=7.63
r163 50 53 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=1.88 $Y=6.25
+ $X2=1.88 $Y2=7.46
r164 46 112 1.6911 $w=3.7e-07 $l=4.405e-06 $layer=MET1_cond $X=5.28 $Y=7.7
+ $X2=9.685 $Y2=7.7
r165 46 82 0.0383905 $w=3.7e-07 $l=1e-07 $layer=MET1_cond $X=5.28 $Y=7.7
+ $X2=5.18 $Y2=7.7
r166 45 85 0.0940568 $w=3.7e-07 $l=2.45e-07 $layer=MET1_cond $X=5.28 $Y=0.44
+ $X2=5.525 $Y2=0.44
r167 45 122 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=0.44
+ $X2=4.8 $Y2=0.44
r168 44 100 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=8.465 $Y=0.425
+ $X2=8.465 $Y2=0.51
r169 42 92 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=0.425
+ $X2=6.905 $Y2=0.51
r170 42 43 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=0.425
+ $X2=6.905 $Y2=0.34
r171 41 84 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=5.345 $Y=0.425
+ $X2=5.345 $Y2=0.51
r172 40 81 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=7.715 $X2=5
+ $Y2=7.63
r173 38 68 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=7.715
+ $X2=3.44 $Y2=7.63
r174 38 39 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=7.715
+ $X2=3.44 $Y2=7.8
r175 37 55 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=7.715
+ $X2=1.88 $Y2=7.63
r176 36 43 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=7.2 $Y=0.34
+ $X2=6.905 $Y2=0.34
r177 35 44 9.96617 $w=1.7e-07 $l=3.34813e-07 $layer=LI1_cond $X=8.17 $Y=0.34
+ $X2=8.465 $Y2=0.425
r178 35 36 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=8.17 $Y=0.34
+ $X2=7.2 $Y2=0.34
r179 34 41 9.96617 $w=1.7e-07 $l=3.34813e-07 $layer=LI1_cond $X=5.64 $Y=0.34
+ $X2=5.345 $Y2=0.425
r180 33 43 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.61 $Y=0.34
+ $X2=6.905 $Y2=0.34
r181 33 34 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=6.61 $Y=0.34
+ $X2=5.64 $Y2=0.34
r182 32 39 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.735 $Y=7.8
+ $X2=3.44 $Y2=7.8
r183 31 40 9.96617 $w=1.7e-07 $l=3.34813e-07 $layer=LI1_cond $X=4.705 $Y=7.8
+ $X2=5 $Y2=7.715
r184 31 32 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=4.705 $Y=7.8
+ $X2=3.735 $Y2=7.8
r185 27 115 0.77205 $w=2.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.57 $Y=0.565
+ $X2=3.57 $Y2=0.45
r186 27 29 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.57 $Y=0.565
+ $X2=3.57 $Y2=0.88
r187 26 37 9.96617 $w=1.7e-07 $l=3.34813e-07 $layer=LI1_cond $X=2.175 $Y=7.8
+ $X2=1.88 $Y2=7.715
r188 25 39 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.145 $Y=7.8
+ $X2=3.44 $Y2=7.8
r189 25 26 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=3.145 $Y=7.8
+ $X2=2.175 $Y2=7.8
r190 8 108 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=9.32
+ $Y=6.855 $X2=9.505 $Y2=7
r191 7 105 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=8.325
+ $Y=0.535 $X2=8.465 $Y2=1.89
r192 7 103 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.325
+ $Y=0.535 $X2=8.465 $Y2=0.68
r193 6 97 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.535 $X2=6.905 $Y2=1.89
r194 6 95 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.535 $X2=6.905 $Y2=0.68
r195 5 89 91 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.535 $X2=5.345 $Y2=1.89
r196 5 87 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.535 $X2=5.345 $Y2=0.68
r197 4 79 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=4.86
+ $Y=6.105 $X2=5 $Y2=7.46
r198 4 76 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.86
+ $Y=6.105 $X2=5 $Y2=6.25
r199 3 29 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.43
+ $Y=0.755 $X2=3.57 $Y2=0.88
r200 2 66 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=3.3
+ $Y=6.105 $X2=3.44 $Y2=7.46
r201 2 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.3
+ $Y=6.105 $X2=3.44 $Y2=6.25
r202 1 53 91 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_NDIFF $count=2 $X=1.755
+ $Y=6.105 $X2=1.88 $Y2=7.46
r203 1 50 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.755
+ $Y=6.105 $X2=1.88 $Y2=6.25
.ends

