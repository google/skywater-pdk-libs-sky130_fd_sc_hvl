* File: sky130_fd_sc_hvl__inv_2.spice
* Created: Wed Sep  2 09:06:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__inv_2.pex.spice"
.subckt sky130_fd_sc_hvl__inv_2  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_Y_M1001_d N_A_M1001_g N_VGND_M1001_s N_VNB_M1001_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.21375 PD=1.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5 SA=250000 SB=250001
+ A=0.375 P=2.5 MULT=1
MM1003 N_Y_M1001_d N_A_M1003_g N_VGND_M1003_s N_VNB_M1001_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.21375 PD=1.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5 SA=250001 SB=250000
+ A=0.375 P=2.5 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.4275 AS=0.21 PD=3.57 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250000 SB=250001
+ A=0.75 P=4 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_Y_M1000_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.4275 AS=0.21 PD=3.57 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001 SB=250000
+ A=0.75 P=4 MULT=1
DX4_noxref N_VNB_M1001_b N_VPB_M1000_b NWDIODE A=7.956 P=11.32
*
.include "sky130_fd_sc_hvl__inv_2.pxi.spice"
*
.ends
*
*
