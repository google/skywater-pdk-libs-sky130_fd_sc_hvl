* NGSPICE file created from sky130_fd_sc_hvl__xnor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__xnor2_1 A B VGND VNB VPB VPWR Y
M1000 a_539_443# A VPWR VPB phv w=1.5e+06u l=500000u
+  ad=3.15e+11p pd=3.42e+06u as=1.3125e+12p ps=1.075e+07u
M1001 Y B a_539_443# VPB phv w=1.5e+06u l=500000u
+  ad=1.2675e+12p pd=4.69e+06u as=0p ps=0u
M1002 Y a_30_107# a_523_107# VNB nhv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=4.3125e+11p ps=4.15e+06u
M1003 VPWR A a_30_107# VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=4.2e+11p ps=3.56e+06u
M1004 a_222_107# B a_30_107# VNB nhv w=750000u l=500000u
+  ad=1.575e+11p pd=1.92e+06u as=3.45e+11p ps=2.42e+06u
M1005 VGND A a_222_107# VNB nhv w=750000u l=500000u
+  ad=4.35e+11p pd=4.16e+06u as=0p ps=0u
M1006 VGND B a_523_107# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_30_107# Y VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_523_107# A VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_30_107# B VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends

