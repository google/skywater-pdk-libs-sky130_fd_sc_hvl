* File: sky130_fd_sc_hvl__or3_1.pex.spice
* Created: Wed Sep  2 09:09:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__OR3_1%VNB 5 7 11 25
r32 7 25 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=0.057
+ $X2=1.92 $Y2=0.058
r33 7 11 0.00185547 $w=3.84e-06 $l=5.7e-08 $layer=MET1_cond $X=1.92 $Y=0.057
+ $X2=1.92 $Y2=0
r34 5 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r35 5 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__OR3_1%VPB 4 6 14 21
r19 10 21 0.00185547 $w=3.84e-06 $l=5.7e-08 $layer=MET1_cond $X=1.92 $Y=4.07
+ $X2=1.92 $Y2=4.013
r20 10 14 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=4.07
+ $X2=3.6 $Y2=4.07
r21 9 14 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=3.6
+ $Y2=4.07
r22 9 10 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r23 6 21 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=4.012
+ $X2=1.92 $Y2=4.013
r24 4 14 45.5 $w=1.7e-07 $l=3.64225e-06 $layer=licon1_NTAP_notbjt $count=4 $X=0
+ $Y=3.985 $X2=3.6 $Y2=4.07
r25 4 9 45.5 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=4 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__OR3_1%C 3 7 8 9 13
c25 13 0 1.09826e-19 $X=0.665 $Y=0.745
r26 13 16 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=0.665 $Y=0.745
+ $X2=0.665 $Y2=1.28
r27 8 9 18.7737 $w=3.08e-07 $l=5.05e-07 $layer=LI1_cond $X=0.695 $Y=1.235
+ $X2=1.2 $Y2=1.235
r28 8 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.695
+ $Y=1.28 $X2=0.695 $Y2=1.28
r29 6 16 43.8724 $w=5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.665 $Y=1.69 $X2=0.665
+ $Y2=1.28
r30 6 7 50.0028 $w=5.35e-07 $l=5e-07 $layer=POLY_cond $X=0.682 $Y=1.69 $X2=0.682
+ $Y2=2.19
r31 3 7 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.7 $Y=2.53 $X2=0.7
+ $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_HVL__OR3_1%B 1 2 3 4 18 22 24
r25 21 24 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.455 $Y=1.995
+ $X2=1.455 $Y2=2.53
r26 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=1.995 $X2=1.37 $Y2=1.995
r27 18 21 133.757 $w=5e-07 $l=1.25e-06 $layer=POLY_cond $X=1.455 $Y=0.745
+ $X2=1.455 $Y2=1.995
r28 3 4 4.85376 $w=9.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.07 $Y=2.775 $X2=1.07
+ $Y2=3.145
r29 2 3 4.85376 $w=9.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.07 $Y=2.405 $X2=1.07
+ $Y2=2.775
r30 1 2 4.85376 $w=9.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.07 $Y=2.035 $X2=1.07
+ $Y2=2.405
r31 1 22 0.524731 $w=9.28e-07 $l=4e-08 $layer=LI1_cond $X=1.07 $Y=2.035 $X2=1.07
+ $Y2=1.995
.ends

.subckt PM_SKY130_FD_SC_HVL__OR3_1%A 3 7 9 12
c31 12 0 1.38666e-20 $X=2.08 $Y=1.28
r32 12 15 29.5733 $w=5.7e-07 $l=3.05e-07 $layer=POLY_cond $X=2.2 $Y=1.28 $X2=2.2
+ $Y2=1.585
r33 12 14 19.2482 $w=5.7e-07 $l=1.95e-07 $layer=POLY_cond $X=2.2 $Y=1.28 $X2=2.2
+ $Y2=1.085
r34 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.28 $X2=2.08 $Y2=1.28
r35 7 14 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.235 $Y=0.745 $X2=2.235
+ $Y2=1.085
r36 3 15 101.121 $w=5e-07 $l=9.45e-07 $layer=POLY_cond $X=2.165 $Y=2.53
+ $X2=2.165 $Y2=1.585
.ends

.subckt PM_SKY130_FD_SC_HVL__OR3_1%A_30_107# 1 2 3 12 16 20 24 26 29 30 32 36 38
+ 39 43
c69 39 0 1.38666e-20 $X=3.09 $Y=1.645
c70 36 0 1.09826e-19 $X=1.845 $Y=0.745
r71 43 47 32.4104 $w=5.2e-07 $l=3.15e-07 $layer=POLY_cond $X=3.165 $Y=1.77
+ $X2=3.165 $Y2=2.085
r72 43 46 36.5261 $w=5.2e-07 $l=3.55e-07 $layer=POLY_cond $X=3.165 $Y=1.77
+ $X2=3.165 $Y2=1.415
r73 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.77 $X2=3.09 $Y2=1.77
r74 39 42 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.09 $Y=1.645
+ $X2=3.09 $Y2=1.77
r75 33 36 5.41509 $w=4.13e-07 $l=1.95e-07 $layer=LI1_cond $X=1.65 $Y=0.702
+ $X2=1.845 $Y2=0.702
r76 31 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=1.645
+ $X2=1.65 $Y2=1.645
r77 30 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=1.645
+ $X2=3.09 $Y2=1.645
r78 30 31 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=2.925 $Y=1.645
+ $X2=1.735 $Y2=1.645
r79 29 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=1.56 $X2=1.65
+ $Y2=1.645
r80 28 33 6.00275 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=1.65 $Y=0.91
+ $X2=1.65 $Y2=0.702
r81 28 29 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.65 $Y=0.91
+ $X2=1.65 $Y2=1.56
r82 27 32 2.49072 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.395 $Y=1.645
+ $X2=0.27 $Y2=1.645
r83 26 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.565 $Y=1.645
+ $X2=1.65 $Y2=1.645
r84 26 27 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=1.565 $Y=1.645
+ $X2=0.395 $Y2=1.645
r85 22 32 3.95216 $w=2.32e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=1.73
+ $X2=0.27 $Y2=1.645
r86 22 24 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=0.27 $Y=1.73 $X2=0.27
+ $Y2=2.53
r87 18 32 3.95216 $w=2.32e-07 $l=9.35682e-08 $layer=LI1_cond $X=0.252 $Y=1.56
+ $X2=0.27 $Y2=1.645
r88 18 20 43.6856 $w=2.13e-07 $l=8.15e-07 $layer=LI1_cond $X=0.252 $Y=1.56
+ $X2=0.252 $Y2=0.745
r89 16 46 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.175 $Y=0.91
+ $X2=3.175 $Y2=1.415
r90 12 47 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.155 $Y=2.965
+ $X2=3.155 $Y2=2.085
r91 3 24 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=2.32 $X2=0.31 $Y2=2.53
r92 2 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.705
+ $Y=0.535 $X2=1.845 $Y2=0.745
r93 1 20 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.535 $X2=0.275 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__OR3_1%VPWR 1 4 11 15
r21 11 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.195 $Y=3.59
+ $X2=3.195 $Y2=3.59
r22 11 12 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.755 $Y=3.59
+ $X2=1.755 $Y2=3.59
r23 9 11 6.39887 $w=1.592e-06 $l=8.35e-07 $layer=LI1_cond $X=2.45 $Y=2.755
+ $X2=2.45 $Y2=3.59
r24 7 9 3.18028 $w=1.592e-06 $l=4.15e-07 $layer=LI1_cond $X=2.45 $Y=2.34
+ $X2=2.45 $Y2=2.755
r25 4 15 0.489479 $w=3.7e-07 $l=1.275e-06 $layer=MET1_cond $X=1.92 $Y=3.63
+ $X2=3.195 $Y2=3.63
r26 4 12 0.0633444 $w=3.7e-07 $l=1.65e-07 $layer=MET1_cond $X=1.92 $Y=3.63
+ $X2=1.755 $Y2=3.63
r27 1 11 400 $w=1.7e-07 $l=1.43436e-06 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=2.32 $X2=2.765 $Y2=3.59
r28 1 9 400 $w=1.7e-07 $l=5.84359e-07 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=2.32 $X2=2.765 $Y2=2.755
r29 1 7 600 $w=1.7e-07 $l=3.59861e-07 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=2.32 $X2=2.765 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__OR3_1%X 1 2 7 8 9 10 11 12 13 22
r14 13 40 20.1113 $w=2.53e-07 $l=4.45e-07 $layer=LI1_cond $X=3.587 $Y=3.145
+ $X2=3.587 $Y2=3.59
r15 12 13 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=2.775
+ $X2=3.587 $Y2=3.145
r16 11 12 19.6593 $w=2.53e-07 $l=4.35e-07 $layer=LI1_cond $X=3.587 $Y=2.34
+ $X2=3.587 $Y2=2.775
r17 10 11 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=3.587 $Y=2.035
+ $X2=3.587 $Y2=2.34
r18 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=1.665
+ $X2=3.587 $Y2=2.035
r19 8 9 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=1.295
+ $X2=3.587 $Y2=1.665
r20 7 8 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=0.925
+ $X2=3.587 $Y2=1.295
r21 7 22 11.0725 $w=2.53e-07 $l=2.45e-07 $layer=LI1_cond $X=3.587 $Y=0.925
+ $X2=3.587 $Y2=0.68
r22 2 40 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=2.215 $X2=3.545 $Y2=3.59
r23 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=2.215 $X2=3.545 $Y2=2.34
r24 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.425
+ $Y=0.535 $X2=3.565 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__OR3_1%VGND 1 2 7 10 17 18
r34 21 23 8.92596 $w=6.68e-07 $l=5e-07 $layer=LI1_cond $X=2.955 $Y=0.66
+ $X2=2.955 $Y2=1.16
r35 17 21 3.21335 $w=6.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.955 $Y=0.48
+ $X2=2.955 $Y2=0.66
r36 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.135 $Y=0.48
+ $X2=3.135 $Y2=0.48
r37 10 14 4.05582 $w=8.53e-07 $l=2.65e-07 $layer=LI1_cond $X=0.957 $Y=0.48
+ $X2=0.957 $Y2=0.745
r38 10 11 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.25 $Y=0.48
+ $X2=1.25 $Y2=0.48
r39 7 18 0.466445 $w=3.7e-07 $l=1.215e-06 $layer=MET1_cond $X=1.92 $Y=0.44
+ $X2=3.135 $Y2=0.44
r40 7 11 0.257217 $w=3.7e-07 $l=6.7e-07 $layer=MET1_cond $X=1.92 $Y=0.44
+ $X2=1.25 $Y2=0.44
r41 2 23 182 $w=1.7e-07 $l=7.60345e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.535 $X2=2.785 $Y2=1.16
r42 2 21 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.535 $X2=2.785 $Y2=0.66
r43 1 14 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.915
+ $Y=0.535 $X2=1.055 $Y2=0.745
.ends

