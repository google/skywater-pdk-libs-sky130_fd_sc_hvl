* File: sky130_fd_sc_hvl__nand2_1.pex.spice
* Created: Fri Aug 28 09:37:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__NAND2_1%VNB 5 7 11 25
r14 7 25 5.20833e-05 $w=2.4e-06 $l=1e-09 $layer=MET1_cond $X=1.2 $Y=0.057
+ $X2=1.2 $Y2=0.058
r15 7 11 0.00296875 $w=2.4e-06 $l=5.7e-08 $layer=MET1_cond $X=1.2 $Y=0.057
+ $X2=1.2 $Y2=0
r16 5 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r17 5 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND2_1%VPB 4 6 14 21
r20 10 21 0.00296875 $w=2.4e-06 $l=5.7e-08 $layer=MET1_cond $X=1.2 $Y=4.07
+ $X2=1.2 $Y2=4.013
r21 10 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=4.07
+ $X2=2.16 $Y2=4.07
r22 9 14 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=2.16 $Y2=4.07
r23 9 10 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r24 6 21 5.20833e-05 $w=2.4e-06 $l=1e-09 $layer=MET1_cond $X=1.2 $Y=4.012
+ $X2=1.2 $Y2=4.013
r25 4 14 72.8 $w=1.7e-07 $l=2.20209e-06 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=2.16 $Y2=4.07
r26 4 9 72.8 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND2_1%B 1 2 6 10 12
c20 6 0 1.03339e-19 $X=0.915 $Y=0.93
r21 9 12 127.872 $w=5e-07 $l=1.195e-06 $layer=POLY_cond $X=0.915 $Y=1.77
+ $X2=0.915 $Y2=2.965
r22 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.85
+ $Y=1.77 $X2=0.85 $Y2=1.77
r23 6 9 89.8849 $w=5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.915 $Y=0.93 $X2=0.915
+ $Y2=1.77
r24 2 10 3.89137 $w=3.83e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.742
+ $X2=0.85 $Y2=1.742
r25 1 2 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.742 $X2=0.72
+ $Y2=1.742
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND2_1%A 3 7 9 15
r28 13 15 34.1596 $w=6.5e-07 $l=4.15e-07 $layer=POLY_cond $X=1.695 $Y=1.76
+ $X2=2.11 $Y2=1.76
r29 11 13 5.76186 $w=6.5e-07 $l=7e-08 $layer=POLY_cond $X=1.625 $Y=1.76
+ $X2=1.695 $Y2=1.76
r30 9 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.69 $X2=2.11 $Y2=1.69
r31 5 13 8.99251 $w=5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.695 $Y=2.085
+ $X2=1.695 $Y2=1.76
r32 5 7 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.695 $Y=2.085 $X2=1.695
+ $Y2=2.965
r33 1 11 8.99251 $w=5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.625 $Y=1.435
+ $X2=1.625 $Y2=1.76
r34 1 3 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.625 $Y=1.435 $X2=1.625
+ $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND2_1%VPWR 1 2 7 10 20 25
r22 23 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.135 $Y=3.59
+ $X2=2.135 $Y2=3.59
r23 20 23 25.3406 $w=5.88e-07 $l=1.25e-06 $layer=LI1_cond $X=1.955 $Y=2.34
+ $X2=1.955 $Y2=3.59
r24 14 17 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.205 $Y=3.63
+ $X2=0.925 $Y2=3.63
r25 13 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.925 $Y=3.59
+ $X2=0.925 $Y2=3.59
r26 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.205 $Y=3.59
+ $X2=0.205 $Y2=3.59
r27 10 13 16.0526 $w=9.48e-07 $l=1.25e-06 $layer=LI1_cond $X=0.565 $Y=2.34
+ $X2=0.565 $Y2=3.59
r28 7 25 0.358952 $w=3.7e-07 $l=9.35e-07 $layer=MET1_cond $X=1.2 $Y=3.63
+ $X2=2.135 $Y2=3.63
r29 7 17 0.105574 $w=3.7e-07 $l=2.75e-07 $layer=MET1_cond $X=1.2 $Y=3.63
+ $X2=0.925 $Y2=3.63
r30 2 23 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.945
+ $Y=2.215 $X2=2.085 $Y2=3.59
r31 2 20 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.945
+ $Y=2.215 $X2=2.085 $Y2=2.34
r32 1 13 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.38
+ $Y=2.215 $X2=0.525 $Y2=3.59
r33 1 10 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.38
+ $Y=2.215 $X2=0.525 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND2_1%Y 1 2 9 13 15 20 22
c35 13 0 1.03339e-19 $X=2.015 $Y=1.175
r36 22 25 0.456684 $w=1.68e-07 $l=7e-09 $layer=LI1_cond $X=1.68 $Y=1.26
+ $X2=1.687 $Y2=1.26
r37 22 25 0.911234 $w=2.13e-07 $l=1.7e-08 $layer=LI1_cond $X=1.687 $Y=1.362
+ $X2=1.687 $Y2=1.345
r38 20 22 8.73713 $w=2.13e-07 $l=1.63e-07 $layer=LI1_cond $X=1.687 $Y=1.525
+ $X2=1.687 $Y2=1.362
r39 13 25 21.3989 $w=1.68e-07 $l=3.28e-07 $layer=LI1_cond $X=2.015 $Y=1.26
+ $X2=1.687 $Y2=1.26
r40 13 15 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.015 $Y=1.175
+ $X2=2.015 $Y2=0.68
r41 9 11 57.6222 $w=2.48e-07 $l=1.25e-06 $layer=LI1_cond $X=1.345 $Y=2.34
+ $X2=1.345 $Y2=3.59
r42 7 20 22.3123 $w=1.68e-07 $l=3.42e-07 $layer=LI1_cond $X=1.345 $Y=1.61
+ $X2=1.687 $Y2=1.61
r43 7 9 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=1.345 $Y=1.695
+ $X2=1.345 $Y2=2.34
r44 2 11 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.165
+ $Y=2.215 $X2=1.305 $Y2=3.59
r45 2 9 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.165
+ $Y=2.215 $X2=1.305 $Y2=2.34
r46 1 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.875
+ $Y=0.555 $X2=2.015 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND2_1%VGND 1 4 7
r13 7 13 1.8626 $w=1.308e-06 $l=2e-07 $layer=LI1_cond $X=0.745 $Y=0.48 $X2=0.745
+ $Y2=0.68
r14 7 8 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.205 $Y=0.48
+ $X2=0.205 $Y2=0.48
r15 4 8 0.381986 $w=3.7e-07 $l=9.95e-07 $layer=MET1_cond $X=1.2 $Y=0.44
+ $X2=0.205 $Y2=0.44
r16 4 7 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.285 $Y=0.48
+ $X2=1.285 $Y2=0.48
r17 1 13 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.38
+ $Y=0.555 $X2=0.525 $Y2=0.68
.ends

