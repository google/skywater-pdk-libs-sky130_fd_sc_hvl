# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__sdfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__sdfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  19.68000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 1.175000 4.675000 2.150000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.611250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.955000 0.495000 16.285000 2.025000 ;
        RECT 15.955000 2.025000 16.545000 2.515000 ;
        RECT 16.215000 2.515000 16.545000 3.455000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.220000 0.495000 19.555000 3.755000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.930000 1.975000 2.440000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.550000 2.755000 1.750000 ;
        RECT 0.565000 1.750000 0.895000 2.220000 ;
        RECT 2.425000 1.750000 2.755000 2.745000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 10.685000 1.895000 11.395000 2.120000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  1.050000 0.365000  2.000000 0.995000 ;
        RECT  3.860000 0.365000  4.785000 0.995000 ;
        RECT  6.175000 0.365000  7.065000 1.075000 ;
        RECT 10.495000 0.365000 11.445000 0.915000 ;
        RECT 13.915000 0.365000 14.865000 1.325000 ;
        RECT 16.465000 0.365000 17.415000 1.325000 ;
        RECT 18.140000 0.365000 19.040000 1.325000 ;
      LAYER mcon ;
        RECT  1.080000 0.395000  1.250000 0.565000 ;
        RECT  1.440000 0.395000  1.610000 0.565000 ;
        RECT  1.800000 0.395000  1.970000 0.565000 ;
        RECT  3.875000 0.395000  4.045000 0.565000 ;
        RECT  4.235000 0.395000  4.405000 0.565000 ;
        RECT  4.595000 0.395000  4.765000 0.565000 ;
        RECT  6.175000 0.395000  6.345000 0.565000 ;
        RECT  6.535000 0.395000  6.705000 0.565000 ;
        RECT  6.895000 0.395000  7.065000 0.565000 ;
        RECT 10.525000 0.395000 10.695000 0.565000 ;
        RECT 10.885000 0.395000 11.055000 0.565000 ;
        RECT 11.245000 0.395000 11.415000 0.565000 ;
        RECT 13.945000 0.395000 14.115000 0.565000 ;
        RECT 14.305000 0.395000 14.475000 0.565000 ;
        RECT 14.665000 0.395000 14.835000 0.565000 ;
        RECT 16.495000 0.395000 16.665000 0.565000 ;
        RECT 16.855000 0.395000 17.025000 0.565000 ;
        RECT 17.215000 0.395000 17.385000 0.565000 ;
        RECT 18.145000 0.395000 18.315000 0.565000 ;
        RECT 18.505000 0.395000 18.675000 0.565000 ;
        RECT 18.865000 0.395000 19.035000 0.565000 ;
      LAYER met1 ;
        RECT 0.000000 0.255000 19.680000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 19.680000 0.085000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
        RECT 15.995000 -0.085000 16.165000 0.085000 ;
        RECT 16.475000 -0.085000 16.645000 0.085000 ;
        RECT 16.955000 -0.085000 17.125000 0.085000 ;
        RECT 17.435000 -0.085000 17.605000 0.085000 ;
        RECT 17.915000 -0.085000 18.085000 0.085000 ;
        RECT 18.395000 -0.085000 18.565000 0.085000 ;
        RECT 18.875000 -0.085000 19.045000 0.085000 ;
        RECT 19.355000 -0.085000 19.525000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.115000 19.680000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 19.680000 4.155000 ;
      LAYER mcon ;
        RECT  0.155000 3.985000  0.325000 4.155000 ;
        RECT  0.635000 3.985000  0.805000 4.155000 ;
        RECT  1.115000 3.985000  1.285000 4.155000 ;
        RECT  1.595000 3.985000  1.765000 4.155000 ;
        RECT  2.075000 3.985000  2.245000 4.155000 ;
        RECT  2.555000 3.985000  2.725000 4.155000 ;
        RECT  3.035000 3.985000  3.205000 4.155000 ;
        RECT  3.515000 3.985000  3.685000 4.155000 ;
        RECT  3.995000 3.985000  4.165000 4.155000 ;
        RECT  4.475000 3.985000  4.645000 4.155000 ;
        RECT  4.955000 3.985000  5.125000 4.155000 ;
        RECT  5.435000 3.985000  5.605000 4.155000 ;
        RECT  5.915000 3.985000  6.085000 4.155000 ;
        RECT  6.395000 3.985000  6.565000 4.155000 ;
        RECT  6.875000 3.985000  7.045000 4.155000 ;
        RECT  7.355000 3.985000  7.525000 4.155000 ;
        RECT  7.835000 3.985000  8.005000 4.155000 ;
        RECT  8.315000 3.985000  8.485000 4.155000 ;
        RECT  8.795000 3.985000  8.965000 4.155000 ;
        RECT  9.275000 3.985000  9.445000 4.155000 ;
        RECT  9.755000 3.985000  9.925000 4.155000 ;
        RECT 10.235000 3.985000 10.405000 4.155000 ;
        RECT 10.715000 3.985000 10.885000 4.155000 ;
        RECT 11.195000 3.985000 11.365000 4.155000 ;
        RECT 11.675000 3.985000 11.845000 4.155000 ;
        RECT 12.155000 3.985000 12.325000 4.155000 ;
        RECT 12.635000 3.985000 12.805000 4.155000 ;
        RECT 13.115000 3.985000 13.285000 4.155000 ;
        RECT 13.595000 3.985000 13.765000 4.155000 ;
        RECT 14.075000 3.985000 14.245000 4.155000 ;
        RECT 14.555000 3.985000 14.725000 4.155000 ;
        RECT 15.035000 3.985000 15.205000 4.155000 ;
        RECT 15.515000 3.985000 15.685000 4.155000 ;
        RECT 15.995000 3.985000 16.165000 4.155000 ;
        RECT 16.475000 3.985000 16.645000 4.155000 ;
        RECT 16.955000 3.985000 17.125000 4.155000 ;
        RECT 17.435000 3.985000 17.605000 4.155000 ;
        RECT 17.915000 3.985000 18.085000 4.155000 ;
        RECT 18.395000 3.985000 18.565000 4.155000 ;
        RECT 18.875000 3.985000 19.045000 4.155000 ;
        RECT 19.355000 3.985000 19.525000 4.155000 ;
      LAYER met1 ;
        RECT 0.000000 3.955000 19.680000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.630000 2.620000  1.220000 3.705000 ;
        RECT  1.750000 3.335000  2.700000 3.755000 ;
        RECT  6.320000 3.465000  7.210000 3.755000 ;
        RECT 10.535000 2.650000 11.125000 3.705000 ;
        RECT 14.520000 2.695000 15.425000 3.735000 ;
        RECT 17.075000 2.025000 17.665000 3.705000 ;
        RECT 18.380000 2.175000 18.970000 3.755000 ;
      LAYER mcon ;
        RECT  0.660000 3.505000  0.830000 3.675000 ;
        RECT  1.020000 3.505000  1.190000 3.675000 ;
        RECT  1.780000 3.505000  1.950000 3.675000 ;
        RECT  2.140000 3.505000  2.310000 3.675000 ;
        RECT  2.500000 3.505000  2.670000 3.675000 ;
        RECT  6.320000 3.505000  6.490000 3.675000 ;
        RECT  6.680000 3.505000  6.850000 3.675000 ;
        RECT  7.040000 3.505000  7.210000 3.675000 ;
        RECT 10.565000 3.505000 10.735000 3.675000 ;
        RECT 10.925000 3.505000 11.095000 3.675000 ;
        RECT 14.525000 3.505000 14.695000 3.675000 ;
        RECT 14.885000 3.505000 15.055000 3.675000 ;
        RECT 15.245000 3.505000 15.415000 3.675000 ;
        RECT 17.105000 3.505000 17.275000 3.675000 ;
        RECT 17.465000 3.505000 17.635000 3.675000 ;
        RECT 18.410000 3.505000 18.580000 3.675000 ;
        RECT 18.770000 3.505000 18.940000 3.675000 ;
      LAYER met1 ;
        RECT 0.000000 3.445000 19.680000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.110000 1.175000  3.330000 1.345000 ;
      RECT  0.110000 1.345000  0.280000 2.555000 ;
      RECT  0.110000 2.555000  0.440000 3.015000 ;
      RECT  0.540000 0.495000  0.870000 1.175000 ;
      RECT  1.400000 2.925000  3.680000 3.095000 ;
      RECT  1.400000 3.095000  1.570000 3.755000 ;
      RECT  2.810000 0.495000  3.140000 0.825000 ;
      RECT  2.810000 0.825000  3.680000 0.995000 ;
      RECT  2.880000 3.275000  3.210000 3.610000 ;
      RECT  2.880000 3.610000  4.030000 3.780000 ;
      RECT  3.065000 1.345000  3.330000 1.845000 ;
      RECT  3.430000 3.095000  3.680000 3.430000 ;
      RECT  3.510000 0.995000  3.680000 2.330000 ;
      RECT  3.510000 2.330000  5.135000 2.500000 ;
      RECT  3.860000 2.680000  5.240000 2.850000 ;
      RECT  3.860000 2.850000  4.030000 3.610000 ;
      RECT  4.210000 3.030000  4.540000 3.635000 ;
      RECT  4.210000 3.635000  6.140000 3.805000 ;
      RECT  4.965000 0.265000  5.995000 0.435000 ;
      RECT  4.965000 0.435000  5.135000 2.330000 ;
      RECT  4.990000 2.850000  5.240000 3.430000 ;
      RECT  5.315000 0.615000  5.645000 1.605000 ;
      RECT  5.315000 1.605000  7.120000 1.775000 ;
      RECT  5.420000 1.775000  5.790000 3.455000 ;
      RECT  5.825000 0.435000  5.995000 1.255000 ;
      RECT  5.825000 1.255000  8.165000 1.425000 ;
      RECT  5.970000 1.955000  7.470000 2.125000 ;
      RECT  5.970000 2.125000  6.140000 3.115000 ;
      RECT  5.970000 3.115000  7.560000 3.285000 ;
      RECT  5.970000 3.285000  6.140000 3.635000 ;
      RECT  6.320000 2.305000  7.910000 2.555000 ;
      RECT  7.245000 0.590000  9.725000 0.760000 ;
      RECT  7.245000 0.760000  7.575000 1.075000 ;
      RECT  7.300000 1.425000  7.470000 1.955000 ;
      RECT  7.390000 3.285000  9.435000 3.455000 ;
      RECT  7.740000 2.135000  8.785000 2.305000 ;
      RECT  7.740000 2.555000  7.910000 2.855000 ;
      RECT  7.740000 2.855000  8.655000 3.105000 ;
      RECT  7.835000 0.940000  8.165000 1.255000 ;
      RECT  8.090000 2.485000  9.005000 2.675000 ;
      RECT  8.615000 0.940000  8.945000 1.360000 ;
      RECT  8.615000 1.360000  8.785000 2.135000 ;
      RECT  8.835000 2.675000  9.005000 2.750000 ;
      RECT  8.835000 2.750000 10.355000 2.920000 ;
      RECT  9.070000 1.545000 12.130000 1.715000 ;
      RECT  9.070000 1.715000  9.400000 2.215000 ;
      RECT  9.105000 3.100000  9.435000 3.285000 ;
      RECT  9.395000 0.760000  9.725000 1.360000 ;
      RECT  9.675000 1.715000  9.845000 2.320000 ;
      RECT  9.675000 2.320000 10.005000 2.570000 ;
      RECT  9.985000 0.495000 10.315000 1.545000 ;
      RECT 10.025000 1.895000 10.355000 2.140000 ;
      RECT 10.185000 2.140000 10.355000 2.300000 ;
      RECT 10.185000 2.300000 11.565000 2.470000 ;
      RECT 10.185000 2.470000 10.355000 2.750000 ;
      RECT 10.495000 1.095000 11.875000 1.265000 ;
      RECT 10.495000 1.265000 10.825000 1.365000 ;
      RECT 11.315000 2.470000 11.565000 3.110000 ;
      RECT 11.625000 0.475000 13.610000 0.645000 ;
      RECT 11.625000 0.645000 11.875000 1.095000 ;
      RECT 11.785000 2.205000 12.115000 3.635000 ;
      RECT 11.785000 3.635000 14.340000 3.805000 ;
      RECT 11.800000 1.445000 12.130000 1.545000 ;
      RECT 11.800000 1.715000 12.130000 2.025000 ;
      RECT 12.150000 0.825000 12.480000 1.245000 ;
      RECT 12.310000 1.245000 12.480000 3.285000 ;
      RECT 12.310000 3.285000 13.795000 3.455000 ;
      RECT 12.660000 2.205000 12.990000 3.105000 ;
      RECT 12.820000 0.825000 13.260000 1.325000 ;
      RECT 12.820000 1.325000 12.990000 1.915000 ;
      RECT 12.820000 1.915000 15.135000 2.085000 ;
      RECT 12.820000 2.085000 12.990000 2.205000 ;
      RECT 13.280000 1.505000 13.610000 1.735000 ;
      RECT 13.440000 0.645000 13.610000 1.505000 ;
      RECT 13.440000 2.265000 13.795000 3.285000 ;
      RECT 14.010000 2.695000 14.340000 3.635000 ;
      RECT 14.465000 2.265000 15.775000 2.515000 ;
      RECT 14.805000 1.545000 15.135000 1.915000 ;
      RECT 15.315000 0.495000 15.775000 2.265000 ;
      RECT 15.605000 2.515000 15.775000 2.695000 ;
      RECT 15.605000 2.695000 15.995000 3.635000 ;
      RECT 15.605000 3.635000 16.895000 3.805000 ;
      RECT 16.725000 1.505000 17.055000 1.835000 ;
      RECT 16.725000 1.835000 16.895000 3.635000 ;
      RECT 17.630000 0.495000 17.960000 1.505000 ;
      RECT 17.630000 1.505000 19.040000 1.675000 ;
      RECT 17.870000 2.025000 18.200000 2.815000 ;
      RECT 18.030000 1.675000 19.040000 1.835000 ;
      RECT 18.030000 1.835000 18.200000 2.025000 ;
    LAYER mcon ;
      RECT  5.435000 3.060000  5.605000 3.230000 ;
      RECT 13.595000 3.060000 13.765000 3.230000 ;
    LAYER met1 ;
      RECT  5.375000 3.030000  5.665000 3.075000 ;
      RECT  5.375000 3.075000 13.825000 3.215000 ;
      RECT  5.375000 3.215000  5.665000 3.260000 ;
      RECT 13.535000 3.030000 13.825000 3.075000 ;
      RECT 13.535000 3.215000 13.825000 3.260000 ;
  END
END sky130_fd_sc_hvl__sdfxbp_1
