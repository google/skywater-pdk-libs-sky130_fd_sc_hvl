# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__sdfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__sdfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.88000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 2.205000 2.755000 2.520000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.660000 0.615000 14.020000 1.505000 ;
        RECT 13.660000 2.195000 14.020000 3.735000 ;
        RECT 13.850000 1.505000 14.755000 1.780000 ;
        RECT 13.850000 1.780000 14.020000 2.195000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.600000 2.215000 4.195000 2.765000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.445000 1.795000 1.855000 ;
        RECT 0.605000 1.855000 3.050000 2.025000 ;
        RECT 2.720000 1.095000 3.050000 1.855000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.345000 1.175000 4.675000 1.685000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 14.880000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 14.880000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 14.880000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 14.880000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.880000 0.085000 ;
      RECT  0.000000  3.985000 14.880000 4.155000 ;
      RECT  0.125000  0.515000  0.455000 1.095000 ;
      RECT  0.125000  1.095000  2.305000 1.265000 ;
      RECT  0.125000  1.265000  0.380000 3.425000 ;
      RECT  0.905000  0.365000  1.855000 0.915000 ;
      RECT  0.910000  2.925000  1.860000 3.705000 ;
      RECT  1.975000  1.265000  2.305000 1.675000 ;
      RECT  2.395000  0.495000  2.725000 0.745000 ;
      RECT  2.395000  0.745000  3.400000 0.915000 ;
      RECT  2.400000  2.925000  3.400000 3.095000 ;
      RECT  2.400000  3.095000  2.730000 3.425000 ;
      RECT  3.230000  0.915000  3.400000 1.865000 ;
      RECT  3.230000  1.865000  6.780000 2.035000 ;
      RECT  3.230000  2.035000  3.400000 2.925000 ;
      RECT  3.580000  0.365000  4.485000 0.995000 ;
      RECT  3.635000  2.945000  4.585000 3.735000 ;
      RECT  4.665000  0.515000  5.025000 0.975000 ;
      RECT  4.765000  2.595000  5.605000 2.765000 ;
      RECT  4.765000  2.765000  5.095000 3.735000 ;
      RECT  4.855000  0.975000  5.025000 1.155000 ;
      RECT  4.855000  1.155000  5.870000 1.325000 ;
      RECT  5.215000  0.365000  5.805000 0.975000 ;
      RECT  5.275000  2.215000  5.605000 2.595000 ;
      RECT  5.315000  2.945000  5.905000 3.735000 ;
      RECT  5.540000  1.325000  5.870000 1.685000 ;
      RECT  5.995000  0.265000  8.210000 0.435000 ;
      RECT  5.995000  0.435000  6.325000 0.975000 ;
      RECT  6.095000  2.945000  6.425000 3.335000 ;
      RECT  6.095000  3.335000  7.325000 3.505000 ;
      RECT  6.095000  3.505000  6.425000 3.735000 ;
      RECT  6.565000  0.615000  6.895000 0.995000 ;
      RECT  6.565000  0.995000  6.780000 1.865000 ;
      RECT  6.610000  2.035000  6.780000 2.695000 ;
      RECT  6.610000  2.695000  6.975000 3.155000 ;
      RECT  6.960000  2.225000  7.325000 2.515000 ;
      RECT  7.075000  0.435000  7.245000 2.225000 ;
      RECT  7.155000  2.515000  7.325000 3.335000 ;
      RECT  7.425000  0.615000  7.755000 0.995000 ;
      RECT  7.505000  0.995000  7.755000 1.605000 ;
      RECT  7.505000  1.605000  9.685000 1.775000 ;
      RECT  7.505000  1.775000  7.675000 2.675000 ;
      RECT  7.505000  2.675000  7.755000 3.175000 ;
      RECT  7.880000  1.955000  8.210000 2.495000 ;
      RECT  7.935000  0.435000  8.210000 1.255000 ;
      RECT  7.935000  1.255000 10.295000 1.425000 ;
      RECT  8.040000  2.495000  8.210000 3.155000 ;
      RECT  8.040000  3.155000 10.490000 3.325000 ;
      RECT  8.620000  1.955000 10.645000 2.125000 ;
      RECT  8.620000  2.125000  8.950000 2.555000 ;
      RECT  8.680000  0.365000  9.630000 1.075000 ;
      RECT  9.030000  3.505000  9.980000 3.755000 ;
      RECT  9.810000  0.495000 10.140000 0.905000 ;
      RECT  9.810000  0.905000 10.645000 1.075000 ;
      RECT  9.810000  2.125000  9.980000 2.675000 ;
      RECT  9.810000  2.675000 10.140000 2.975000 ;
      RECT 10.045000  1.425000 10.295000 1.775000 ;
      RECT 10.160000  2.305000 10.490000 2.495000 ;
      RECT 10.320000  2.495000 10.490000 3.155000 ;
      RECT 10.320000  3.325000 11.450000 3.495000 ;
      RECT 10.475000  1.075000 10.645000 1.955000 ;
      RECT 10.670000  2.675000 11.075000 3.145000 ;
      RECT 10.825000  0.495000 11.800000 0.665000 ;
      RECT 10.825000  0.665000 11.075000 2.675000 ;
      RECT 11.255000  1.085000 11.450000 3.325000 ;
      RECT 11.630000  0.665000 11.800000 2.345000 ;
      RECT 11.630000  2.345000 12.930000 2.515000 ;
      RECT 11.980000  0.365000 12.930000 1.305000 ;
      RECT 11.980000  1.485000 13.440000 1.655000 ;
      RECT 11.980000  1.655000 12.310000 2.155000 ;
      RECT 11.980000  2.695000 12.930000 3.735000 ;
      RECT 12.600000  1.845000 12.930000 2.345000 ;
      RECT 13.110000  0.515000 13.440000 1.485000 ;
      RECT 13.110000  1.655000 13.440000 1.685000 ;
      RECT 13.110000  1.685000 13.670000 2.015000 ;
      RECT 13.110000  2.015000 13.440000 3.735000 ;
      RECT 14.200000  0.365000 14.790000 1.325000 ;
      RECT 14.200000  2.195000 14.790000 3.735000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.935000  0.395000  1.105000 0.565000 ;
      RECT  0.940000  3.505000  1.110000 3.675000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.295000  0.395000  1.465000 0.565000 ;
      RECT  1.300000  3.505000  1.470000 3.675000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  1.655000  0.395000  1.825000 0.565000 ;
      RECT  1.660000  3.505000  1.830000 3.675000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.590000  0.395000  3.760000 0.565000 ;
      RECT  3.665000  3.505000  3.835000 3.675000 ;
      RECT  3.950000  0.395000  4.120000 0.565000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.025000  3.505000  4.195000 3.675000 ;
      RECT  4.310000  0.395000  4.480000 0.565000 ;
      RECT  4.385000  3.505000  4.555000 3.675000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.245000  0.395000  5.415000 0.565000 ;
      RECT  5.345000  3.505000  5.515000 3.675000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.605000  0.395000  5.775000 0.565000 ;
      RECT  5.705000  3.505000  5.875000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.710000  0.395000  8.880000 0.565000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.060000  3.535000  9.230000 3.705000 ;
      RECT  9.070000  0.395000  9.240000 0.565000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.420000  3.535000  9.590000 3.705000 ;
      RECT  9.430000  0.395000  9.600000 0.565000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.780000  3.535000  9.950000 3.705000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.010000  0.395000 12.180000 0.565000 ;
      RECT 12.010000  3.505000 12.180000 3.675000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.370000  0.395000 12.540000 0.565000 ;
      RECT 12.370000  3.505000 12.540000 3.675000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 12.730000  0.395000 12.900000 0.565000 ;
      RECT 12.730000  3.505000 12.900000 3.675000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.230000  0.395000 14.400000 0.565000 ;
      RECT 14.230000  3.505000 14.400000 3.675000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.590000  0.395000 14.760000 0.565000 ;
      RECT 14.590000  3.505000 14.760000 3.675000 ;
  END
END sky130_fd_sc_hvl__sdfxtp_1
END LIBRARY
