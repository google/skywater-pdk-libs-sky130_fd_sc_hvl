* File: sky130_fd_sc_hvl__lsbufhv2lv_1.spice
* Created: Fri Aug 28 09:36:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__lsbufhv2lv_1.pex.spice"
.subckt sky130_fd_sc_hvl__lsbufhv2lv_1  VNB VPB LVPWR A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* LVPWR	LVPWR
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_389_141#_M1011_g N_X_M1011_s N_VNB_M1011_b NSHORT
+ L=0.15 W=0.74 AD=0.1961 AS=0.1961 PD=2.01 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_30_1337#_M1002_g N_A_30_207#_M1002_s N_VNB_M1011_b NHV
+ L=0.5 W=0.42 AD=0.128423 AS=0.1197 PD=0.904615 PS=1.41 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g N_A_30_1337#_M1009_s N_VNB_M1011_b NHV L=0.5
+ W=0.42 AD=0.128423 AS=0.1197 PD=0.904615 PS=1.41 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250003 A=0.21 P=1.84 MULT=1
MM1004 N_VGND_M1002_d N_A_30_207#_M1004_g N_A_389_141#_M1004_s N_VNB_M1011_b NHV
+ L=0.5 W=0.75 AD=0.229327 AS=0.105 PD=1.61538 PS=1.03 NRD=17.4762 NRS=0 M=1
+ R=1.5 SA=250001 SB=250001 A=0.375 P=2.5 MULT=1
MM1005 N_A_389_1337#_M1005_d N_A_30_1337#_M1005_g N_VGND_M1009_d N_VNB_M1011_b
+ NHV L=0.5 W=0.75 AD=0.105 AS=0.229327 PD=1.03 PS=1.61538 NRD=0 NRS=17.4762 M=1
+ R=1.5 SA=250001 SB=250002 A=0.375 P=2.5 MULT=1
MM1006 N_VGND_M1006_d N_A_30_207#_M1006_g N_A_389_141#_M1004_s N_VNB_M1011_b NHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1007 N_VGND_M1007_d N_A_30_207#_M1007_g N_A_389_141#_M1007_s N_VNB_M1011_b NHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1010 N_VGND_M1010_d N_A_30_207#_M1010_g N_A_389_141#_M1010_s N_VNB_M1011_b NHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1008 N_A_389_1337#_M1008_d N_A_30_1337#_M1008_g N_VGND_M1008_s N_VNB_M1011_b
+ NHV L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1012 N_A_389_1337#_M1005_d N_A_30_1337#_M1012_g N_VGND_M1012_s N_VNB_M1011_b
+ NHV L=0.5 W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250001 A=0.375 P=2.5 MULT=1
MM1014 N_A_389_1337#_M1014_d N_A_30_1337#_M1014_g N_VGND_M1012_s N_VNB_M1011_b
+ NHV L=0.5 W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250002 SB=250000 A=0.375 P=2.5 MULT=1
MM1003 N_LVPWR_M1003_d N_A_389_141#_M1003_g N_X_M1003_s N_LVPWR_M1003_b PHIGHVT
+ L=0.15 W=1.12 AD=0.1568 AS=0.2968 PD=1.4 PS=2.77 NRD=0 NRS=0 M=1 R=7.46667
+ SA=75000.2 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1001 N_LVPWR_M1001_d N_A_389_1337#_M1001_g N_A_389_141#_M1001_s
+ N_LVPWR_M1003_b PHIGHVT L=0.15 W=1.12 AD=0.2968 AS=0.2968 PD=2.77 PS=2.77
+ NRD=0 NRS=0 M=1 R=7.46667 SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1013 N_A_389_1337#_M1013_d N_A_389_141#_M1013_g N_LVPWR_M1003_d
+ N_LVPWR_M1003_b PHIGHVT L=0.15 W=1.12 AD=0.2968 AS=0.1568 PD=2.77 PS=1.4 NRD=0
+ NRS=0 M=1 R=7.46667 SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1015 N_A_30_207#_M1015_d N_A_30_1337#_M1015_g N_VPWR_M1015_s N_VPB_M1015_b PHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.1197 PD=1.37 PS=1.41 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1000 N_A_30_1337#_M1000_d N_A_M1000_g N_VPWR_M1000_s N_VPB_M1015_b PHV L=0.5
+ W=0.42 AD=0.1113 AS=0.1197 PD=1.37 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250000 A=0.21 P=1.84 MULT=1
DX16_noxref N_VNB_M1011_b N_VPB_M1015_b NWDIODE A=8.1282 P=12.46
DX17_noxref N_VNB_M1011_b N_LVPWR_M1003_b NWDIODE A=5.3655 P=10.24
DX18_noxref N_VNB_M1011_b N_VPB_X18_noxref_D1 NWDIODE A=6.5113 P=11.72
*
.include "sky130_fd_sc_hvl__lsbufhv2lv_1.pxi.spice"
*
.ends
*
*
