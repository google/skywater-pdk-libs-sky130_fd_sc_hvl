* File: sky130_fd_sc_hvl__buf_2.spice
* Created: Fri Aug 28 09:33:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__buf_2.pex.spice"
.subckt sky130_fd_sc_hvl__buf_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_X_M1002_d N_A_129_279#_M1002_g N_VGND_M1002_s N_VNB_M1002_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.21375 PD=1.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1005 N_X_M1002_d N_A_129_279#_M1005_g N_VGND_M1005_s N_VNB_M1002_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.194904 PD=1.03 PS=1.60256 NRD=0 NRS=0 M=1 R=1.5 SA=250001
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1004 N_A_129_279#_M1004_d N_A_M1004_g N_VGND_M1005_s N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.109146 PD=1.37 PS=0.897436 NRD=0 NRS=59.7132 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1001 N_X_M1001_d N_A_129_279#_M1001_g N_VPWR_M1001_s N_VPB_M1001_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.4275 PD=1.78 PS=3.57 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250001 A=0.75 P=4 MULT=1
MM1003 N_X_M1001_d N_A_129_279#_M1003_g N_VPWR_M1003_s N_VPB_M1001_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.3925 PD=1.78 PS=2.66667 NRD=0 NRS=0 M=1 R=3 SA=250001
+ SB=250001 A=0.75 P=4 MULT=1
MM1000 N_A_129_279#_M1000_d N_A_M1000_g N_VPWR_M1003_s N_VPB_M1001_b PHV L=0.5
+ W=0.75 AD=0.21375 AS=0.19625 PD=2.07 PS=1.33333 NRD=0 NRS=56.0203 M=1 R=1.5
+ SA=250002 SB=250000 A=0.375 P=2.5 MULT=1
DX6_noxref N_VNB_M1002_b N_VPB_M1001_b NWDIODE A=10.452 P=13.24
*
.include "sky130_fd_sc_hvl__buf_2.pxi.spice"
*
.ends
*
*
