* NGSPICE file created from sky130_fd_sc_hvl__lsbufhv2hv_hl_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__lsbufhv2hv_hl_1 A LOWHVPWR VGND VNB VPB VPWR X
M1000 a_762_107# a_662_81# X VNB nhv w=750000u l=500000u
+  ad=3.0405e+11p pd=2.5e+06u as=1.9875e+11p ps=2.03e+06u
M1001 a_662_81# A LOWHVPWR LOWHVPWR phv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=5.1e+11p ps=3.79e+06u
M1002 a_662_81# A a_762_107# VNB nhv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1003 LOWHVPWR a_662_81# X LOWHVPWR phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=4.275e+11p ps=3.57e+06u
.ends

