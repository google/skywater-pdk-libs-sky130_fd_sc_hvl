* File: sky130_fd_sc_hvl__sdlxtp_1.pxi.spice
* Created: Fri Aug 28 09:40:44 2020
* 
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%VNB N_VNB_M1004_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__SDLXTP_1%VNB
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%VPB N_VPB_M1018_b VPB N_VPB_c_95_p VPB
+ PM_SKY130_FD_SC_HVL__SDLXTP_1%VPB
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%SCE N_SCE_M1018_g N_SCE_M1004_g N_SCE_c_218_n
+ N_SCE_M1010_g N_SCE_M1008_g N_SCE_c_211_n N_SCE_c_212_n N_SCE_c_213_n
+ N_SCE_c_214_n N_SCE_c_215_n SCE SCE SCE N_SCE_c_222_n N_SCE_c_216_n
+ N_SCE_c_226_n N_SCE_c_217_n PM_SKY130_FD_SC_HVL__SDLXTP_1%SCE
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%A_30_587# N_A_30_587#_M1004_s
+ N_A_30_587#_M1018_s N_A_30_587#_c_285_n N_A_30_587#_c_287_n
+ N_A_30_587#_c_288_n N_A_30_587#_c_289_n N_A_30_587#_c_290_n
+ N_A_30_587#_c_311_n N_A_30_587#_c_296_n N_A_30_587#_c_297_n
+ N_A_30_587#_c_291_n N_A_30_587#_M1016_g N_A_30_587#_M1003_g
+ PM_SKY130_FD_SC_HVL__SDLXTP_1%A_30_587#
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%D N_D_M1015_g N_D_M1017_g D D D N_D_c_375_n
+ N_D_c_384_n PM_SKY130_FD_SC_HVL__SDLXTP_1%D
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%SCD N_SCD_M1009_g N_SCD_c_412_n SCD SCD SCD
+ N_SCD_c_413_n N_SCD_M1012_g PM_SKY130_FD_SC_HVL__SDLXTP_1%SCD
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%GATE N_GATE_M1006_g N_GATE_M1023_g
+ N_GATE_c_455_n GATE GATE GATE GATE N_GATE_c_453_n N_GATE_c_454_n
+ PM_SKY130_FD_SC_HVL__SDLXTP_1%GATE
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%A_1214_107# N_A_1214_107#_M1005_d
+ N_A_1214_107#_M1014_d N_A_1214_107#_c_501_n N_A_1214_107#_M1000_g
+ N_A_1214_107#_c_491_n N_A_1214_107#_c_505_n N_A_1214_107#_c_492_n
+ N_A_1214_107#_c_494_n N_A_1214_107#_c_516_p N_A_1214_107#_c_496_n
+ N_A_1214_107#_c_512_p N_A_1214_107#_c_519_p N_A_1214_107#_c_506_n
+ N_A_1214_107#_c_507_n N_A_1214_107#_c_497_n N_A_1214_107#_c_498_n
+ N_A_1214_107#_M1002_g PM_SKY130_FD_SC_HVL__SDLXTP_1%A_1214_107#
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%A_944_107# N_A_944_107#_M1006_d
+ N_A_944_107#_M1023_d N_A_944_107#_c_593_n N_A_944_107#_M1014_g
+ N_A_944_107#_c_596_n N_A_944_107#_c_582_n N_A_944_107#_M1007_g
+ N_A_944_107#_M1019_g N_A_944_107#_c_601_n N_A_944_107#_c_585_n
+ N_A_944_107#_c_586_n N_A_944_107#_c_587_n N_A_944_107#_c_588_n
+ N_A_944_107#_c_590_n N_A_944_107#_c_633_n N_A_944_107#_M1005_g
+ PM_SKY130_FD_SC_HVL__SDLXTP_1%A_944_107#
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%A_1678_81# N_A_1678_81#_M1013_s
+ N_A_1678_81#_M1011_s N_A_1678_81#_c_693_n N_A_1678_81#_M1022_g
+ N_A_1678_81#_M1001_g N_A_1678_81#_c_695_n N_A_1678_81#_c_696_n
+ N_A_1678_81#_c_702_n N_A_1678_81#_c_697_n N_A_1678_81#_c_703_n
+ N_A_1678_81#_c_710_n N_A_1678_81#_c_704_n N_A_1678_81#_c_698_n
+ N_A_1678_81#_c_699_n PM_SKY130_FD_SC_HVL__SDLXTP_1%A_1678_81#
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%A_1480_107# N_A_1480_107#_M1002_d
+ N_A_1480_107#_M1007_d N_A_1480_107#_M1011_g N_A_1480_107#_M1013_g
+ N_A_1480_107#_M1021_g N_A_1480_107#_M1020_g N_A_1480_107#_c_773_n
+ N_A_1480_107#_c_787_n N_A_1480_107#_c_788_n N_A_1480_107#_c_775_n
+ N_A_1480_107#_c_776_n N_A_1480_107#_c_791_n N_A_1480_107#_c_777_n
+ N_A_1480_107#_c_778_n N_A_1480_107#_c_779_n N_A_1480_107#_c_794_n
+ N_A_1480_107#_c_780_n N_A_1480_107#_c_853_n N_A_1480_107#_c_781_n
+ N_A_1480_107#_c_782_n PM_SKY130_FD_SC_HVL__SDLXTP_1%A_1480_107#
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%VPWR N_VPWR_M1018_d N_VPWR_M1012_d
+ N_VPWR_M1014_s N_VPWR_M1001_d N_VPWR_M1011_d VPWR N_VPWR_c_893_n
+ N_VPWR_c_896_n N_VPWR_c_899_n N_VPWR_c_902_n N_VPWR_c_905_n N_VPWR_c_908_n
+ PM_SKY130_FD_SC_HVL__SDLXTP_1%VPWR
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%A_489_107# N_A_489_107#_M1016_d
+ N_A_489_107#_M1002_s N_A_489_107#_M1017_d N_A_489_107#_M1007_s
+ N_A_489_107#_c_991_n N_A_489_107#_c_984_n N_A_489_107#_c_994_n
+ N_A_489_107#_c_995_n N_A_489_107#_c_1019_n N_A_489_107#_c_985_n
+ N_A_489_107#_c_1028_n N_A_489_107#_c_986_n N_A_489_107#_c_997_n
+ N_A_489_107#_c_1049_n N_A_489_107#_c_998_n N_A_489_107#_c_1001_n
+ N_A_489_107#_c_1003_n N_A_489_107#_c_1004_n N_A_489_107#_c_1005_n
+ N_A_489_107#_c_1006_n N_A_489_107#_c_1007_n N_A_489_107#_c_1010_n
+ N_A_489_107#_c_1013_n N_A_489_107#_c_987_n N_A_489_107#_c_1014_n
+ N_A_489_107#_c_989_n N_A_489_107#_c_1015_n N_A_489_107#_c_990_n
+ PM_SKY130_FD_SC_HVL__SDLXTP_1%A_489_107#
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%Q N_Q_M1020_d N_Q_M1021_d Q Q Q Q Q Q Q
+ N_Q_c_1137_n PM_SKY130_FD_SC_HVL__SDLXTP_1%Q
x_PM_SKY130_FD_SC_HVL__SDLXTP_1%VGND N_VGND_M1004_d N_VGND_M1009_d
+ N_VGND_M1005_s N_VGND_M1022_d N_VGND_M1013_d VGND N_VGND_c_1152_n
+ N_VGND_c_1154_n N_VGND_c_1156_n N_VGND_c_1158_n N_VGND_c_1160_n
+ N_VGND_c_1162_n PM_SKY130_FD_SC_HVL__SDLXTP_1%VGND
cc_1 N_VNB_M1004_b N_SCE_M1004_g 0.0469269f $X=-0.33 $Y=-0.265 $X2=0.705
+ $Y2=0.745
cc_2 N_VNB_c_2_p N_SCE_M1004_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.705 $Y2=0.745
cc_3 N_VNB_M1004_b N_SCE_M1008_g 0.0468022f $X=-0.33 $Y=-0.265 $X2=2.975
+ $Y2=0.745
cc_4 N_VNB_c_2_p N_SCE_M1008_g 0.0023273f $X=0.24 $Y=0 $X2=2.975 $Y2=0.745
cc_5 N_VNB_M1004_b N_SCE_c_211_n 0.0507418f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=1.585
cc_6 N_VNB_M1004_b N_SCE_c_212_n 0.00867929f $X=-0.33 $Y=-0.265 $X2=2.6 $Y2=1.92
cc_7 N_VNB_M1004_b N_SCE_c_213_n 0.00548442f $X=-0.33 $Y=-0.265 $X2=2.685
+ $Y2=1.835
cc_8 N_VNB_M1004_b N_SCE_c_214_n 0.00262112f $X=-0.33 $Y=-0.265 $X2=2.82
+ $Y2=1.53
cc_9 N_VNB_M1004_b N_SCE_c_215_n 0.0645996f $X=-0.33 $Y=-0.265 $X2=2.82 $Y2=1.53
cc_10 N_VNB_M1004_b N_SCE_c_216_n 0.0289088f $X=-0.33 $Y=-0.265 $X2=0.75
+ $Y2=2.27
cc_11 N_VNB_M1004_b N_SCE_c_217_n 0.0052153f $X=-0.33 $Y=-0.265 $X2=1.795
+ $Y2=2.305
cc_12 N_VNB_M1004_b N_A_30_587#_c_285_n 0.0360511f $X=-0.33 $Y=-0.265 $X2=1.56
+ $Y2=3.31
cc_13 N_VNB_c_2_p N_A_30_587#_c_285_n 8.66888e-19 $X=0.24 $Y=0 $X2=1.56 $Y2=3.31
cc_14 N_VNB_M1004_b N_A_30_587#_c_287_n 0.0285069f $X=-0.33 $Y=-0.265 $X2=2.975
+ $Y2=0.745
cc_15 N_VNB_M1004_b N_A_30_587#_c_288_n 0.0123137f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=1.585
cc_16 N_VNB_M1004_b N_A_30_587#_c_289_n 0.00648436f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=1.585
cc_17 N_VNB_M1004_b N_A_30_587#_c_290_n 0.00994965f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1004_b N_A_30_587#_c_291_n 0.00678108f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.425
cc_19 N_VNB_M1004_b N_A_30_587#_M1016_g 0.113954f $X=-0.33 $Y=-0.265 $X2=0.75
+ $Y2=2.27
cc_20 N_VNB_c_2_p N_A_30_587#_M1016_g 0.0023273f $X=0.24 $Y=0 $X2=0.75 $Y2=2.27
cc_21 N_VNB_M1004_b N_D_M1015_g 0.114444f $X=-0.33 $Y=-0.265 $X2=0.685 $Y2=3.145
cc_22 N_VNB_c_2_p N_D_M1015_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.685 $Y2=3.145
cc_23 N_VNB_M1004_b N_SCD_M1009_g 0.0467133f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=3.145
cc_24 N_VNB_c_2_p N_SCD_M1009_g 0.00200614f $X=0.24 $Y=0 $X2=0.685 $Y2=3.145
cc_25 N_VNB_M1004_b N_SCD_c_412_n 0.0522425f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_26 N_VNB_M1004_b N_SCD_c_413_n 0.0278019f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=1.585
cc_27 N_VNB_M1004_b N_GATE_M1006_g 0.048209f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=3.145
cc_28 N_VNB_c_2_p N_GATE_M1006_g 0.00123813f $X=0.24 $Y=0 $X2=0.685 $Y2=3.145
cc_29 N_VNB_M1004_b N_GATE_c_453_n 0.0522482f $X=-0.33 $Y=-0.265 $X2=2.685
+ $Y2=1.695
cc_30 N_VNB_M1004_b N_GATE_c_454_n 0.0307656f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_31 N_VNB_M1004_b N_A_1214_107#_c_491_n 0.00488841f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_32 N_VNB_M1004_b N_A_1214_107#_c_492_n 0.0669937f $X=-0.33 $Y=-0.265
+ $X2=2.685 $Y2=1.835
cc_33 N_VNB_c_2_p N_A_1214_107#_c_492_n 0.00289338f $X=0.24 $Y=0 $X2=2.685
+ $Y2=1.835
cc_34 N_VNB_M1004_b N_A_1214_107#_c_494_n 0.0288875f $X=-0.33 $Y=-0.265
+ $X2=2.685 $Y2=1.57
cc_35 N_VNB_c_2_p N_A_1214_107#_c_494_n 0.00122664f $X=0.24 $Y=0 $X2=2.685
+ $Y2=1.57
cc_36 N_VNB_M1004_b N_A_1214_107#_c_496_n 0.0058657f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=2.32
cc_37 N_VNB_M1004_b N_A_1214_107#_c_497_n 0.00912578f $X=-0.33 $Y=-0.265
+ $X2=0.75 $Y2=2.27
cc_38 N_VNB_M1004_b N_A_1214_107#_c_498_n 0.0212012f $X=-0.33 $Y=-0.265
+ $X2=0.685 $Y2=2.625
cc_39 N_VNB_M1004_b N_A_1214_107#_M1002_g 0.122116f $X=-0.33 $Y=-0.265 $X2=0.75
+ $Y2=2.61
cc_40 N_VNB_c_2_p N_A_1214_107#_M1002_g 5.98017e-19 $X=0.24 $Y=0 $X2=0.75
+ $Y2=2.61
cc_41 N_VNB_M1004_b N_A_944_107#_c_582_n 0.0450477f $X=-0.33 $Y=-0.265 $X2=2.975
+ $Y2=0.745
cc_42 N_VNB_M1004_b N_A_944_107#_M1019_g 0.0800738f $X=-0.33 $Y=-0.265 $X2=2.6
+ $Y2=1.92
cc_43 N_VNB_c_2_p N_A_944_107#_M1019_g 0.0023273f $X=0.24 $Y=0 $X2=2.6 $Y2=1.92
cc_44 N_VNB_M1004_b N_A_944_107#_c_585_n 0.00516217f $X=-0.33 $Y=-0.265 $X2=2.82
+ $Y2=1.57
cc_45 N_VNB_M1004_b N_A_944_107#_c_586_n 0.0122361f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_M1004_b N_A_944_107#_c_587_n 0.0276223f $X=-0.33 $Y=-0.265 $X2=1.115
+ $Y2=2.32
cc_47 N_VNB_M1004_b N_A_944_107#_c_588_n 0.017505f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.425
cc_48 N_VNB_c_2_p N_A_944_107#_c_588_n 7.96506e-19 $X=0.24 $Y=0 $X2=0.685
+ $Y2=2.425
cc_49 N_VNB_M1004_b N_A_944_107#_c_590_n 0.00209233f $X=-0.33 $Y=-0.265 $X2=0.75
+ $Y2=2.27
cc_50 N_VNB_M1004_b N_A_944_107#_M1005_g 0.139526f $X=-0.33 $Y=-0.265 $X2=1.34
+ $Y2=2.625
cc_51 N_VNB_c_2_p N_A_944_107#_M1005_g 0.00116831f $X=0.24 $Y=0 $X2=1.34
+ $Y2=2.625
cc_52 N_VNB_M1004_b N_A_1678_81#_c_693_n 0.0397912f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_53 N_VNB_M1004_b N_A_1678_81#_M1001_g 0.0130479f $X=-0.33 $Y=-0.265 $X2=2.975
+ $Y2=0.745
cc_54 N_VNB_M1004_b N_A_1678_81#_c_695_n 0.003789f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_55 N_VNB_M1004_b N_A_1678_81#_c_696_n 0.0102722f $X=-0.33 $Y=-0.265 $X2=2.6
+ $Y2=1.92
cc_56 N_VNB_M1004_b N_A_1678_81#_c_697_n 0.003199f $X=-0.33 $Y=-0.265 $X2=2.685
+ $Y2=1.57
cc_57 N_VNB_M1004_b N_A_1678_81#_c_698_n 0.00302906f $X=-0.33 $Y=-0.265 $X2=0.75
+ $Y2=2.27
cc_58 N_VNB_M1004_b N_A_1678_81#_c_699_n 0.119952f $X=-0.33 $Y=-0.265 $X2=0.75
+ $Y2=2.61
cc_59 N_VNB_M1004_b N_A_1480_107#_M1013_g 0.0457815f $X=-0.33 $Y=-0.265
+ $X2=2.975 $Y2=0.745
cc_60 N_VNB_M1004_b N_A_1480_107#_M1020_g 0.0497485f $X=-0.33 $Y=-0.265
+ $X2=2.685 $Y2=1.835
cc_61 N_VNB_c_2_p N_A_1480_107#_M1020_g 0.00102867f $X=0.24 $Y=0 $X2=2.685
+ $Y2=1.835
cc_62 N_VNB_M1004_b N_A_1480_107#_c_773_n 0.00953558f $X=-0.33 $Y=-0.265
+ $X2=2.82 $Y2=1.53
cc_63 N_VNB_c_2_p N_A_1480_107#_c_773_n 6.32535e-19 $X=0.24 $Y=0 $X2=2.82
+ $Y2=1.53
cc_64 N_VNB_M1004_b N_A_1480_107#_c_775_n 0.00344775f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_65 N_VNB_M1004_b N_A_1480_107#_c_776_n 0.00378325f $X=-0.33 $Y=-0.265
+ $X2=0.685 $Y2=2.425
cc_66 N_VNB_M1004_b N_A_1480_107#_c_777_n 0.0113523f $X=-0.33 $Y=-0.265
+ $X2=0.685 $Y2=2.625
cc_67 N_VNB_M1004_b N_A_1480_107#_c_778_n 0.00413102f $X=-0.33 $Y=-0.265
+ $X2=0.75 $Y2=2.625
cc_68 N_VNB_M1004_b N_A_1480_107#_c_779_n 6.14009e-19 $X=-0.33 $Y=-0.265
+ $X2=0.75 $Y2=2.61
cc_69 N_VNB_M1004_b N_A_1480_107#_c_780_n 4.83292e-19 $X=-0.33 $Y=-0.265
+ $X2=2.94 $Y2=1.53
cc_70 N_VNB_M1004_b N_A_1480_107#_c_781_n 0.00386664f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_71 N_VNB_M1004_b N_A_1480_107#_c_782_n 0.0993206f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_72 N_VNB_M1004_b N_A_489_107#_c_984_n 0.00889136f $X=-0.33 $Y=-0.265
+ $X2=0.695 $Y2=1.585
cc_73 N_VNB_M1004_b N_A_489_107#_c_985_n 0.00341124f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_74 N_VNB_M1004_b N_A_489_107#_c_986_n 0.0088334f $X=-0.33 $Y=-0.265 $X2=2.82
+ $Y2=1.53
cc_75 N_VNB_M1004_b N_A_489_107#_c_987_n 0.0109104f $X=-0.33 $Y=-0.265 $X2=2.94
+ $Y2=1.53
cc_76 N_VNB_c_2_p N_A_489_107#_c_987_n 8.65969e-19 $X=0.24 $Y=0 $X2=2.94
+ $Y2=1.53
cc_77 N_VNB_M1004_b N_A_489_107#_c_989_n 0.00936525f $X=-0.33 $Y=-0.265 $X2=0.75
+ $Y2=2.305
cc_78 N_VNB_M1004_b N_A_489_107#_c_990_n 0.0106999f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_79 N_VNB_M1004_b N_Q_c_1137_n 0.0634697f $X=-0.33 $Y=-0.265 $X2=2.685
+ $Y2=1.57
cc_80 N_VNB_c_2_p N_Q_c_1137_n 8.4323e-19 $X=0.24 $Y=0 $X2=2.685 $Y2=1.57
cc_81 N_VNB_M1004_b N_VGND_c_1152_n 0.0496364f $X=-0.33 $Y=-0.265 $X2=1.795
+ $Y2=1.92
cc_82 N_VNB_c_2_p N_VGND_c_1152_n 0.00269373f $X=0.24 $Y=0 $X2=1.795 $Y2=1.92
cc_83 N_VNB_M1004_b N_VGND_c_1154_n 0.0326631f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=2.32
cc_84 N_VNB_c_2_p N_VGND_c_1154_n 0.00167165f $X=0.24 $Y=0 $X2=0.635 $Y2=2.32
cc_85 N_VNB_M1004_b N_VGND_c_1156_n 0.0398898f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.27
cc_86 N_VNB_c_2_p N_VGND_c_1156_n 0.00167079f $X=0.24 $Y=0 $X2=0.685 $Y2=2.27
cc_87 N_VNB_M1004_b N_VGND_c_1158_n 0.0593794f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_88 N_VNB_c_2_p N_VGND_c_1158_n 0.00270289f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_89 N_VNB_M1004_b N_VGND_c_1160_n 0.0577136f $X=-0.33 $Y=-0.265 $X2=0.75
+ $Y2=2.305
cc_90 N_VNB_c_2_p N_VGND_c_1160_n 0.00269049f $X=0.24 $Y=0 $X2=0.75 $Y2=2.305
cc_91 N_VNB_M1004_b N_VGND_c_1162_n 0.170998f $X=-0.33 $Y=-0.265 $X2=1.68
+ $Y2=2.305
cc_92 N_VNB_c_2_p N_VGND_c_1162_n 1.23199f $X=0.24 $Y=0 $X2=1.68 $Y2=2.305
cc_93 N_VPB_M1018_b N_SCE_c_218_n 0.0394936f $X=-0.33 $Y=1.885 $X2=1.56
+ $Y2=2.825
cc_94 VPB N_SCE_c_218_n 0.00282611f $X=0 $Y=3.955 $X2=1.56 $Y2=2.825
cc_95 N_VPB_c_95_p N_SCE_c_218_n 0.012804f $X=11.28 $Y=4.07 $X2=1.56 $Y2=2.825
cc_96 N_VPB_M1018_b N_SCE_c_212_n 0.00632721f $X=-0.33 $Y=1.885 $X2=2.6 $Y2=1.92
cc_97 N_VPB_M1018_b N_SCE_c_222_n 0.0396819f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.425
cc_98 VPB N_SCE_c_222_n 4.80548e-19 $X=0 $Y=3.955 $X2=0.685 $Y2=2.425
cc_99 N_VPB_c_95_p N_SCE_c_222_n 0.00338556f $X=11.28 $Y=4.07 $X2=0.685
+ $Y2=2.425
cc_100 N_VPB_M1018_b N_SCE_c_216_n 0.0521971f $X=-0.33 $Y=1.885 $X2=0.75
+ $Y2=2.27
cc_101 N_VPB_M1018_b N_SCE_c_226_n 0.093224f $X=-0.33 $Y=1.885 $X2=1.34 $Y2=2.61
cc_102 N_VPB_M1018_b N_SCE_c_217_n 0.00149264f $X=-0.33 $Y=1.885 $X2=1.795
+ $Y2=2.305
cc_103 N_VPB_M1018_b N_A_30_587#_c_287_n 0.0747542f $X=-0.33 $Y=1.885 $X2=2.975
+ $Y2=0.745
cc_104 N_VPB_c_95_p N_A_30_587#_c_287_n 0.00357885f $X=11.28 $Y=4.07 $X2=2.975
+ $Y2=0.745
cc_105 N_VPB_M1018_b N_A_30_587#_c_296_n 0.0058196f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_106 N_VPB_M1018_b N_A_30_587#_c_297_n 0.120375f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_107 VPB N_A_30_587#_c_297_n 0.00282611f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_108 N_VPB_c_95_p N_A_30_587#_c_297_n 0.0147142f $X=11.28 $Y=4.07 $X2=0 $Y2=0
cc_109 N_VPB_M1018_b N_A_30_587#_c_291_n 3.61802e-19 $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.425
cc_110 N_VPB_M1018_b N_D_M1015_g 0.00660615f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=3.145
cc_111 N_VPB_M1018_b N_D_M1017_g 0.0871796f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_112 VPB N_D_M1017_g 0.00282611f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_113 N_VPB_c_95_p N_D_M1017_g 0.0149809f $X=11.28 $Y=4.07 $X2=0 $Y2=0
cc_114 N_VPB_M1018_b N_D_c_375_n 0.0837085f $X=-0.33 $Y=1.885 $X2=0.695
+ $Y2=1.585
cc_115 N_VPB_M1018_b N_SCD_c_413_n 0.116153f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=1.585
cc_116 VPB N_SCD_c_413_n 0.00282611f $X=0 $Y=3.955 $X2=0.685 $Y2=1.585
cc_117 N_VPB_c_95_p N_SCD_c_413_n 0.00942901f $X=11.28 $Y=4.07 $X2=0.685
+ $Y2=1.585
cc_118 N_VPB_M1018_b N_GATE_c_455_n 0.0697791f $X=-0.33 $Y=1.885 $X2=1.56
+ $Y2=3.31
cc_119 VPB N_GATE_c_455_n 0.00282611f $X=0 $Y=3.955 $X2=1.56 $Y2=3.31
cc_120 N_VPB_c_95_p N_GATE_c_455_n 0.0112134f $X=11.28 $Y=4.07 $X2=1.56 $Y2=3.31
cc_121 N_VPB_M1018_b N_GATE_c_453_n 0.0664792f $X=-0.33 $Y=1.885 $X2=2.685
+ $Y2=1.695
cc_122 N_VPB_M1018_b N_A_1214_107#_c_501_n 0.0602896f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_123 N_VPB_M1018_b N_A_1214_107#_M1000_g 0.0453453f $X=-0.33 $Y=1.885 $X2=1.56
+ $Y2=3.31
cc_124 VPB N_A_1214_107#_M1000_g 0.00196852f $X=0 $Y=3.955 $X2=1.56 $Y2=3.31
cc_125 N_VPB_c_95_p N_A_1214_107#_M1000_g 0.00883031f $X=11.28 $Y=4.07 $X2=1.56
+ $Y2=3.31
cc_126 N_VPB_M1018_b N_A_1214_107#_c_505_n 0.0111669f $X=-0.33 $Y=1.885
+ $X2=1.795 $Y2=1.92
cc_127 N_VPB_M1018_b N_A_1214_107#_c_506_n 0.00347787f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_128 N_VPB_M1018_b N_A_1214_107#_c_507_n 0.00408753f $X=-0.33 $Y=1.885
+ $X2=0.685 $Y2=2.425
cc_129 N_VPB_M1018_b N_A_1214_107#_c_498_n 0.00365362f $X=-0.33 $Y=1.885
+ $X2=0.685 $Y2=2.625
cc_130 N_VPB_M1018_b N_A_944_107#_c_593_n 0.0425912f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_131 VPB N_A_944_107#_c_593_n 4.92992e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_132 N_VPB_c_95_p N_A_944_107#_c_593_n 0.00294781f $X=11.28 $Y=4.07 $X2=0
+ $Y2=0
cc_133 N_VPB_M1018_b N_A_944_107#_c_596_n 0.108865f $X=-0.33 $Y=1.885 $X2=1.56
+ $Y2=3.31
cc_134 N_VPB_M1018_b N_A_944_107#_c_582_n 0.0915199f $X=-0.33 $Y=1.885 $X2=2.975
+ $Y2=0.745
cc_135 N_VPB_M1018_b N_A_944_107#_M1007_g 0.0758064f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_136 VPB N_A_944_107#_M1007_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_137 N_VPB_c_95_p N_A_944_107#_M1007_g 0.0190881f $X=11.28 $Y=4.07 $X2=0 $Y2=0
cc_138 N_VPB_M1018_b N_A_944_107#_c_601_n 0.0696022f $X=-0.33 $Y=1.885 $X2=2.685
+ $Y2=1.835
cc_139 N_VPB_M1018_b N_A_944_107#_c_586_n 0.0240522f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_140 N_VPB_M1018_b N_A_944_107#_M1005_g 0.0143845f $X=-0.33 $Y=1.885 $X2=1.34
+ $Y2=2.625
cc_141 N_VPB_M1018_b N_A_1678_81#_M1001_g 0.126183f $X=-0.33 $Y=1.885 $X2=2.975
+ $Y2=0.745
cc_142 N_VPB_c_95_p N_A_1678_81#_M1001_g 0.0018103f $X=11.28 $Y=4.07 $X2=2.975
+ $Y2=0.745
cc_143 N_VPB_M1018_b N_A_1678_81#_c_702_n 0.00231579f $X=-0.33 $Y=1.885
+ $X2=2.685 $Y2=1.695
cc_144 N_VPB_M1018_b N_A_1678_81#_c_703_n 0.00180874f $X=-0.33 $Y=1.885 $X2=2.82
+ $Y2=1.53
cc_145 N_VPB_M1018_b N_A_1678_81#_c_704_n 0.0128136f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_146 N_VPB_M1018_b N_A_1480_107#_M1011_g 0.0437171f $X=-0.33 $Y=1.885 $X2=1.56
+ $Y2=3.31
cc_147 N_VPB_M1018_b N_A_1480_107#_M1021_g 0.0424813f $X=-0.33 $Y=1.885
+ $X2=0.695 $Y2=1.585
cc_148 VPB N_A_1480_107#_M1021_g 0.00970178f $X=0 $Y=3.955 $X2=0.695 $Y2=1.585
cc_149 N_VPB_c_95_p N_A_1480_107#_M1021_g 0.0162989f $X=11.28 $Y=4.07 $X2=0.695
+ $Y2=1.585
cc_150 N_VPB_M1018_b N_A_1480_107#_c_787_n 0.00803094f $X=-0.33 $Y=1.885
+ $X2=1.115 $Y2=2.32
cc_151 N_VPB_M1018_b N_A_1480_107#_c_788_n 0.00539731f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_152 VPB N_A_1480_107#_c_788_n 0.00104693f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_153 N_VPB_c_95_p N_A_1480_107#_c_788_n 0.0172373f $X=11.28 $Y=4.07 $X2=0
+ $Y2=0
cc_154 N_VPB_M1018_b N_A_1480_107#_c_791_n 0.00928095f $X=-0.33 $Y=1.885
+ $X2=0.685 $Y2=2.27
cc_155 N_VPB_M1018_b N_A_1480_107#_c_778_n 0.00499514f $X=-0.33 $Y=1.885
+ $X2=0.75 $Y2=2.625
cc_156 N_VPB_M1018_b N_A_1480_107#_c_779_n 0.00264604f $X=-0.33 $Y=1.885
+ $X2=0.75 $Y2=2.61
cc_157 N_VPB_M1018_b N_A_1480_107#_c_794_n 0.00992348f $X=-0.33 $Y=1.885
+ $X2=1.34 $Y2=2.625
cc_158 N_VPB_M1018_b N_A_1480_107#_c_781_n 0.00476546f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_159 N_VPB_M1018_b N_A_1480_107#_c_782_n 0.0453947f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_160 N_VPB_M1018_b N_VPWR_c_893_n 0.007562f $X=-0.33 $Y=1.885 $X2=1.795
+ $Y2=1.92
cc_161 VPB N_VPWR_c_893_n 0.00307235f $X=0 $Y=3.955 $X2=1.795 $Y2=1.92
cc_162 N_VPB_c_95_p N_VPWR_c_893_n 0.0402284f $X=11.28 $Y=4.07 $X2=1.795
+ $Y2=1.92
cc_163 N_VPB_M1018_b N_VPWR_c_896_n 0.00243384f $X=-0.33 $Y=1.885 $X2=0.75
+ $Y2=2.27
cc_164 VPB N_VPWR_c_896_n 0.00375116f $X=0 $Y=3.955 $X2=0.75 $Y2=2.27
cc_165 N_VPB_c_95_p N_VPWR_c_896_n 0.0420982f $X=11.28 $Y=4.07 $X2=0.75 $Y2=2.27
cc_166 N_VPB_M1018_b N_VPWR_c_899_n 0.0078136f $X=-0.33 $Y=1.885 $X2=0.75
+ $Y2=2.61
cc_167 VPB N_VPWR_c_899_n 4.76796e-19 $X=0 $Y=3.955 $X2=0.75 $Y2=2.61
cc_168 N_VPB_c_95_p N_VPWR_c_899_n 0.00726526f $X=11.28 $Y=4.07 $X2=0.75
+ $Y2=2.61
cc_169 N_VPB_M1018_b N_VPWR_c_902_n 0.0151561f $X=-0.33 $Y=1.885 $X2=2.94
+ $Y2=1.085
cc_170 VPB N_VPWR_c_902_n 0.00268927f $X=0 $Y=3.955 $X2=2.94 $Y2=1.085
cc_171 N_VPB_c_95_p N_VPWR_c_902_n 0.0410163f $X=11.28 $Y=4.07 $X2=2.94
+ $Y2=1.085
cc_172 N_VPB_M1018_b N_VPWR_c_905_n 0.0239961f $X=-0.33 $Y=1.885 $X2=1.68
+ $Y2=2.305
cc_173 VPB N_VPWR_c_905_n 0.00335473f $X=0 $Y=3.955 $X2=1.68 $Y2=2.305
cc_174 N_VPB_c_95_p N_VPWR_c_905_n 0.0490696f $X=11.28 $Y=4.07 $X2=1.68
+ $Y2=2.305
cc_175 N_VPB_M1018_b N_VPWR_c_908_n 0.125921f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_908_n 1.22607f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_177 N_VPB_c_95_p N_VPWR_c_908_n 0.0576181f $X=11.28 $Y=4.07 $X2=0 $Y2=0
cc_178 N_VPB_M1018_b N_A_489_107#_c_991_n 0.00236203f $X=-0.33 $Y=1.885
+ $X2=0.685 $Y2=1.585
cc_179 VPB N_A_489_107#_c_991_n 7.69934e-19 $X=0 $Y=3.955 $X2=0.685 $Y2=1.585
cc_180 N_VPB_c_95_p N_A_489_107#_c_991_n 0.0114811f $X=11.28 $Y=4.07 $X2=0.685
+ $Y2=1.585
cc_181 N_VPB_M1018_b N_A_489_107#_c_994_n 0.00960226f $X=-0.33 $Y=1.885
+ $X2=1.795 $Y2=1.92
cc_182 N_VPB_M1018_b N_A_489_107#_c_995_n 0.00595173f $X=-0.33 $Y=1.885
+ $X2=2.685 $Y2=1.695
cc_183 N_VPB_M1018_b N_A_489_107#_c_986_n 0.0137518f $X=-0.33 $Y=1.885 $X2=2.82
+ $Y2=1.53
cc_184 N_VPB_M1018_b N_A_489_107#_c_997_n 0.0014452f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_185 N_VPB_M1018_b N_A_489_107#_c_998_n 0.00710874f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_186 VPB N_A_489_107#_c_998_n 0.00248257f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_187 N_VPB_c_95_p N_A_489_107#_c_998_n 0.0459346f $X=11.28 $Y=4.07 $X2=0 $Y2=0
cc_188 VPB N_A_489_107#_c_1001_n 8.17382e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_189 N_VPB_c_95_p N_A_489_107#_c_1001_n 0.0107872f $X=11.28 $Y=4.07 $X2=0
+ $Y2=0
cc_190 N_VPB_M1018_b N_A_489_107#_c_1003_n 0.0244999f $X=-0.33 $Y=1.885
+ $X2=0.685 $Y2=2.425
cc_191 N_VPB_M1018_b N_A_489_107#_c_1004_n 0.0135652f $X=-0.33 $Y=1.885
+ $X2=0.685 $Y2=2.27
cc_192 N_VPB_M1018_b N_A_489_107#_c_1005_n 0.00919848f $X=-0.33 $Y=1.885
+ $X2=0.75 $Y2=2.27
cc_193 N_VPB_M1018_b N_A_489_107#_c_1006_n 0.00145965f $X=-0.33 $Y=1.885
+ $X2=0.685 $Y2=2.625
cc_194 N_VPB_M1018_b N_A_489_107#_c_1007_n 0.0157969f $X=-0.33 $Y=1.885 $X2=0.75
+ $Y2=2.625
cc_195 VPB N_A_489_107#_c_1007_n 0.0037738f $X=0 $Y=3.955 $X2=0.75 $Y2=2.625
cc_196 N_VPB_c_95_p N_A_489_107#_c_1007_n 0.064276f $X=11.28 $Y=4.07 $X2=0.75
+ $Y2=2.625
cc_197 N_VPB_M1018_b N_A_489_107#_c_1010_n 0.00210815f $X=-0.33 $Y=1.885
+ $X2=0.75 $Y2=2.61
cc_198 VPB N_A_489_107#_c_1010_n 5.37289e-19 $X=0 $Y=3.955 $X2=0.75 $Y2=2.61
cc_199 N_VPB_c_95_p N_A_489_107#_c_1010_n 0.00939255f $X=11.28 $Y=4.07 $X2=0.75
+ $Y2=2.61
cc_200 N_VPB_M1018_b N_A_489_107#_c_1013_n 0.00700687f $X=-0.33 $Y=1.885
+ $X2=1.34 $Y2=2.61
cc_201 N_VPB_M1018_b N_A_489_107#_c_1014_n 0.00152933f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_202 N_VPB_M1018_b N_A_489_107#_c_1015_n 0.0102605f $X=-0.33 $Y=1.885 $X2=1.68
+ $Y2=2.305
cc_203 N_VPB_M1018_b N_A_489_107#_c_990_n 0.0119876f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_204 N_VPB_M1018_b N_Q_c_1137_n 0.0670661f $X=-0.33 $Y=1.885 $X2=2.685
+ $Y2=1.57
cc_205 VPB N_Q_c_1137_n 0.00107758f $X=0 $Y=3.955 $X2=2.685 $Y2=1.57
cc_206 N_VPB_c_95_p N_Q_c_1137_n 0.0177658f $X=11.28 $Y=4.07 $X2=2.685 $Y2=1.57
cc_207 N_SCE_M1004_g N_A_30_587#_c_285_n 0.0159945f $X=0.705 $Y=0.745 $X2=0
+ $Y2=0
cc_208 N_SCE_c_211_n N_A_30_587#_c_285_n 0.00664239f $X=0.695 $Y=1.585 $X2=0
+ $Y2=0
cc_209 N_SCE_c_211_n N_A_30_587#_c_287_n 0.0601516f $X=0.695 $Y=1.585 $X2=0
+ $Y2=0
cc_210 N_SCE_c_217_n N_A_30_587#_c_287_n 0.0668666f $X=1.795 $Y=2.305 $X2=0
+ $Y2=0
cc_211 N_SCE_c_211_n N_A_30_587#_c_288_n 0.0313291f $X=0.695 $Y=1.585 $X2=0
+ $Y2=0
cc_212 N_SCE_c_217_n N_A_30_587#_c_288_n 0.0477546f $X=1.795 $Y=2.305 $X2=0
+ $Y2=0
cc_213 N_SCE_c_212_n N_A_30_587#_c_289_n 0.00930681f $X=2.6 $Y=1.92 $X2=11.28
+ $Y2=0
cc_214 N_SCE_c_214_n N_A_30_587#_c_289_n 0.0261157f $X=2.82 $Y=1.53 $X2=11.28
+ $Y2=0
cc_215 N_SCE_c_215_n N_A_30_587#_c_289_n 0.0273928f $X=2.82 $Y=1.53 $X2=11.28
+ $Y2=0
cc_216 N_SCE_c_211_n N_A_30_587#_c_290_n 0.00643921f $X=0.695 $Y=1.585 $X2=5.76
+ $Y2=0.057
cc_217 N_SCE_c_212_n N_A_30_587#_c_311_n 0.0247098f $X=2.6 $Y=1.92 $X2=5.76
+ $Y2=0.058
cc_218 N_SCE_c_214_n N_A_30_587#_c_311_n 0.0108722f $X=2.82 $Y=1.53 $X2=5.76
+ $Y2=0.058
cc_219 N_SCE_c_215_n N_A_30_587#_c_311_n 0.00124261f $X=2.82 $Y=1.53 $X2=5.76
+ $Y2=0.058
cc_220 N_SCE_c_212_n N_A_30_587#_c_296_n 0.00816237f $X=2.6 $Y=1.92 $X2=0 $Y2=0
cc_221 N_SCE_c_214_n N_A_30_587#_c_296_n 0.00221894f $X=2.82 $Y=1.53 $X2=0 $Y2=0
cc_222 N_SCE_c_215_n N_A_30_587#_c_296_n 0.00104415f $X=2.82 $Y=1.53 $X2=0 $Y2=0
cc_223 N_SCE_c_212_n N_A_30_587#_c_297_n 0.00201857f $X=2.6 $Y=1.92 $X2=0 $Y2=0
cc_224 N_SCE_c_214_n N_A_30_587#_c_297_n 0.00120844f $X=2.82 $Y=1.53 $X2=0 $Y2=0
cc_225 N_SCE_c_215_n N_A_30_587#_c_297_n 0.0297566f $X=2.82 $Y=1.53 $X2=0 $Y2=0
cc_226 N_SCE_c_212_n N_A_30_587#_c_291_n 0.00327323f $X=2.6 $Y=1.92 $X2=0 $Y2=0
cc_227 N_SCE_c_213_n N_A_30_587#_c_291_n 0.00586729f $X=2.685 $Y=1.835 $X2=0
+ $Y2=0
cc_228 N_SCE_c_214_n N_A_30_587#_c_291_n 0.0172129f $X=2.82 $Y=1.53 $X2=0 $Y2=0
cc_229 N_SCE_c_215_n N_A_30_587#_c_291_n 0.0161209f $X=2.82 $Y=1.53 $X2=0 $Y2=0
cc_230 N_SCE_M1008_g N_A_30_587#_M1016_g 0.0160132f $X=2.975 $Y=0.745 $X2=0
+ $Y2=0
cc_231 N_SCE_c_212_n N_A_30_587#_M1016_g 0.00431326f $X=2.6 $Y=1.92 $X2=0 $Y2=0
cc_232 N_SCE_c_213_n N_A_30_587#_M1016_g 0.00201124f $X=2.685 $Y=1.835 $X2=0
+ $Y2=0
cc_233 N_SCE_c_214_n N_A_30_587#_M1016_g 0.00266436f $X=2.82 $Y=1.53 $X2=0 $Y2=0
cc_234 N_SCE_c_215_n N_A_30_587#_M1016_g 0.0414695f $X=2.82 $Y=1.53 $X2=0 $Y2=0
cc_235 N_SCE_M1004_g N_D_M1015_g 0.0425237f $X=0.705 $Y=0.745 $X2=0 $Y2=0
cc_236 N_SCE_c_216_n N_D_M1015_g 0.0301591f $X=0.75 $Y=2.27 $X2=0 $Y2=0
cc_237 N_SCE_c_217_n N_D_M1015_g 0.0230251f $X=1.795 $Y=2.305 $X2=0 $Y2=0
cc_238 N_SCE_c_226_n N_D_M1017_g 0.0948437f $X=1.34 $Y=2.61 $X2=0 $Y2=0
cc_239 N_SCE_c_217_n N_D_M1017_g 0.00521373f $X=1.795 $Y=2.305 $X2=0 $Y2=0
cc_240 N_SCE_c_212_n N_D_c_375_n 0.0307893f $X=2.6 $Y=1.92 $X2=11.28 $Y2=0
cc_241 N_SCE_c_226_n N_D_c_375_n 0.0336088f $X=1.34 $Y=2.61 $X2=11.28 $Y2=0
cc_242 N_SCE_c_217_n N_D_c_375_n 0.0369845f $X=1.795 $Y=2.305 $X2=11.28 $Y2=0
cc_243 N_SCE_c_212_n N_D_c_384_n 0.0238596f $X=2.6 $Y=1.92 $X2=0 $Y2=0
cc_244 N_SCE_c_226_n N_D_c_384_n 0.00388085f $X=1.34 $Y=2.61 $X2=0 $Y2=0
cc_245 N_SCE_c_217_n N_D_c_384_n 0.0360125f $X=1.795 $Y=2.305 $X2=0 $Y2=0
cc_246 N_SCE_M1008_g N_SCD_M1009_g 0.0403136f $X=2.975 $Y=0.745 $X2=0 $Y2=0
cc_247 N_SCE_c_215_n N_SCD_c_412_n 0.0403136f $X=2.82 $Y=1.53 $X2=0 $Y2=0
cc_248 N_SCE_c_215_n N_SCD_c_413_n 0.0047642f $X=2.82 $Y=1.53 $X2=0 $Y2=0
cc_249 N_SCE_c_218_n N_VPWR_c_893_n 0.033628f $X=1.56 $Y=2.825 $X2=0 $Y2=0
cc_250 N_SCE_c_222_n N_VPWR_c_893_n 0.0452269f $X=0.685 $Y=2.425 $X2=0 $Y2=0
cc_251 N_SCE_c_226_n N_VPWR_c_893_n 0.00487654f $X=1.34 $Y=2.61 $X2=0 $Y2=0
cc_252 N_SCE_c_217_n N_VPWR_c_893_n 0.0602571f $X=1.795 $Y=2.305 $X2=0 $Y2=0
cc_253 N_SCE_c_218_n N_VPWR_c_908_n 0.0206647f $X=1.56 $Y=2.825 $X2=0 $Y2=0
cc_254 N_SCE_c_222_n N_VPWR_c_908_n 0.0078567f $X=0.685 $Y=2.425 $X2=0 $Y2=0
cc_255 N_SCE_M1008_g N_A_489_107#_c_984_n 0.0260633f $X=2.975 $Y=0.745 $X2=11.28
+ $Y2=0
cc_256 N_SCE_c_212_n N_A_489_107#_c_995_n 0.00653246f $X=2.6 $Y=1.92 $X2=0 $Y2=0
cc_257 N_SCE_M1008_g N_A_489_107#_c_1019_n 0.0011108f $X=2.975 $Y=0.745 $X2=0
+ $Y2=0
cc_258 N_SCE_M1008_g N_A_489_107#_c_987_n 0.00825293f $X=2.975 $Y=0.745 $X2=0
+ $Y2=0
cc_259 N_SCE_c_215_n N_A_489_107#_c_987_n 0.00166757f $X=2.82 $Y=1.53 $X2=0
+ $Y2=0
cc_260 N_SCE_M1004_g N_VGND_c_1152_n 0.0358184f $X=0.705 $Y=0.745 $X2=0 $Y2=0
cc_261 N_SCE_M1008_g N_VGND_c_1154_n 0.00158455f $X=2.975 $Y=0.745 $X2=0 $Y2=0
cc_262 N_SCE_M1004_g N_VGND_c_1162_n 0.00618666f $X=0.705 $Y=0.745 $X2=0 $Y2=0
cc_263 N_SCE_M1008_g N_VGND_c_1162_n 0.0151022f $X=2.975 $Y=0.745 $X2=0 $Y2=0
cc_264 N_A_30_587#_c_288_n N_D_M1015_g 0.0318386f $X=1.965 $Y=1.26 $X2=0 $Y2=0
cc_265 N_A_30_587#_c_311_n N_D_M1015_g 0.00286609f $X=2.13 $Y=1.18 $X2=0 $Y2=0
cc_266 N_A_30_587#_M1016_g N_D_M1015_g 0.0966721f $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_267 N_A_30_587#_c_296_n N_D_M1017_g 0.00105308f $X=3.115 $Y=2.07 $X2=0 $Y2=0
cc_268 N_A_30_587#_c_288_n N_D_c_375_n 9.69651e-19 $X=1.965 $Y=1.26 $X2=11.28
+ $Y2=0
cc_269 N_A_30_587#_c_289_n N_D_c_375_n 4.11296e-19 $X=3.165 $Y=1.18 $X2=11.28
+ $Y2=0
cc_270 N_A_30_587#_c_311_n N_D_c_375_n 2.8044e-19 $X=2.13 $Y=1.18 $X2=11.28
+ $Y2=0
cc_271 N_A_30_587#_c_296_n N_D_c_375_n 0.00108666f $X=3.115 $Y=2.07 $X2=11.28
+ $Y2=0
cc_272 N_A_30_587#_c_297_n N_D_c_375_n 0.0604181f $X=3.115 $Y=2.07 $X2=11.28
+ $Y2=0
cc_273 N_A_30_587#_M1016_g N_D_c_375_n 0.0329045f $X=2.195 $Y=0.745 $X2=11.28
+ $Y2=0
cc_274 N_A_30_587#_c_296_n N_D_c_384_n 0.00853905f $X=3.115 $Y=2.07 $X2=0 $Y2=0
cc_275 N_A_30_587#_c_297_n N_D_c_384_n 0.00233979f $X=3.115 $Y=2.07 $X2=0 $Y2=0
cc_276 N_A_30_587#_c_289_n N_SCD_c_412_n 0.00131336f $X=3.165 $Y=1.18 $X2=0
+ $Y2=0
cc_277 N_A_30_587#_c_291_n N_SCD_c_412_n 0.00502504f $X=3.142 $Y=1.905 $X2=0
+ $Y2=0
cc_278 N_A_30_587#_c_297_n SCD 6.82618e-19 $X=3.115 $Y=2.07 $X2=0 $Y2=0
cc_279 N_A_30_587#_c_291_n SCD 0.072765f $X=3.142 $Y=1.905 $X2=0 $Y2=0
cc_280 N_A_30_587#_c_297_n N_SCD_c_413_n 0.129804f $X=3.115 $Y=2.07 $X2=0 $Y2=0
cc_281 N_A_30_587#_c_291_n N_SCD_c_413_n 0.00946251f $X=3.142 $Y=1.905 $X2=0
+ $Y2=0
cc_282 N_A_30_587#_c_287_n N_VPWR_c_893_n 0.017513f $X=0.295 $Y=3.145 $X2=0
+ $Y2=0
cc_283 N_A_30_587#_c_297_n N_VPWR_c_896_n 0.00901155f $X=3.115 $Y=2.07 $X2=0
+ $Y2=0
cc_284 N_A_30_587#_c_287_n N_VPWR_c_908_n 0.0110536f $X=0.295 $Y=3.145 $X2=0
+ $Y2=0
cc_285 N_A_30_587#_c_297_n N_VPWR_c_908_n 0.0157473f $X=3.115 $Y=2.07 $X2=0
+ $Y2=0
cc_286 N_A_30_587#_c_297_n N_A_489_107#_c_991_n 0.0221785f $X=3.115 $Y=2.07
+ $X2=0 $Y2=0
cc_287 N_A_30_587#_c_289_n N_A_489_107#_c_984_n 0.0361079f $X=3.165 $Y=1.18
+ $X2=11.28 $Y2=0
cc_288 N_A_30_587#_c_296_n N_A_489_107#_c_994_n 0.0279607f $X=3.115 $Y=2.07
+ $X2=0 $Y2=0
cc_289 N_A_30_587#_c_297_n N_A_489_107#_c_994_n 0.0309179f $X=3.115 $Y=2.07
+ $X2=0 $Y2=0
cc_290 N_A_30_587#_c_297_n N_A_489_107#_c_995_n 0.00324065f $X=3.115 $Y=2.07
+ $X2=0 $Y2=0
cc_291 N_A_30_587#_c_289_n N_A_489_107#_c_1019_n 0.00615029f $X=3.165 $Y=1.18
+ $X2=0 $Y2=0
cc_292 N_A_30_587#_c_289_n N_A_489_107#_c_1028_n 0.00768578f $X=3.165 $Y=1.18
+ $X2=5.76 $Y2=0.058
cc_293 N_A_30_587#_c_291_n N_A_489_107#_c_1028_n 0.00608785f $X=3.142 $Y=1.905
+ $X2=5.76 $Y2=0.058
cc_294 N_A_30_587#_c_289_n N_A_489_107#_c_987_n 0.018802f $X=3.165 $Y=1.18 $X2=0
+ $Y2=0
cc_295 N_A_30_587#_M1016_g N_A_489_107#_c_987_n 0.011462f $X=2.195 $Y=0.745
+ $X2=0 $Y2=0
cc_296 N_A_30_587#_c_285_n N_VGND_c_1152_n 0.0361847f $X=0.315 $Y=0.745 $X2=0
+ $Y2=0
cc_297 N_A_30_587#_c_288_n N_VGND_c_1152_n 0.0686854f $X=1.965 $Y=1.26 $X2=0
+ $Y2=0
cc_298 N_A_30_587#_M1016_g N_VGND_c_1152_n 0.00407355f $X=2.195 $Y=0.745 $X2=0
+ $Y2=0
cc_299 N_A_30_587#_c_285_n N_VGND_c_1162_n 0.0344602f $X=0.315 $Y=0.745 $X2=0
+ $Y2=0
cc_300 N_A_30_587#_c_288_n N_VGND_c_1162_n 0.0195359f $X=1.965 $Y=1.26 $X2=0
+ $Y2=0
cc_301 N_A_30_587#_c_289_n N_VGND_c_1162_n 0.00571924f $X=3.165 $Y=1.18 $X2=0
+ $Y2=0
cc_302 N_A_30_587#_c_311_n N_VGND_c_1162_n 0.0112852f $X=2.13 $Y=1.18 $X2=0
+ $Y2=0
cc_303 N_A_30_587#_M1016_g N_VGND_c_1162_n 0.0173471f $X=2.195 $Y=0.745 $X2=0
+ $Y2=0
cc_304 N_D_M1017_g N_VPWR_c_893_n 0.00309089f $X=2.27 $Y=3.31 $X2=0 $Y2=0
cc_305 N_D_c_384_n N_VPWR_c_893_n 0.00829215f $X=2.205 $Y=2.27 $X2=0 $Y2=0
cc_306 N_D_M1017_g N_VPWR_c_908_n 0.0211812f $X=2.27 $Y=3.31 $X2=0 $Y2=0
cc_307 N_D_c_384_n N_VPWR_c_908_n 0.0158931f $X=2.205 $Y=2.27 $X2=0 $Y2=0
cc_308 N_D_M1017_g N_A_489_107#_c_991_n 0.00438833f $X=2.27 $Y=3.31 $X2=0 $Y2=0
cc_309 N_D_c_384_n N_A_489_107#_c_991_n 0.0164829f $X=2.205 $Y=2.27 $X2=0 $Y2=0
cc_310 N_D_M1017_g N_A_489_107#_c_995_n 0.00172221f $X=2.27 $Y=3.31 $X2=0 $Y2=0
cc_311 N_D_c_384_n N_A_489_107#_c_995_n 0.0124553f $X=2.205 $Y=2.27 $X2=0 $Y2=0
cc_312 N_D_M1015_g N_A_489_107#_c_987_n 0.0014684f $X=1.485 $Y=0.745 $X2=0 $Y2=0
cc_313 N_D_M1015_g N_VGND_c_1152_n 0.0445503f $X=1.485 $Y=0.745 $X2=0 $Y2=0
cc_314 N_D_M1015_g N_VGND_c_1162_n 0.00461913f $X=1.485 $Y=0.745 $X2=0 $Y2=0
cc_315 N_SCD_M1009_g N_GATE_M1006_g 0.0140267f $X=3.685 $Y=0.745 $X2=0 $Y2=0
cc_316 N_SCD_c_413_n N_GATE_c_455_n 0.0151736f $X=3.695 $Y=1.69 $X2=0 $Y2=0
cc_317 N_SCD_c_412_n GATE 6.55407e-19 $X=3.722 $Y=1.585 $X2=0.24 $Y2=0
cc_318 N_SCD_c_413_n N_GATE_c_453_n 0.0555728f $X=3.695 $Y=1.69 $X2=0 $Y2=0
cc_319 N_SCD_c_412_n N_GATE_c_454_n 0.0555728f $X=3.722 $Y=1.585 $X2=5.76
+ $Y2=0.057
cc_320 N_SCD_c_413_n N_VPWR_c_896_n 0.0478675f $X=3.695 $Y=1.69 $X2=0 $Y2=0
cc_321 N_SCD_c_413_n N_VPWR_c_908_n 0.00103564f $X=3.695 $Y=1.69 $X2=0 $Y2=0
cc_322 N_SCD_c_413_n N_A_489_107#_c_991_n 0.00110691f $X=3.695 $Y=1.69 $X2=0
+ $Y2=0
cc_323 N_SCD_M1009_g N_A_489_107#_c_984_n 0.0162966f $X=3.685 $Y=0.745 $X2=11.28
+ $Y2=0
cc_324 SCD N_A_489_107#_c_994_n 0.0249507f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_325 N_SCD_c_413_n N_A_489_107#_c_994_n 0.0298224f $X=3.695 $Y=1.69 $X2=0
+ $Y2=0
cc_326 N_SCD_M1009_g N_A_489_107#_c_1019_n 0.00756837f $X=3.685 $Y=0.745 $X2=0
+ $Y2=0
cc_327 N_SCD_c_412_n N_A_489_107#_c_1019_n 0.00364997f $X=3.722 $Y=1.585 $X2=0
+ $Y2=0
cc_328 N_SCD_c_412_n N_A_489_107#_c_985_n 0.0211472f $X=3.722 $Y=1.585 $X2=5.76
+ $Y2=0.057
cc_329 SCD N_A_489_107#_c_985_n 0.0126247f $X=3.515 $Y=1.58 $X2=5.76 $Y2=0.057
cc_330 N_SCD_c_412_n N_A_489_107#_c_1028_n 0.00636132f $X=3.722 $Y=1.585
+ $X2=5.76 $Y2=0.058
cc_331 SCD N_A_489_107#_c_1028_n 0.013489f $X=3.515 $Y=1.58 $X2=5.76 $Y2=0.058
cc_332 N_SCD_c_412_n N_A_489_107#_c_986_n 0.0163822f $X=3.722 $Y=1.585 $X2=0
+ $Y2=0
cc_333 SCD N_A_489_107#_c_986_n 0.0731014f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_334 N_SCD_c_413_n N_A_489_107#_c_1049_n 8.7508e-19 $X=3.695 $Y=1.69 $X2=0
+ $Y2=0
cc_335 N_SCD_c_413_n N_A_489_107#_c_1001_n 6.53242e-19 $X=3.695 $Y=1.69 $X2=0
+ $Y2=0
cc_336 N_SCD_M1009_g N_A_489_107#_c_987_n 9.82117e-19 $X=3.685 $Y=0.745 $X2=0
+ $Y2=0
cc_337 N_SCD_M1009_g N_VGND_c_1154_n 0.018911f $X=3.685 $Y=0.745 $X2=0 $Y2=0
cc_338 N_SCD_c_412_n N_VGND_c_1154_n 0.00222517f $X=3.722 $Y=1.585 $X2=0 $Y2=0
cc_339 N_SCD_M1009_g N_VGND_c_1162_n 0.0140288f $X=3.685 $Y=0.745 $X2=0 $Y2=0
cc_340 N_GATE_M1006_g N_A_944_107#_c_585_n 0.00452969f $X=4.47 $Y=0.745 $X2=5.76
+ $Y2=0.058
cc_341 GATE N_A_944_107#_c_585_n 0.00210485f $X=4.475 $Y=1.21 $X2=5.76 $Y2=0.058
cc_342 N_GATE_c_454_n N_A_944_107#_c_585_n 0.00360198f $X=4.52 $Y=1.31 $X2=5.76
+ $Y2=0.058
cc_343 GATE N_A_944_107#_c_586_n 0.0819998f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_344 N_GATE_c_454_n N_A_944_107#_c_586_n 0.0500296f $X=4.52 $Y=1.31 $X2=0
+ $Y2=0
cc_345 N_GATE_M1006_g N_A_944_107#_c_588_n 0.0109008f $X=4.47 $Y=0.745 $X2=0
+ $Y2=0
cc_346 N_GATE_c_454_n N_A_944_107#_c_588_n 0.00343943f $X=4.52 $Y=1.31 $X2=0
+ $Y2=0
cc_347 GATE N_A_944_107#_c_590_n 0.013626f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_348 N_GATE_c_454_n N_A_944_107#_c_590_n 0.00511205f $X=4.52 $Y=1.31 $X2=0
+ $Y2=0
cc_349 N_GATE_c_455_n N_VPWR_c_896_n 0.0120389f $X=4.505 $Y=2.825 $X2=0 $Y2=0
cc_350 N_GATE_c_455_n N_VPWR_c_908_n 0.0124669f $X=4.505 $Y=2.825 $X2=0 $Y2=0
cc_351 N_GATE_M1006_g N_A_489_107#_c_1019_n 8.69805e-19 $X=4.47 $Y=0.745 $X2=0
+ $Y2=0
cc_352 GATE N_A_489_107#_c_985_n 0.0142339f $X=4.475 $Y=1.21 $X2=5.76 $Y2=0.057
cc_353 N_GATE_c_454_n N_A_489_107#_c_985_n 0.00150857f $X=4.52 $Y=1.31 $X2=5.76
+ $Y2=0.057
cc_354 GATE N_A_489_107#_c_986_n 0.0856077f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_355 N_GATE_c_454_n N_A_489_107#_c_986_n 0.0113919f $X=4.52 $Y=1.31 $X2=0
+ $Y2=0
cc_356 N_GATE_c_455_n N_A_489_107#_c_997_n 0.0265372f $X=4.505 $Y=2.825 $X2=0
+ $Y2=0
cc_357 GATE N_A_489_107#_c_997_n 0.0226451f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_358 N_GATE_c_455_n N_A_489_107#_c_1049_n 0.029741f $X=4.505 $Y=2.825 $X2=0
+ $Y2=0
cc_359 N_GATE_c_455_n N_A_489_107#_c_998_n 0.00894016f $X=4.505 $Y=2.825 $X2=0
+ $Y2=0
cc_360 N_GATE_c_455_n N_A_489_107#_c_1001_n 0.00523064f $X=4.505 $Y=2.825 $X2=0
+ $Y2=0
cc_361 N_GATE_c_455_n N_A_489_107#_c_1003_n 0.00387557f $X=4.505 $Y=2.825 $X2=0
+ $Y2=0
cc_362 N_GATE_M1006_g N_VGND_c_1154_n 0.0366571f $X=4.47 $Y=0.745 $X2=0 $Y2=0
cc_363 GATE N_VGND_c_1154_n 0.00674369f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_364 N_GATE_M1006_g N_VGND_c_1156_n 0.00285804f $X=4.47 $Y=0.745 $X2=0 $Y2=0
cc_365 N_GATE_M1006_g N_VGND_c_1162_n 0.00966044f $X=4.47 $Y=0.745 $X2=0 $Y2=0
cc_366 GATE N_VGND_c_1162_n 0.00731361f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_367 N_A_1214_107#_c_505_n N_A_944_107#_c_593_n 0.0178141f $X=6.41 $Y=2.75
+ $X2=0 $Y2=0
cc_368 N_A_1214_107#_c_498_n N_A_944_107#_c_593_n 0.00228416f $X=6.41 $Y=2.585
+ $X2=0 $Y2=0
cc_369 N_A_1214_107#_c_505_n N_A_944_107#_c_596_n 0.0082365f $X=6.41 $Y=2.75
+ $X2=0.24 $Y2=0
cc_370 N_A_1214_107#_c_512_p N_A_944_107#_c_596_n 8.4955e-19 $X=7.275 $Y=1.67
+ $X2=0.24 $Y2=0
cc_371 N_A_1214_107#_c_498_n N_A_944_107#_c_596_n 0.0216459f $X=6.41 $Y=2.585
+ $X2=0.24 $Y2=0
cc_372 N_A_1214_107#_M1002_g N_A_944_107#_c_596_n 0.0222601f $X=7.15 $Y=0.745
+ $X2=0.24 $Y2=0
cc_373 N_A_1214_107#_c_501_n N_A_944_107#_c_582_n 0.013819f $X=8.37 $Y=2.775
+ $X2=0 $Y2=0
cc_374 N_A_1214_107#_c_516_p N_A_944_107#_c_582_n 7.42695e-19 $X=7.19 $Y=1.25
+ $X2=0 $Y2=0
cc_375 N_A_1214_107#_c_496_n N_A_944_107#_c_582_n 0.0361045f $X=7.84 $Y=1.67
+ $X2=0 $Y2=0
cc_376 N_A_1214_107#_c_512_p N_A_944_107#_c_582_n 3.63082e-19 $X=7.275 $Y=1.67
+ $X2=0 $Y2=0
cc_377 N_A_1214_107#_c_519_p N_A_944_107#_c_582_n 0.0353296f $X=7.925 $Y=2.215
+ $X2=0 $Y2=0
cc_378 N_A_1214_107#_c_506_n N_A_944_107#_c_582_n 0.016194f $X=8.01 $Y=2.345
+ $X2=0 $Y2=0
cc_379 N_A_1214_107#_c_507_n N_A_944_107#_c_582_n 0.00592006f $X=8.405 $Y=2.38
+ $X2=0 $Y2=0
cc_380 N_A_1214_107#_M1002_g N_A_944_107#_c_582_n 0.0355809f $X=7.15 $Y=0.745
+ $X2=0 $Y2=0
cc_381 N_A_1214_107#_c_501_n N_A_944_107#_M1007_g 0.0229191f $X=8.37 $Y=2.775
+ $X2=0 $Y2=0
cc_382 N_A_1214_107#_c_505_n N_A_944_107#_M1007_g 8.24241e-19 $X=6.41 $Y=2.75
+ $X2=0 $Y2=0
cc_383 N_A_1214_107#_c_492_n N_A_944_107#_M1019_g 2.52933e-19 $X=7.105 $Y=0.35
+ $X2=0 $Y2=0
cc_384 N_A_1214_107#_c_516_p N_A_944_107#_M1019_g 0.00205622f $X=7.19 $Y=1.25
+ $X2=0 $Y2=0
cc_385 N_A_1214_107#_M1002_g N_A_944_107#_M1019_g 0.032203f $X=7.15 $Y=0.745
+ $X2=0 $Y2=0
cc_386 N_A_1214_107#_c_498_n N_A_944_107#_c_601_n 0.0150874f $X=6.41 $Y=2.585
+ $X2=5.76 $Y2=0
cc_387 N_A_1214_107#_c_498_n N_A_944_107#_c_633_n 0.0314765f $X=6.41 $Y=2.585
+ $X2=0 $Y2=0
cc_388 N_A_1214_107#_c_491_n N_A_944_107#_M1005_g 0.00805751f $X=6.21 $Y=0.745
+ $X2=0 $Y2=0
cc_389 N_A_1214_107#_c_494_n N_A_944_107#_M1005_g 0.00157105f $X=6.415 $Y=0.35
+ $X2=0 $Y2=0
cc_390 N_A_1214_107#_c_497_n N_A_944_107#_M1005_g 0.00560284f $X=6.23 $Y=0.975
+ $X2=0 $Y2=0
cc_391 N_A_1214_107#_c_498_n N_A_944_107#_M1005_g 0.0317217f $X=6.41 $Y=2.585
+ $X2=0 $Y2=0
cc_392 N_A_1214_107#_c_501_n N_A_1678_81#_M1001_g 0.0873839f $X=8.37 $Y=2.775
+ $X2=0 $Y2=0
cc_393 N_A_1214_107#_c_507_n N_A_1678_81#_M1001_g 2.51395e-19 $X=8.405 $Y=2.38
+ $X2=0 $Y2=0
cc_394 N_A_1214_107#_c_501_n N_A_1678_81#_c_699_n 0.00530376f $X=8.37 $Y=2.775
+ $X2=0 $Y2=0
cc_395 N_A_1214_107#_c_516_p N_A_1480_107#_c_773_n 0.0258964f $X=7.19 $Y=1.25
+ $X2=5.76 $Y2=0.058
cc_396 N_A_1214_107#_M1002_g N_A_1480_107#_c_773_n 0.00157677f $X=7.15 $Y=0.745
+ $X2=5.76 $Y2=0.058
cc_397 N_A_1214_107#_M1000_g N_A_1480_107#_c_787_n 0.00631423f $X=8.37 $Y=3.175
+ $X2=0 $Y2=0
cc_398 N_A_1214_107#_c_506_n N_A_1480_107#_c_787_n 0.0144434f $X=8.01 $Y=2.345
+ $X2=0 $Y2=0
cc_399 N_A_1214_107#_c_507_n N_A_1480_107#_c_787_n 0.00163176f $X=8.405 $Y=2.38
+ $X2=0 $Y2=0
cc_400 N_A_1214_107#_M1000_g N_A_1480_107#_c_788_n 0.00668305f $X=8.37 $Y=3.175
+ $X2=0 $Y2=0
cc_401 N_A_1214_107#_c_496_n N_A_1480_107#_c_775_n 0.0126237f $X=7.84 $Y=1.67
+ $X2=0 $Y2=0
cc_402 N_A_1214_107#_c_516_p N_A_1480_107#_c_776_n 0.0131377f $X=7.19 $Y=1.25
+ $X2=0 $Y2=0
cc_403 N_A_1214_107#_c_496_n N_A_1480_107#_c_776_n 0.0125551f $X=7.84 $Y=1.67
+ $X2=0 $Y2=0
cc_404 N_A_1214_107#_M1002_g N_A_1480_107#_c_776_n 0.00163512f $X=7.15 $Y=0.745
+ $X2=0 $Y2=0
cc_405 N_A_1214_107#_c_501_n N_A_1480_107#_c_791_n 0.015212f $X=8.37 $Y=2.775
+ $X2=0 $Y2=0
cc_406 N_A_1214_107#_M1000_g N_A_1480_107#_c_791_n 0.025395f $X=8.37 $Y=3.175
+ $X2=0 $Y2=0
cc_407 N_A_1214_107#_c_507_n N_A_1480_107#_c_791_n 0.0372062f $X=8.405 $Y=2.38
+ $X2=0 $Y2=0
cc_408 N_A_1214_107#_c_496_n N_A_1480_107#_c_777_n 0.0130053f $X=7.84 $Y=1.67
+ $X2=0 $Y2=0
cc_409 N_A_1214_107#_c_519_p N_A_1480_107#_c_777_n 0.00541191f $X=7.925 $Y=2.215
+ $X2=0 $Y2=0
cc_410 N_A_1214_107#_c_501_n N_A_1480_107#_c_778_n 0.00314557f $X=8.37 $Y=2.775
+ $X2=0 $Y2=0
cc_411 N_A_1214_107#_c_507_n N_A_1480_107#_c_778_n 0.0131973f $X=8.405 $Y=2.38
+ $X2=0 $Y2=0
cc_412 N_A_1214_107#_c_501_n N_A_1480_107#_c_779_n 0.00381302f $X=8.37 $Y=2.775
+ $X2=0 $Y2=0
cc_413 N_A_1214_107#_c_519_p N_A_1480_107#_c_779_n 0.0131378f $X=7.925 $Y=2.215
+ $X2=0 $Y2=0
cc_414 N_A_1214_107#_c_507_n N_A_1480_107#_c_779_n 0.0121659f $X=8.405 $Y=2.38
+ $X2=0 $Y2=0
cc_415 N_A_1214_107#_c_501_n N_A_1480_107#_c_794_n 0.00590994f $X=8.37 $Y=2.775
+ $X2=0 $Y2=0
cc_416 N_A_1214_107#_c_507_n N_A_1480_107#_c_794_n 0.0197395f $X=8.405 $Y=2.38
+ $X2=0 $Y2=0
cc_417 N_A_1214_107#_M1000_g N_VPWR_c_902_n 0.00788454f $X=8.37 $Y=3.175 $X2=0
+ $Y2=0
cc_418 N_A_1214_107#_M1000_g N_VPWR_c_908_n 0.0310706f $X=8.37 $Y=3.175 $X2=0
+ $Y2=0
cc_419 N_A_1214_107#_c_505_n N_VPWR_c_908_n 0.0118571f $X=6.41 $Y=2.75 $X2=0
+ $Y2=0
cc_420 N_A_1214_107#_c_498_n N_A_489_107#_c_1004_n 0.0123662f $X=6.41 $Y=2.585
+ $X2=0 $Y2=0
cc_421 N_A_1214_107#_c_498_n N_A_489_107#_c_1006_n 0.0681055f $X=6.41 $Y=2.585
+ $X2=0 $Y2=0
cc_422 N_A_1214_107#_c_505_n N_A_489_107#_c_1007_n 0.0220429f $X=6.41 $Y=2.75
+ $X2=0 $Y2=0
cc_423 N_A_1214_107#_c_491_n N_A_489_107#_c_989_n 0.0288784f $X=6.21 $Y=0.745
+ $X2=0 $Y2=0
cc_424 N_A_1214_107#_c_492_n N_A_489_107#_c_989_n 0.0209364f $X=7.105 $Y=0.35
+ $X2=0 $Y2=0
cc_425 N_A_1214_107#_c_516_p N_A_489_107#_c_989_n 0.0639142f $X=7.19 $Y=1.25
+ $X2=0 $Y2=0
cc_426 N_A_1214_107#_M1002_g N_A_489_107#_c_989_n 0.0066279f $X=7.15 $Y=0.745
+ $X2=0 $Y2=0
cc_427 N_A_1214_107#_c_505_n N_A_489_107#_c_1015_n 0.0331012f $X=6.41 $Y=2.75
+ $X2=0 $Y2=0
cc_428 N_A_1214_107#_c_505_n N_A_489_107#_c_990_n 0.0331012f $X=6.41 $Y=2.75
+ $X2=0 $Y2=0
cc_429 N_A_1214_107#_c_512_p N_A_489_107#_c_990_n 0.0123662f $X=7.275 $Y=1.67
+ $X2=0 $Y2=0
cc_430 N_A_1214_107#_c_498_n N_A_489_107#_c_990_n 0.0711162f $X=6.41 $Y=2.585
+ $X2=0 $Y2=0
cc_431 N_A_1214_107#_M1002_g N_A_489_107#_c_990_n 0.0270811f $X=7.15 $Y=0.745
+ $X2=0 $Y2=0
cc_432 N_A_1214_107#_c_491_n N_VGND_c_1156_n 0.0283847f $X=6.21 $Y=0.745 $X2=0
+ $Y2=0
cc_433 N_A_1214_107#_c_494_n N_VGND_c_1156_n 0.00330668f $X=6.415 $Y=0.35 $X2=0
+ $Y2=0
cc_434 N_A_1214_107#_c_498_n N_VGND_c_1156_n 7.35778e-19 $X=6.41 $Y=2.585 $X2=0
+ $Y2=0
cc_435 N_A_1214_107#_c_491_n N_VGND_c_1162_n 0.0365733f $X=6.21 $Y=0.745 $X2=0
+ $Y2=0
cc_436 N_A_1214_107#_c_492_n N_VGND_c_1162_n 0.0350102f $X=7.105 $Y=0.35 $X2=0
+ $Y2=0
cc_437 N_A_1214_107#_c_494_n N_VGND_c_1162_n 0.0121556f $X=6.415 $Y=0.35 $X2=0
+ $Y2=0
cc_438 N_A_1214_107#_c_516_p N_VGND_c_1162_n 0.0209621f $X=7.19 $Y=1.25 $X2=0
+ $Y2=0
cc_439 N_A_1214_107#_M1002_g N_VGND_c_1162_n 0.0181231f $X=7.15 $Y=0.745 $X2=0
+ $Y2=0
cc_440 N_A_944_107#_M1019_g N_A_1678_81#_c_693_n 0.0450296f $X=7.93 $Y=0.745
+ $X2=0 $Y2=0
cc_441 N_A_944_107#_c_582_n N_A_1678_81#_M1001_g 0.0026662f $X=7.475 $Y=2.515
+ $X2=0 $Y2=0
cc_442 N_A_944_107#_M1019_g N_A_1678_81#_c_710_n 2.62155e-19 $X=7.93 $Y=0.745
+ $X2=0 $Y2=0
cc_443 N_A_944_107#_c_582_n N_A_1678_81#_c_699_n 0.0450296f $X=7.475 $Y=2.515
+ $X2=0 $Y2=0
cc_444 N_A_944_107#_M1019_g N_A_1480_107#_c_773_n 0.0152268f $X=7.93 $Y=0.745
+ $X2=5.76 $Y2=0.058
cc_445 N_A_944_107#_c_582_n N_A_1480_107#_c_787_n 0.00443378f $X=7.475 $Y=2.515
+ $X2=0 $Y2=0
cc_446 N_A_944_107#_M1007_g N_A_1480_107#_c_787_n 0.0139459f $X=7.475 $Y=3.34
+ $X2=0 $Y2=0
cc_447 N_A_944_107#_M1007_g N_A_1480_107#_c_788_n 0.0174441f $X=7.475 $Y=3.34
+ $X2=0 $Y2=0
cc_448 N_A_944_107#_M1019_g N_A_1480_107#_c_775_n 0.0318296f $X=7.93 $Y=0.745
+ $X2=0 $Y2=0
cc_449 N_A_944_107#_c_582_n N_A_1480_107#_c_776_n 0.00199138f $X=7.475 $Y=2.515
+ $X2=0 $Y2=0
cc_450 N_A_944_107#_M1019_g N_A_1480_107#_c_776_n 0.00247317f $X=7.93 $Y=0.745
+ $X2=0 $Y2=0
cc_451 N_A_944_107#_M1019_g N_A_1480_107#_c_777_n 0.0112361f $X=7.93 $Y=0.745
+ $X2=0 $Y2=0
cc_452 N_A_944_107#_c_582_n N_A_1480_107#_c_779_n 0.00302757f $X=7.475 $Y=2.515
+ $X2=0 $Y2=0
cc_453 N_A_944_107#_c_593_n N_VPWR_c_899_n 0.00715793f $X=6.02 $Y=2.515 $X2=0
+ $Y2=0
cc_454 N_A_944_107#_c_601_n N_VPWR_c_899_n 0.00445234f $X=5.92 $Y=2.265 $X2=0
+ $Y2=0
cc_455 N_A_944_107#_M1023_d N_VPWR_c_908_n 0.00479598f $X=4.79 $Y=2.935 $X2=0
+ $Y2=0
cc_456 N_A_944_107#_c_593_n N_VPWR_c_908_n 0.0204412f $X=6.02 $Y=2.515 $X2=0
+ $Y2=0
cc_457 N_A_944_107#_M1007_g N_VPWR_c_908_n 0.0274961f $X=7.475 $Y=3.34 $X2=0
+ $Y2=0
cc_458 N_A_944_107#_c_586_n N_VPWR_c_908_n 0.0117486f $X=4.93 $Y=3.175 $X2=0
+ $Y2=0
cc_459 N_A_944_107#_c_586_n N_A_489_107#_c_986_n 0.00522802f $X=4.93 $Y=3.175
+ $X2=0 $Y2=0
cc_460 N_A_944_107#_c_586_n N_A_489_107#_c_997_n 0.0129653f $X=4.93 $Y=3.175
+ $X2=0 $Y2=0
cc_461 N_A_944_107#_c_586_n N_A_489_107#_c_1049_n 0.0230778f $X=4.93 $Y=3.175
+ $X2=0 $Y2=0
cc_462 N_A_944_107#_M1023_d N_A_489_107#_c_998_n 0.00215778f $X=4.79 $Y=2.935
+ $X2=0 $Y2=0
cc_463 N_A_944_107#_c_586_n N_A_489_107#_c_998_n 0.0110919f $X=4.93 $Y=3.175
+ $X2=0 $Y2=0
cc_464 N_A_944_107#_c_593_n N_A_489_107#_c_1003_n 0.00280691f $X=6.02 $Y=2.515
+ $X2=0 $Y2=0
cc_465 N_A_944_107#_c_601_n N_A_489_107#_c_1003_n 0.00316556f $X=5.92 $Y=2.265
+ $X2=0 $Y2=0
cc_466 N_A_944_107#_c_586_n N_A_489_107#_c_1003_n 0.0751475f $X=4.93 $Y=3.175
+ $X2=0 $Y2=0
cc_467 N_A_944_107#_c_601_n N_A_489_107#_c_1004_n 0.0383384f $X=5.92 $Y=2.265
+ $X2=0 $Y2=0
cc_468 N_A_944_107#_c_633_n N_A_489_107#_c_1004_n 0.012841f $X=5.755 $Y=1.34
+ $X2=0 $Y2=0
cc_469 N_A_944_107#_c_586_n N_A_489_107#_c_1005_n 0.0137874f $X=4.93 $Y=3.175
+ $X2=0 $Y2=0
cc_470 N_A_944_107#_c_593_n N_A_489_107#_c_1006_n 0.0429996f $X=6.02 $Y=2.515
+ $X2=0 $Y2=0
cc_471 N_A_944_107#_c_601_n N_A_489_107#_c_1006_n 0.00556771f $X=5.92 $Y=2.265
+ $X2=0 $Y2=0
cc_472 N_A_944_107#_c_593_n N_A_489_107#_c_1007_n 0.00673315f $X=6.02 $Y=2.515
+ $X2=0 $Y2=0
cc_473 N_A_944_107#_M1007_g N_A_489_107#_c_1007_n 0.00458401f $X=7.475 $Y=3.34
+ $X2=0 $Y2=0
cc_474 N_A_944_107#_c_593_n N_A_489_107#_c_1013_n 0.0020308f $X=6.02 $Y=2.515
+ $X2=0 $Y2=0
cc_475 N_A_944_107#_M1007_g N_A_489_107#_c_1013_n 0.0125158f $X=7.475 $Y=3.34
+ $X2=0 $Y2=0
cc_476 N_A_944_107#_M1005_g N_A_489_107#_c_989_n 5.7526e-19 $X=5.82 $Y=0.745
+ $X2=0 $Y2=0
cc_477 N_A_944_107#_c_596_n N_A_489_107#_c_1015_n 0.00756804f $X=7.225 $Y=2.265
+ $X2=0 $Y2=0
cc_478 N_A_944_107#_M1007_g N_A_489_107#_c_1015_n 0.00870633f $X=7.475 $Y=3.34
+ $X2=0 $Y2=0
cc_479 N_A_944_107#_c_593_n N_A_489_107#_c_990_n 0.00202053f $X=6.02 $Y=2.515
+ $X2=0 $Y2=0
cc_480 N_A_944_107#_c_596_n N_A_489_107#_c_990_n 0.048027f $X=7.225 $Y=2.265
+ $X2=0 $Y2=0
cc_481 N_A_944_107#_c_582_n N_A_489_107#_c_990_n 0.00618906f $X=7.475 $Y=2.515
+ $X2=0 $Y2=0
cc_482 N_A_944_107#_M1007_g N_A_489_107#_c_990_n 0.014088f $X=7.475 $Y=3.34
+ $X2=0 $Y2=0
cc_483 N_A_944_107#_c_588_n N_VGND_c_1154_n 0.0257598f $X=4.86 $Y=0.745 $X2=0
+ $Y2=0
cc_484 N_A_944_107#_c_585_n N_VGND_c_1156_n 0.00150218f $X=4.93 $Y=1.175 $X2=0
+ $Y2=0
cc_485 N_A_944_107#_c_587_n N_VGND_c_1156_n 0.0298111f $X=5.59 $Y=1.26 $X2=0
+ $Y2=0
cc_486 N_A_944_107#_c_588_n N_VGND_c_1156_n 0.0368304f $X=4.86 $Y=0.745 $X2=0
+ $Y2=0
cc_487 N_A_944_107#_c_633_n N_VGND_c_1156_n 0.0158209f $X=5.755 $Y=1.34 $X2=0
+ $Y2=0
cc_488 N_A_944_107#_M1005_g N_VGND_c_1156_n 0.0322328f $X=5.82 $Y=0.745 $X2=0
+ $Y2=0
cc_489 N_A_944_107#_M1019_g N_VGND_c_1158_n 0.00731985f $X=7.93 $Y=0.745 $X2=0
+ $Y2=0
cc_490 N_A_944_107#_M1019_g N_VGND_c_1162_n 0.0168423f $X=7.93 $Y=0.745 $X2=0
+ $Y2=0
cc_491 N_A_944_107#_c_587_n N_VGND_c_1162_n 0.00773943f $X=5.59 $Y=1.26 $X2=0
+ $Y2=0
cc_492 N_A_944_107#_c_588_n N_VGND_c_1162_n 0.0277681f $X=4.86 $Y=0.745 $X2=0
+ $Y2=0
cc_493 N_A_944_107#_c_633_n N_VGND_c_1162_n 0.00480816f $X=5.755 $Y=1.34 $X2=0
+ $Y2=0
cc_494 N_A_944_107#_M1005_g N_VGND_c_1162_n 0.010759f $X=5.82 $Y=0.745 $X2=0
+ $Y2=0
cc_495 N_A_1678_81#_M1001_g N_A_1480_107#_M1011_g 0.0225109f $X=9.08 $Y=3.175
+ $X2=0 $Y2=0
cc_496 N_A_1678_81#_c_702_n N_A_1480_107#_M1011_g 0.0285799f $X=10.38 $Y=2.27
+ $X2=0 $Y2=0
cc_497 N_A_1678_81#_c_703_n N_A_1480_107#_M1011_g 0.00224589f $X=10.465 $Y=2.185
+ $X2=0 $Y2=0
cc_498 N_A_1678_81#_c_704_n N_A_1480_107#_M1011_g 0.0143362f $X=9.55 $Y=2.27
+ $X2=0 $Y2=0
cc_499 N_A_1678_81#_c_696_n N_A_1480_107#_M1013_g 0.0175744f $X=9.58 $Y=1.075
+ $X2=0 $Y2=0
cc_500 N_A_1678_81#_c_697_n N_A_1480_107#_M1013_g 0.0123129f $X=10.38 $Y=1.49
+ $X2=0 $Y2=0
cc_501 N_A_1678_81#_c_699_n N_A_1480_107#_M1013_g 0.00688645f $X=9.08 $Y=1.41
+ $X2=0 $Y2=0
cc_502 N_A_1678_81#_c_702_n N_A_1480_107#_M1021_g 0.00162228f $X=10.38 $Y=2.27
+ $X2=11.28 $Y2=0
cc_503 N_A_1678_81#_c_703_n N_A_1480_107#_M1021_g 0.00150592f $X=10.465 $Y=2.185
+ $X2=11.28 $Y2=0
cc_504 N_A_1678_81#_c_693_n N_A_1480_107#_c_773_n 8.5452e-19 $X=8.64 $Y=1.065
+ $X2=5.76 $Y2=0.058
cc_505 N_A_1678_81#_c_710_n N_A_1480_107#_c_775_n 0.0137299f $X=8.705 $Y=1.23
+ $X2=0 $Y2=0
cc_506 N_A_1678_81#_c_699_n N_A_1480_107#_c_775_n 0.00156493f $X=9.08 $Y=1.41
+ $X2=0 $Y2=0
cc_507 N_A_1678_81#_M1001_g N_A_1480_107#_c_791_n 0.0119534f $X=9.08 $Y=3.175
+ $X2=0 $Y2=0
cc_508 N_A_1678_81#_c_704_n N_A_1480_107#_c_791_n 7.8365e-19 $X=9.55 $Y=2.27
+ $X2=0 $Y2=0
cc_509 N_A_1678_81#_M1001_g N_A_1480_107#_c_777_n 0.00141763f $X=9.08 $Y=3.175
+ $X2=0 $Y2=0
cc_510 N_A_1678_81#_c_710_n N_A_1480_107#_c_777_n 0.0294737f $X=8.705 $Y=1.23
+ $X2=0 $Y2=0
cc_511 N_A_1678_81#_c_699_n N_A_1480_107#_c_777_n 0.00578462f $X=9.08 $Y=1.41
+ $X2=0 $Y2=0
cc_512 N_A_1678_81#_c_710_n N_A_1480_107#_c_778_n 0.0157522f $X=8.705 $Y=1.23
+ $X2=0 $Y2=0
cc_513 N_A_1678_81#_c_699_n N_A_1480_107#_c_778_n 0.00886323f $X=9.08 $Y=1.41
+ $X2=0 $Y2=0
cc_514 N_A_1678_81#_M1001_g N_A_1480_107#_c_794_n 0.0272818f $X=9.08 $Y=3.175
+ $X2=0 $Y2=0
cc_515 N_A_1678_81#_c_704_n N_A_1480_107#_c_794_n 0.016701f $X=9.55 $Y=2.27
+ $X2=0 $Y2=0
cc_516 N_A_1678_81#_M1001_g N_A_1480_107#_c_780_n 0.00639982f $X=9.08 $Y=3.175
+ $X2=0 $Y2=0
cc_517 N_A_1678_81#_c_695_n N_A_1480_107#_c_780_n 0.00270798f $X=9.415 $Y=1.49
+ $X2=0 $Y2=0
cc_518 N_A_1678_81#_c_710_n N_A_1480_107#_c_780_n 0.00986478f $X=8.705 $Y=1.23
+ $X2=0 $Y2=0
cc_519 N_A_1678_81#_c_699_n N_A_1480_107#_c_780_n 0.00244186f $X=9.08 $Y=1.41
+ $X2=0 $Y2=0
cc_520 N_A_1678_81#_M1001_g N_A_1480_107#_c_853_n 3.92856e-19 $X=9.08 $Y=3.175
+ $X2=0 $Y2=0
cc_521 N_A_1678_81#_c_697_n N_A_1480_107#_c_853_n 0.0220177f $X=10.38 $Y=1.49
+ $X2=0 $Y2=0
cc_522 N_A_1678_81#_c_703_n N_A_1480_107#_c_853_n 0.0177091f $X=10.465 $Y=2.185
+ $X2=0 $Y2=0
cc_523 N_A_1678_81#_M1001_g N_A_1480_107#_c_781_n 0.0340235f $X=9.08 $Y=3.175
+ $X2=0 $Y2=0
cc_524 N_A_1678_81#_c_695_n N_A_1480_107#_c_781_n 0.0245013f $X=9.415 $Y=1.49
+ $X2=0 $Y2=0
cc_525 N_A_1678_81#_c_702_n N_A_1480_107#_c_781_n 0.0320585f $X=10.38 $Y=2.27
+ $X2=0 $Y2=0
cc_526 N_A_1678_81#_c_697_n N_A_1480_107#_c_781_n 0.00598559f $X=10.38 $Y=1.49
+ $X2=0 $Y2=0
cc_527 N_A_1678_81#_c_704_n N_A_1480_107#_c_781_n 0.0257001f $X=9.55 $Y=2.27
+ $X2=0 $Y2=0
cc_528 N_A_1678_81#_c_698_n N_A_1480_107#_c_781_n 0.0202343f $X=9.58 $Y=1.49
+ $X2=0 $Y2=0
cc_529 N_A_1678_81#_c_702_n N_A_1480_107#_c_782_n 0.00332534f $X=10.38 $Y=2.27
+ $X2=0 $Y2=0
cc_530 N_A_1678_81#_c_697_n N_A_1480_107#_c_782_n 0.0304195f $X=10.38 $Y=1.49
+ $X2=0 $Y2=0
cc_531 N_A_1678_81#_c_703_n N_A_1480_107#_c_782_n 0.0380626f $X=10.465 $Y=2.185
+ $X2=0 $Y2=0
cc_532 N_A_1678_81#_c_698_n N_A_1480_107#_c_782_n 0.00483699f $X=9.58 $Y=1.49
+ $X2=0 $Y2=0
cc_533 N_A_1678_81#_c_699_n N_A_1480_107#_c_782_n 0.0225109f $X=9.08 $Y=1.41
+ $X2=0 $Y2=0
cc_534 N_A_1678_81#_c_702_n N_VPWR_M1011_d 0.00389681f $X=10.38 $Y=2.27
+ $X2=-0.33 $Y2=-0.265
cc_535 N_A_1678_81#_M1001_g N_VPWR_c_902_n 0.0614541f $X=9.08 $Y=3.175 $X2=0
+ $Y2=0
cc_536 N_A_1678_81#_c_704_n N_VPWR_c_902_n 0.0138343f $X=9.55 $Y=2.27 $X2=0
+ $Y2=0
cc_537 N_A_1678_81#_M1001_g N_VPWR_c_905_n 0.00880927f $X=9.08 $Y=3.175 $X2=0
+ $Y2=0
cc_538 N_A_1678_81#_c_702_n N_VPWR_c_905_n 0.0445012f $X=10.38 $Y=2.27 $X2=0
+ $Y2=0
cc_539 N_A_1678_81#_c_704_n N_VPWR_c_905_n 0.0106243f $X=9.55 $Y=2.27 $X2=0
+ $Y2=0
cc_540 N_A_1678_81#_c_702_n N_Q_c_1137_n 0.00324147f $X=10.38 $Y=2.27 $X2=0
+ $Y2=0
cc_541 N_A_1678_81#_c_697_n N_Q_c_1137_n 0.00555768f $X=10.38 $Y=1.49 $X2=0
+ $Y2=0
cc_542 N_A_1678_81#_c_703_n N_Q_c_1137_n 0.0181192f $X=10.465 $Y=2.185 $X2=0
+ $Y2=0
cc_543 N_A_1678_81#_c_693_n N_VGND_c_1158_n 0.048961f $X=8.64 $Y=1.065 $X2=0
+ $Y2=0
cc_544 N_A_1678_81#_c_695_n N_VGND_c_1158_n 0.00958505f $X=9.415 $Y=1.49 $X2=0
+ $Y2=0
cc_545 N_A_1678_81#_c_696_n N_VGND_c_1158_n 0.00361551f $X=9.58 $Y=1.075 $X2=0
+ $Y2=0
cc_546 N_A_1678_81#_c_710_n N_VGND_c_1158_n 0.0243389f $X=8.705 $Y=1.23 $X2=0
+ $Y2=0
cc_547 N_A_1678_81#_c_699_n N_VGND_c_1158_n 0.00922173f $X=9.08 $Y=1.41 $X2=0
+ $Y2=0
cc_548 N_A_1678_81#_c_696_n N_VGND_c_1160_n 0.0288375f $X=9.58 $Y=1.075 $X2=0
+ $Y2=0
cc_549 N_A_1678_81#_c_697_n N_VGND_c_1160_n 0.0460568f $X=10.38 $Y=1.49 $X2=0
+ $Y2=0
cc_550 N_A_1678_81#_c_696_n N_VGND_c_1162_n 0.0177898f $X=9.58 $Y=1.075 $X2=0
+ $Y2=0
cc_551 N_A_1678_81#_c_710_n N_VGND_c_1162_n 0.00140034f $X=8.705 $Y=1.23 $X2=0
+ $Y2=0
cc_552 N_A_1678_81#_c_699_n N_VGND_c_1162_n 0.00363195f $X=9.08 $Y=1.41 $X2=0
+ $Y2=0
cc_553 N_A_1480_107#_c_787_n N_VPWR_c_902_n 0.00258863f $X=7.865 $Y=3.09 $X2=0
+ $Y2=0
cc_554 N_A_1480_107#_c_788_n N_VPWR_c_902_n 0.0149851f $X=7.865 $Y=3.59 $X2=0
+ $Y2=0
cc_555 N_A_1480_107#_c_791_n N_VPWR_c_902_n 0.0165596f $X=8.75 $Y=2.74 $X2=0
+ $Y2=0
cc_556 N_A_1480_107#_M1011_g N_VPWR_c_905_n 0.0256009f $X=9.94 $Y=2.425 $X2=0
+ $Y2=0
cc_557 N_A_1480_107#_M1021_g N_VPWR_c_905_n 0.0675823f $X=10.835 $Y=2.965 $X2=0
+ $Y2=0
cc_558 N_A_1480_107#_c_782_n N_VPWR_c_905_n 7.06093e-19 $X=10.845 $Y=1.75 $X2=0
+ $Y2=0
cc_559 N_A_1480_107#_M1021_g N_VPWR_c_908_n 0.0130327f $X=10.835 $Y=2.965 $X2=0
+ $Y2=0
cc_560 N_A_1480_107#_c_788_n N_VPWR_c_908_n 0.0457632f $X=7.865 $Y=3.59 $X2=0
+ $Y2=0
cc_561 N_A_1480_107#_c_791_n N_VPWR_c_908_n 5.86364e-19 $X=8.75 $Y=2.74 $X2=0
+ $Y2=0
cc_562 N_A_1480_107#_c_788_n N_A_489_107#_c_1007_n 0.0030198f $X=7.865 $Y=3.59
+ $X2=0 $Y2=0
cc_563 N_A_1480_107#_c_787_n N_A_489_107#_c_1015_n 0.00582067f $X=7.865 $Y=3.09
+ $X2=0 $Y2=0
cc_564 N_A_1480_107#_c_788_n N_A_489_107#_c_1015_n 0.015266f $X=7.865 $Y=3.59
+ $X2=0 $Y2=0
cc_565 N_A_1480_107#_M1021_g N_Q_c_1137_n 0.0404155f $X=10.835 $Y=2.965 $X2=0
+ $Y2=0
cc_566 N_A_1480_107#_M1020_g N_Q_c_1137_n 0.0255176f $X=10.845 $Y=0.91 $X2=0
+ $Y2=0
cc_567 N_A_1480_107#_c_782_n N_Q_c_1137_n 0.0332302f $X=10.845 $Y=1.75 $X2=0
+ $Y2=0
cc_568 N_A_1480_107#_M1013_g N_VGND_c_1158_n 0.00369955f $X=9.97 $Y=1.075 $X2=0
+ $Y2=0
cc_569 N_A_1480_107#_c_773_n N_VGND_c_1158_n 0.0109217f $X=7.54 $Y=0.745 $X2=0
+ $Y2=0
cc_570 N_A_1480_107#_c_775_n N_VGND_c_1158_n 0.00830264f $X=8.19 $Y=1.16 $X2=0
+ $Y2=0
cc_571 N_A_1480_107#_M1013_g N_VGND_c_1160_n 0.0421792f $X=9.97 $Y=1.075 $X2=0
+ $Y2=0
cc_572 N_A_1480_107#_M1020_g N_VGND_c_1160_n 0.0564366f $X=10.845 $Y=0.91 $X2=0
+ $Y2=0
cc_573 N_A_1480_107#_c_782_n N_VGND_c_1160_n 0.00149477f $X=10.845 $Y=1.75 $X2=0
+ $Y2=0
cc_574 N_A_1480_107#_M1002_d N_VGND_c_1162_n 0.00221032f $X=7.4 $Y=0.535 $X2=0
+ $Y2=0
cc_575 N_A_1480_107#_M1013_g N_VGND_c_1162_n 0.00672879f $X=9.97 $Y=1.075 $X2=0
+ $Y2=0
cc_576 N_A_1480_107#_M1020_g N_VGND_c_1162_n 0.0122818f $X=10.845 $Y=0.91 $X2=0
+ $Y2=0
cc_577 N_A_1480_107#_c_773_n N_VGND_c_1162_n 0.0258005f $X=7.54 $Y=0.745 $X2=0
+ $Y2=0
cc_578 N_A_1480_107#_c_775_n N_VGND_c_1162_n 0.0179793f $X=8.19 $Y=1.16 $X2=0
+ $Y2=0
cc_579 N_VPWR_c_908_n A_362_587# 0.00875788f $X=10.73 $Y=3.59 $X2=0 $Y2=3.985
cc_580 N_VPWR_c_908_n N_A_489_107#_M1017_d 0.00221032f $X=10.73 $Y=3.59 $X2=0
+ $Y2=0
cc_581 N_VPWR_c_896_n N_A_489_107#_c_991_n 0.0181714f $X=4.2 $Y=3.59 $X2=11.28
+ $Y2=4.07
cc_582 N_VPWR_c_908_n N_A_489_107#_c_991_n 0.0393884f $X=10.73 $Y=3.59 $X2=11.28
+ $Y2=4.07
cc_583 N_VPWR_c_896_n N_A_489_107#_c_994_n 0.044689f $X=4.2 $Y=3.59 $X2=0 $Y2=0
cc_584 N_VPWR_c_908_n N_A_489_107#_c_994_n 0.0167076f $X=10.73 $Y=3.59 $X2=0
+ $Y2=0
cc_585 N_VPWR_c_896_n N_A_489_107#_c_997_n 0.00617953f $X=4.2 $Y=3.59 $X2=0
+ $Y2=0
cc_586 N_VPWR_c_908_n N_A_489_107#_c_997_n 0.00510093f $X=10.73 $Y=3.59 $X2=0
+ $Y2=0
cc_587 N_VPWR_c_896_n N_A_489_107#_c_1049_n 0.0421578f $X=4.2 $Y=3.59 $X2=0
+ $Y2=0
cc_588 N_VPWR_c_908_n N_A_489_107#_c_1049_n 0.0190049f $X=10.73 $Y=3.59 $X2=0
+ $Y2=0
cc_589 N_VPWR_c_899_n N_A_489_107#_c_998_n 0.00479486f $X=5.63 $Y=2.75 $X2=0
+ $Y2=0
cc_590 N_VPWR_c_908_n N_A_489_107#_c_998_n 0.0282546f $X=10.73 $Y=3.59 $X2=0
+ $Y2=0
cc_591 N_VPWR_c_896_n N_A_489_107#_c_1001_n 0.00555087f $X=4.2 $Y=3.59 $X2=0
+ $Y2=0
cc_592 N_VPWR_c_908_n N_A_489_107#_c_1001_n 0.00656746f $X=10.73 $Y=3.59 $X2=0
+ $Y2=0
cc_593 N_VPWR_c_899_n N_A_489_107#_c_1003_n 0.0738087f $X=5.63 $Y=2.75 $X2=0
+ $Y2=0
cc_594 N_VPWR_c_908_n N_A_489_107#_c_1003_n 0.0194693f $X=10.73 $Y=3.59 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_899_n N_A_489_107#_c_1004_n 0.0130751f $X=5.63 $Y=2.75 $X2=0
+ $Y2=0
cc_596 N_VPWR_c_899_n N_A_489_107#_c_1006_n 0.0415321f $X=5.63 $Y=2.75 $X2=0
+ $Y2=0
cc_597 N_VPWR_c_908_n N_A_489_107#_c_1006_n 0.0186563f $X=10.73 $Y=3.59 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_908_n N_A_489_107#_c_1007_n 0.0430806f $X=10.73 $Y=3.59 $X2=0
+ $Y2=0
cc_599 N_VPWR_c_899_n N_A_489_107#_c_1010_n 0.00753478f $X=5.63 $Y=2.75 $X2=0
+ $Y2=0
cc_600 N_VPWR_c_908_n N_A_489_107#_c_1010_n 0.00654857f $X=10.73 $Y=3.59 $X2=0
+ $Y2=0
cc_601 N_VPWR_c_908_n N_A_489_107#_c_1013_n 0.0433999f $X=10.73 $Y=3.59 $X2=0
+ $Y2=0
cc_602 N_VPWR_c_896_n N_A_489_107#_c_1014_n 0.0128396f $X=4.2 $Y=3.59 $X2=0
+ $Y2=0
cc_603 N_VPWR_c_908_n N_A_489_107#_c_1014_n 6.35456e-19 $X=10.73 $Y=3.59 $X2=0
+ $Y2=0
cc_604 N_VPWR_c_896_n A_660_587# 0.00962253f $X=4.2 $Y=3.59 $X2=0 $Y2=3.985
cc_605 N_VPWR_c_908_n A_660_587# 9.33524e-19 $X=10.73 $Y=3.59 $X2=0 $Y2=3.985
cc_606 N_VPWR_c_902_n A_1724_593# 0.00665056f $X=9.47 $Y=3.175 $X2=0 $Y2=3.985
cc_607 N_VPWR_c_905_n N_Q_c_1137_n 0.075681f $X=10.445 $Y=2.62 $X2=5.76 $Y2=4.07
cc_608 N_VPWR_c_908_n N_Q_c_1137_n 0.0443798f $X=10.73 $Y=3.59 $X2=5.76 $Y2=4.07
cc_609 N_A_489_107#_c_984_n N_VGND_c_1154_n 0.0135272f $X=3.515 $Y=0.83 $X2=0
+ $Y2=0
cc_610 N_A_489_107#_c_1019_n N_VGND_c_1154_n 0.00426018f $X=3.6 $Y=1.175 $X2=0
+ $Y2=0
cc_611 N_A_489_107#_c_985_n N_VGND_c_1154_n 0.0243515f $X=4.03 $Y=1.26 $X2=0
+ $Y2=0
cc_612 N_A_489_107#_c_984_n N_VGND_c_1162_n 0.0325347f $X=3.515 $Y=0.83 $X2=0
+ $Y2=0
cc_613 N_A_489_107#_c_985_n N_VGND_c_1162_n 0.0062907f $X=4.03 $Y=1.26 $X2=0
+ $Y2=0
cc_614 N_A_489_107#_c_987_n N_VGND_c_1162_n 0.0226044f $X=2.585 $Y=0.745 $X2=0
+ $Y2=0
cc_615 N_A_489_107#_c_989_n N_VGND_c_1162_n 0.0217482f $X=6.76 $Y=0.755 $X2=0
+ $Y2=0
cc_616 N_A_489_107#_c_984_n A_645_107# 0.00382847f $X=3.515 $Y=0.83 $X2=0 $Y2=0
cc_617 N_Q_c_1137_n N_VGND_c_1160_n 0.0511958f $X=11.235 $Y=0.68 $X2=0 $Y2=0
cc_618 N_Q_c_1137_n N_VGND_c_1162_n 0.0329326f $X=11.235 $Y=0.68 $X2=0 $Y2=0
cc_619 N_VGND_c_1162_n A_347_107# 0.00286287f $X=10.76 $Y=0.48 $X2=0 $Y2=0
cc_620 N_VGND_c_1162_n A_645_107# 0.00173403f $X=10.76 $Y=0.48 $X2=0 $Y2=0
cc_621 N_VGND_c_1158_n A_1636_107# 0.00576659f $X=9.08 $Y=0.48 $X2=0 $Y2=0
cc_622 N_VGND_c_1162_n A_1636_107# 7.90755e-19 $X=10.76 $Y=0.48 $X2=0 $Y2=0
