* File: sky130_fd_sc_hvl__dlrtp_1.spice
* Created: Wed Sep  2 09:05:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__dlrtp_1.pex.spice"
.subckt sky130_fd_sc_hvl__dlrtp_1  VNB VPB D GATE RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1019 N_VGND_M1019_d N_D_M1019_g N_A_32_107#_M1019_s N_VNB_M1019_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1007 N_A_345_107#_M1007_d N_GATE_M1007_g N_VGND_M1019_d N_VNB_M1019_b NHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1018 N_VGND_M1018_d N_A_345_107#_M1018_g N_A_462_107#_M1018_s N_VNB_M1019_b
+ NHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250003 A=0.21 P=1.84 MULT=1
MM1008 A_775_107# N_A_32_107#_M1008_g N_VGND_M1018_d N_VNB_M1019_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250001 SB=250002 A=0.21 P=1.84 MULT=1
MM1012 N_A_917_107#_M1012_d N_A_462_107#_M1012_g A_775_107# N_VNB_M1019_b NHV
+ L=0.5 W=0.42 AD=0.08295 AS=0.0441 PD=0.815 PS=0.63 NRD=31.2132 NRS=13.566 M=1
+ R=0.84 SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1004 A_1096_107# N_A_345_107#_M1004_g N_A_917_107#_M1012_d N_VNB_M1019_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.08295 PD=0.63 PS=0.815 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1009 N_VGND_M1009_d N_A_1138_81#_M1009_g A_1096_107# N_VNB_M1019_b NHV L=0.5
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250003 SB=250000 A=0.21 P=1.84 MULT=1
MM1000 A_1512_107# N_A_917_107#_M1000_g N_A_1138_81#_M1000_s N_VNB_M1019_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1003 N_VGND_M1003_d N_RESET_B_M1003_g A_1512_107# N_VNB_M1019_b NHV L=0.5
+ W=0.42 AD=0.0933154 AS=0.0441 PD=0.822051 PS=0.63 NRD=31.2132 NRS=13.566 M=1
+ R=0.84 SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1015 N_Q_M1015_d N_A_1138_81#_M1015_g N_VGND_M1003_d N_VNB_M1019_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.166635 PD=2.07 PS=1.46795 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1014 N_VPWR_M1014_d N_D_M1014_g N_A_32_107#_M1014_s N_VPB_M1014_b PHV L=0.5
+ W=0.75 AD=0.105 AS=0.21375 PD=1.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1005 N_A_345_107#_M1005_d N_GATE_M1005_g N_VPWR_M1014_d N_VPB_M1014_b PHV
+ L=0.5 W=0.75 AD=0.21375 AS=0.105 PD=2.07 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A_345_107#_M1001_g N_A_462_107#_M1001_s N_VPB_M1014_b
+ PHV L=0.5 W=0.75 AD=0.105 AS=0.21375 PD=1.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250004 A=0.375 P=2.5 MULT=1
MM1010 A_775_491# N_A_32_107#_M1010_g N_VPWR_M1001_d N_VPB_M1014_b PHV L=0.5
+ W=0.75 AD=0.07875 AS=0.105 PD=0.96 PS=1.03 NRD=12.7206 NRS=0 M=1 R=1.5
+ SA=250001 SB=250003 A=0.375 P=2.5 MULT=1
MM1016 N_A_917_107#_M1016_d N_A_345_107#_M1016_g A_775_491# N_VPB_M1014_b PHV
+ L=0.5 W=0.75 AD=0.166635 AS=0.07875 PD=1.46795 PS=0.96 NRD=0 NRS=12.7206 M=1
+ R=1.5 SA=250002 SB=250002 A=0.375 P=2.5 MULT=1
MM1006 A_1096_491# N_A_462_107#_M1006_g N_A_917_107#_M1016_d N_VPB_M1014_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0933154 PD=0.63 PS=0.822051 NRD=22.729 NRS=54.5687
+ M=1 R=0.84 SA=250002 SB=250003 A=0.21 P=1.84 MULT=1
MM1013 N_VPWR_M1013_d N_A_1138_81#_M1013_g A_1096_491# N_VPB_M1014_b PHV L=0.5
+ W=0.42 AD=0.0933154 AS=0.0441 PD=0.822051 PS=0.63 NRD=54.5687 NRS=22.729 M=1
+ R=0.84 SA=250003 SB=250003 A=0.21 P=1.84 MULT=1
MM1011 N_A_1138_81#_M1011_d N_A_917_107#_M1011_g N_VPWR_M1013_d N_VPB_M1014_b
+ PHV L=0.5 W=0.75 AD=0.105 AS=0.166635 PD=1.03 PS=1.46795 NRD=0 NRS=0 M=1 R=1.5
+ SA=250002 SB=250002 A=0.375 P=2.5 MULT=1
MM1002 N_VPWR_M1002_d N_RESET_B_M1002_g N_A_1138_81#_M1011_d N_VPB_M1014_b PHV
+ L=0.5 W=0.75 AD=0.17 AS=0.105 PD=1.26333 PS=1.03 NRD=29.2803 NRS=0 M=1 R=1.5
+ SA=250003 SB=250001 A=0.375 P=2.5 MULT=1
MM1017 N_Q_M1017_d N_A_1138_81#_M1017_g N_VPWR_M1002_d N_VPB_M1014_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.34 PD=3.57 PS=2.52667 NRD=0 NRS=0 M=1 R=3 SA=250002
+ SB=250000 A=0.75 P=4 MULT=1
DX20_noxref N_VNB_M1019_b N_VPB_M1014_b NWDIODE A=26.676 P=25.72
*
.include "sky130_fd_sc_hvl__dlrtp_1.pxi.spice"
*
.ends
*
*
