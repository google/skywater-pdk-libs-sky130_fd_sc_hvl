* File: sky130_fd_sc_hvl__schmittbuf_1.spice
* Created: Fri Aug 28 09:39:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__schmittbuf_1.pex.spice"
.subckt sky130_fd_sc_hvl__schmittbuf_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_A_217_207#_M1001_d N_A_117_181#_M1001_g N_A_64_207#_M1001_s
+ N_VNB_M1001_b NHV L=0.5 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1007 N_A_217_207#_M1007_d N_A_M1007_g N_A_117_181#_M1007_s N_VNB_M1001_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_217_207#_M1007_d N_VNB_M1001_b NHV L=0.5
+ W=0.42 AD=0.328132 AS=0.0588 PD=1.63685 PS=0.7 NRD=21.7056 NRS=0 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1000 N_X_M1000_d N_A_117_181#_M1000_g N_VGND_M1003_d N_VNB_M1001_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.58595 PD=2.03 PS=2.92295 NRD=0 NRS=0 M=1 R=1.5
+ SA=250002 SB=250000 A=0.375 P=2.5 MULT=1
MM1006 N_A_231_463#_M1006_d N_A_117_181#_M1006_g N_A_78_463#_M1006_s
+ N_VPB_M1006_b PHV L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0
+ NRS=0 M=1 R=1.5 SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1005 N_A_231_463#_M1005_d N_A_M1005_g N_A_117_181#_M1005_s N_VPB_M1006_b PHV
+ L=0.5 W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250002 A=0.375 P=2.5 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_231_463#_M1005_d N_VPB_M1006_b PHV L=0.5
+ W=0.75 AD=0.433716 AS=0.105 PD=2.44488 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250001
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1004 N_X_M1004_d N_A_117_181#_M1004_g N_VPWR_M1002_d N_VPB_M1006_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.867431 PD=3.53 PS=4.88976 NRD=0 NRS=0 M=1 R=3 SA=250002
+ SB=250000 A=0.75 P=4 MULT=1
DX8_noxref N_VNB_M1001_b N_A_78_463#_X8_noxref_D1 NDIODE_H A=0.2552 P=2.05
DX9_noxref N_A_64_207#_X9_noxref_D0 N_VPB_M1006_b PDIODE_H A=0.5104 P=3.81
DX10_noxref N_VNB_M1001_b N_VPB_M1006_b NWDIODE A=15.2149 P=17.26
R0 N_A_78_463#_X8_noxref_D1 N_VGND_M1003_d MRDN_HV M=1 w=0.29 l=1.355 
R1 N_A_64_207#_X9_noxref_D0 N_VPWR_M1002_d MRDP_HV M=1 w=0.29 l=3.11 
*
.include "sky130_fd_sc_hvl__schmittbuf_1.pxi.spice"
*
.ends
*
*
