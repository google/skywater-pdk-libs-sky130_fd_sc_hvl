* File: sky130_fd_sc_hvl__sdfstp_1.spice
* Created: Fri Aug 28 09:40:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__sdfstp_1.pex.spice"
.subckt sky130_fd_sc_hvl__sdfstp_1  VNB VPB SCE D SCD CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1031 N_VGND_M1031_d N_SCE_M1031_g N_A_30_107#_M1031_s N_VNB_M1031_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250004 A=0.21 P=1.84 MULT=1
MM1006 A_339_107# N_D_M1006_g N_VGND_M1031_d N_VNB_M1031_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84 SA=250001
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1007 N_A_481_107#_M1007_d N_A_30_107#_M1007_g A_339_107# N_VNB_M1031_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1039 A_637_107# N_SCE_M1039_g N_A_481_107#_M1007_d N_VNB_M1031_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1001 N_VGND_M1001_d N_SCD_M1001_g A_637_107# N_VNB_M1031_b NHV L=0.5 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250003
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1028 N_A_935_107#_M1028_d N_CLK_M1028_g N_VGND_M1001_d N_VNB_M1031_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250004
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1002 N_A_1201_123#_M1002_d N_A_935_107#_M1002_g N_VGND_M1002_s N_VNB_M1031_b
+ NHV L=0.5 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1034 N_A_1471_113#_M1034_d N_A_935_107#_M1034_g N_A_481_107#_M1034_s
+ N_VNB_M1031_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1024 A_1627_113# N_A_1201_123#_M1024_g N_A_1471_113#_M1034_d N_VNB_M1031_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1025 N_VGND_M1025_d N_A_1669_87#_M1025_g A_1627_113# N_VNB_M1031_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1022 A_2035_107# N_A_1471_113#_M1022_g N_A_1669_87#_M1022_s N_VNB_M1031_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250000 SB=250003 A=0.21 P=1.84 MULT=1
MM1010 N_VGND_M1010_d N_SET_B_M1010_g A_2035_107# N_VNB_M1031_b NHV L=0.5 W=0.42
+ AD=0.0879308 AS=0.0441 PD=0.807692 PS=0.63 NRD=25.7754 NRS=13.566 M=1 R=0.84
+ SA=250001 SB=250002 A=0.21 P=1.84 MULT=1
MM1011 A_2352_107# N_A_1471_113#_M1011_g N_VGND_M1010_d N_VNB_M1031_b NHV L=0.5
+ W=0.75 AD=0.07875 AS=0.157019 PD=0.96 PS=1.44231 NRD=7.5924 NRS=0 M=1 R=1.5
+ SA=250001 SB=250003 A=0.375 P=2.5 MULT=1
MM1013 N_A_2477_543#_M1013_d N_A_1201_123#_M1013_g A_2352_107# N_VNB_M1031_b NHV
+ L=0.5 W=0.75 AD=0.157019 AS=0.07875 PD=1.44231 PS=0.96 NRD=0 NRS=7.5924 M=1
+ R=1.5 SA=250002 SB=250002 A=0.375 P=2.5 MULT=1
MM1036 A_2669_173# N_A_935_107#_M1036_g N_A_2477_543#_M1013_d N_VNB_M1031_b NHV
+ L=0.5 W=0.42 AD=0.04515 AS=0.0879308 PD=0.635 PS=0.807692 NRD=14.2386
+ NRS=25.7754 M=1 R=0.84 SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1014 A_2812_173# N_A_2698_421#_M1014_g A_2669_173# N_VNB_M1031_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.04515 PD=0.63 PS=0.635 NRD=13.566 NRS=14.2386 M=1 R=0.84
+ SA=250003 SB=250002 A=0.21 P=1.84 MULT=1
MM1015 N_VGND_M1015_d N_SET_B_M1015_g A_2812_173# N_VNB_M1031_b NHV L=0.5 W=0.42
+ AD=0.09345 AS=0.0441 PD=0.865 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250003
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1023 N_A_2698_421#_M1023_d N_A_2477_543#_M1023_g N_VGND_M1015_d N_VNB_M1031_b
+ NHV L=0.5 W=0.42 AD=0.1197 AS=0.09345 PD=1.41 PS=0.865 NRD=0 NRS=44.7792 M=1
+ R=0.84 SA=250004 SB=250000 A=0.21 P=1.84 MULT=1
MM1032 N_VGND_M1032_d N_A_2477_543#_M1032_g N_A_3321_173#_M1032_s N_VNB_M1031_b
+ NHV L=0.5 W=0.42 AD=0.0933154 AS=0.1197 PD=0.822051 PS=1.41 NRD=31.2132 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1003 N_Q_M1003_d N_A_3321_173#_M1003_g N_VGND_M1032_d N_VNB_M1031_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.166635 PD=2.07 PS=1.46795 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1012 N_VPWR_M1012_d N_SCE_M1012_g N_A_30_107#_M1012_s N_VPB_M1012_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250004 A=0.21 P=1.84 MULT=1
MM1029 A_339_569# N_SCE_M1029_g N_VPWR_M1012_d N_VPB_M1012_b PHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84 SA=250001
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1030 N_A_481_107#_M1030_d N_D_M1030_g A_339_569# N_VPB_M1012_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1017 A_637_569# N_A_30_107#_M1017_g N_A_481_107#_M1030_d N_VPB_M1012_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1021 N_VPWR_M1021_d N_SCD_M1021_g A_637_569# N_VPB_M1012_b PHV L=0.5 W=0.42
+ AD=0.0933154 AS=0.0441 PD=0.822051 PS=0.63 NRD=52.2958 NRS=22.729 M=1 R=0.84
+ SA=250003 SB=250001 A=0.21 P=1.84 MULT=1
MM1008 N_A_935_107#_M1008_d N_CLK_M1008_g N_VPWR_M1021_d N_VPB_M1012_b PHV L=0.5
+ W=0.75 AD=0.21375 AS=0.166635 PD=2.07 PS=1.46795 NRD=0 NRS=0 M=1 R=1.5
+ SA=250002 SB=250000 A=0.375 P=2.5 MULT=1
MM1037 N_A_1201_123#_M1037_d N_A_935_107#_M1037_g N_VPWR_M1037_s N_VPB_M1012_b
+ PHV L=0.5 W=0.75 AD=0.21375 AS=0.21375 PD=2.07 PS=2.07 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1004 N_A_1471_113#_M1004_d N_A_1201_123#_M1004_g N_A_481_107#_M1004_s
+ N_VPB_M1012_b PHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250007 A=0.21 P=1.84 MULT=1
MM1026 A_1686_543# N_A_935_107#_M1026_g N_A_1471_113#_M1004_d N_VPB_M1012_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250001 SB=250006 A=0.21 P=1.84 MULT=1
MM1000 N_VPWR_M1000_d N_A_1669_87#_M1000_g A_1686_543# N_VPB_M1012_b PHV L=0.5
+ W=0.42 AD=0.0756 AS=0.0441 PD=0.78 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250006 A=0.21 P=1.84 MULT=1
MM1018 N_A_1669_87#_M1018_d N_A_1471_113#_M1018_g N_VPWR_M1000_d N_VPB_M1012_b
+ PHV L=0.5 W=0.42 AD=0.0588 AS=0.0756 PD=0.7 PS=0.78 NRD=0 NRS=36.3664 M=1
+ R=0.84 SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1027 N_VPWR_M1027_d N_SET_B_M1027_g N_A_1669_87#_M1018_d N_VPB_M1012_b PHV
+ L=0.5 W=0.42 AD=0.0979606 AS=0.0588 PD=0.825211 PS=0.7 NRD=81.0413 NRS=0 M=1
+ R=0.84 SA=250003 SB=250004 A=0.21 P=1.84 MULT=1
MM1016 A_2335_543# N_A_1471_113#_M1016_g N_VPWR_M1027_d N_VPB_M1012_b PHV L=0.5
+ W=1 AD=0.105 AS=0.233239 PD=1.21 PS=1.96479 NRD=9.5309 NRS=0 M=1 R=2 SA=250002
+ SB=250002 A=0.5 P=3 MULT=1
MM1019 N_A_2477_543#_M1019_d N_A_935_107#_M1019_g A_2335_543# N_VPB_M1012_b PHV
+ L=0.5 W=1 AD=0.233239 AS=0.105 PD=1.96479 PS=1.21 NRD=0 NRS=9.5309 M=1 R=2
+ SA=250002 SB=250001 A=0.5 P=3 MULT=1
MM1005 A_2656_543# N_A_1201_123#_M1005_g N_A_2477_543#_M1019_d N_VPB_M1012_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0979606 PD=0.63 PS=0.825211 NRD=22.729 NRS=52.2958
+ M=1 R=0.84 SA=250006 SB=250002 A=0.21 P=1.84 MULT=1
MM1009 N_VPWR_M1009_d N_A_2698_421#_M1009_g A_2656_543# N_VPB_M1012_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250006 SB=250001 A=0.21 P=1.84 MULT=1
MM1038 N_A_2477_543#_M1038_d N_SET_B_M1038_g N_VPWR_M1009_d N_VPB_M1012_b PHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250007 SB=250000 A=0.21 P=1.84 MULT=1
MM1020 N_VPWR_M1020_d N_A_2477_543#_M1020_g N_A_2698_421#_M1020_s N_VPB_M1012_b
+ PHV L=0.5 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1033 N_VPWR_M1033_d N_A_2477_543#_M1033_g N_A_3321_173#_M1033_s N_VPB_M1012_b
+ PHV L=0.5 W=0.75 AD=0.148929 AS=0.19875 PD=1.17857 PS=2.03 NRD=24.1806 NRS=0
+ M=1 R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1035 N_Q_M1035_d N_A_3321_173#_M1035_g N_VPWR_M1033_d N_VPB_M1012_b PHV L=0.5
+ W=1 AD=0.265 AS=0.198571 PD=2.53 PS=1.57143 NRD=0 NRS=0 M=1 R=2 SA=250001
+ SB=250000 A=0.5 P=3 MULT=1
DX40_noxref N_VNB_M1031_b N_VPB_M1012_b NWDIODE A=50.388 P=43.96
*
.include "sky130_fd_sc_hvl__sdfstp_1.pxi.spice"
*
.ends
*
*
