# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hvl__dlclkp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN GATE
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.385000 0.940000 2.200000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.630000 0.515000 9.995000 1.215000 ;
        RECT 9.630000 1.895000 9.995000 3.735000 ;
        RECT 9.725000 1.215000 9.995000 1.895000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  1.170000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.360000 1.465000 3.690000 1.975000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 10.080000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 10.080000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 10.080000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 10.080000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.985000 10.080000 4.155000 ;
      RECT 0.110000  2.200000  0.440000 3.445000 ;
      RECT 0.110000  3.445000  1.025000 3.555000 ;
      RECT 0.110000  3.555000  3.330000 3.815000 ;
      RECT 0.140000  0.365000  0.765000 0.625000 ;
      RECT 0.140000  0.625000  0.470000 1.170000 ;
      RECT 1.155000  0.365000  2.810000 0.535000 ;
      RECT 1.155000  0.535000  1.865000 0.670000 ;
      RECT 1.195000  3.165000  2.495000 3.385000 ;
      RECT 1.595000  1.555000  2.105000 1.885000 ;
      RECT 1.670000  0.840000  2.000000 1.555000 ;
      RECT 1.670000  1.885000  2.000000 2.995000 ;
      RECT 2.220000  0.705000  2.470000 1.080000 ;
      RECT 2.275000  1.080000  2.470000 2.145000 ;
      RECT 2.275000  2.145000  3.690000 2.315000 ;
      RECT 2.275000  2.315000  2.495000 3.165000 ;
      RECT 2.640000  0.535000  2.810000 1.125000 ;
      RECT 2.640000  1.125000  4.070000 1.295000 ;
      RECT 2.640000  1.295000  2.970000 1.965000 ;
      RECT 2.665000  3.445000  3.330000 3.555000 ;
      RECT 2.980000  0.255000  3.925000 0.535000 ;
      RECT 2.980000  0.535000  3.650000 0.625000 ;
      RECT 2.980000  0.625000  3.330000 0.955000 ;
      RECT 3.000000  2.485000  3.330000 3.445000 ;
      RECT 3.520000  2.315000  3.690000 3.385000 ;
      RECT 3.520000  3.385000  5.515000 3.555000 ;
      RECT 3.820000  0.705000  4.070000 1.125000 ;
      RECT 3.860000  1.295000  4.070000 3.005000 ;
      RECT 3.860000  3.005000  5.175000 3.215000 ;
      RECT 4.095000  0.255000  4.660000 0.535000 ;
      RECT 4.375000  0.535000  4.660000 1.195000 ;
      RECT 4.375000  1.195000  6.490000 1.365000 ;
      RECT 4.375000  1.365000  4.545000 2.330000 ;
      RECT 4.375000  2.330000  4.660000 2.660000 ;
      RECT 4.715000  1.615000  5.305000 1.945000 ;
      RECT 4.830000  0.255000  6.150000 0.625000 ;
      RECT 5.135000  1.945000  5.305000 2.425000 ;
      RECT 5.135000  2.425000  5.515000 2.595000 ;
      RECT 5.345000  2.595000  5.515000 3.385000 ;
      RECT 5.515000  1.535000  5.845000 1.875000 ;
      RECT 5.515000  1.875000  6.930000 2.085000 ;
      RECT 5.685000  3.445000  8.065000 3.615000 ;
      RECT 5.685000  3.615000  9.460000 3.815000 ;
      RECT 5.820000  0.625000  6.150000 1.025000 ;
      RECT 5.820000  2.330000  6.150000 3.445000 ;
      RECT 6.125000  1.365000  6.490000 1.655000 ;
      RECT 6.320000  0.355000  6.910000 0.670000 ;
      RECT 6.320000  0.670000  6.490000 1.195000 ;
      RECT 6.660000  0.840000  6.930000 1.615000 ;
      RECT 6.660000  1.615000  7.785000 1.825000 ;
      RECT 6.660000  1.825000  6.930000 1.875000 ;
      RECT 6.660000  2.085000  6.930000 2.660000 ;
      RECT 7.080000  0.255000  9.460000 0.625000 ;
      RECT 7.150000  0.885000  8.180000 1.215000 ;
      RECT 7.150000  2.225000  7.480000 3.445000 ;
      RECT 7.455000  1.385000  7.785000 1.615000 ;
      RECT 7.455000  1.825000  7.785000 2.055000 ;
      RECT 7.955000  1.215000  8.180000 1.385000 ;
      RECT 7.955000  1.385000  9.555000 1.555000 ;
      RECT 7.955000  1.555000  8.180000 2.955000 ;
      RECT 8.235000  3.125000  8.600000 3.445000 ;
      RECT 8.350000  1.725000  8.680000 2.025000 ;
      RECT 8.350000  2.025000  8.600000 3.125000 ;
      RECT 8.770000  0.625000  9.100000 1.215000 ;
      RECT 8.770000  2.195000  9.100000 3.445000 ;
      RECT 8.770000  3.445000  9.460000 3.615000 ;
      RECT 8.945000  1.555000  9.555000 1.725000 ;
    LAYER mcon ;
      RECT 0.140000  3.475000 0.310000 3.645000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.175000  0.425000 0.345000 0.595000 ;
      RECT 0.500000  3.475000 0.670000 3.645000 ;
      RECT 0.535000  0.425000 0.705000 0.595000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.860000  3.600000 1.030000 3.770000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.220000  3.600000 1.390000 3.770000 ;
      RECT 1.580000  3.600000 1.750000 3.770000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.995000  3.600000 2.165000 3.770000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.355000  3.600000 2.525000 3.770000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.715000  3.475000 2.885000 3.645000 ;
      RECT 2.995000  0.425000 3.165000 0.595000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.075000  3.475000 3.245000 3.645000 ;
      RECT 3.355000  0.425000 3.525000 0.595000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.715000  0.355000 3.885000 0.525000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.870000  0.355000 5.040000 0.525000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 5.230000  0.355000 5.400000 0.525000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.985000 5.605000 4.155000 ;
      RECT 5.435000  3.985000 5.605000 4.155000 ;
      RECT 5.590000  0.425000 5.760000 0.595000 ;
      RECT 5.715000  3.475000 5.885000 3.645000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.985000 6.085000 4.155000 ;
      RECT 5.915000  3.985000 6.085000 4.155000 ;
      RECT 5.950000  0.425000 6.120000 0.595000 ;
      RECT 6.075000  3.475000 6.245000 3.645000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.985000 6.565000 4.155000 ;
      RECT 6.395000  3.985000 6.565000 4.155000 ;
      RECT 6.435000  3.545000 6.605000 3.715000 ;
      RECT 6.795000  3.545000 6.965000 3.715000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.985000 7.045000 4.155000 ;
      RECT 6.875000  3.985000 7.045000 4.155000 ;
      RECT 7.100000  0.355000 7.270000 0.525000 ;
      RECT 7.155000  3.475000 7.325000 3.645000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.460000  0.355000 7.630000 0.525000 ;
      RECT 7.515000  3.475000 7.685000 3.645000 ;
      RECT 7.820000  0.355000 7.990000 0.525000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 8.180000  0.355000 8.350000 0.525000 ;
      RECT 8.195000  3.615000 8.365000 3.785000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.985000 8.485000 4.155000 ;
      RECT 8.315000  3.985000 8.485000 4.155000 ;
      RECT 8.540000  0.425000 8.710000 0.595000 ;
      RECT 8.555000  3.615000 8.725000 3.785000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.985000 8.965000 4.155000 ;
      RECT 8.795000  3.985000 8.965000 4.155000 ;
      RECT 8.900000  0.425000 9.070000 0.595000 ;
      RECT 8.915000  3.475000 9.085000 3.645000 ;
      RECT 9.260000  0.425000 9.430000 0.595000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.475000 9.445000 3.645000 ;
      RECT 9.275000  3.985000 9.445000 4.155000 ;
      RECT 9.275000  3.985000 9.445000 4.155000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.985000 9.925000 4.155000 ;
      RECT 9.755000  3.985000 9.925000 4.155000 ;
  END
END sky130_fd_sc_hvl__dlclkp_1
