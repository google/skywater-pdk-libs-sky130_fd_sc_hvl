* File: sky130_fd_sc_hvl__buf_1.pxi.spice
* Created: Wed Sep  2 09:03:58 2020
* 
x_PM_SKY130_FD_SC_HVL__BUF_1%VNB N_VNB_M1001_b VNB N_VNB_c_5_p VNB
+ PM_SKY130_FD_SC_HVL__BUF_1%VNB
x_PM_SKY130_FD_SC_HVL__BUF_1%VPB N_VPB_M1000_b VPB N_VPB_c_20_p VPB
+ PM_SKY130_FD_SC_HVL__BUF_1%VPB
x_PM_SKY130_FD_SC_HVL__BUF_1%A_84_81# N_A_84_81#_M1002_d N_A_84_81#_M1003_d
+ N_A_84_81#_M1001_g N_A_84_81#_M1000_g N_A_84_81#_c_36_n N_A_84_81#_c_37_n
+ N_A_84_81#_c_38_n N_A_84_81#_c_72_p N_A_84_81#_c_39_n N_A_84_81#_c_41_n
+ N_A_84_81#_c_42_n N_A_84_81#_c_43_n PM_SKY130_FD_SC_HVL__BUF_1%A_84_81#
x_PM_SKY130_FD_SC_HVL__BUF_1%A A A A A A N_A_M1002_g N_A_c_86_n N_A_M1003_g
+ PM_SKY130_FD_SC_HVL__BUF_1%A
x_PM_SKY130_FD_SC_HVL__BUF_1%X N_X_M1001_s N_X_M1000_s X X X X X X X N_X_c_104_n
+ X N_X_c_110_n PM_SKY130_FD_SC_HVL__BUF_1%X
x_PM_SKY130_FD_SC_HVL__BUF_1%VPWR N_VPWR_M1000_d VPWR N_VPWR_c_125_n
+ PM_SKY130_FD_SC_HVL__BUF_1%VPWR
x_PM_SKY130_FD_SC_HVL__BUF_1%VGND N_VGND_M1001_d VGND N_VGND_c_140_n
+ PM_SKY130_FD_SC_HVL__BUF_1%VGND
cc_1 N_VNB_M1001_b N_A_84_81#_c_36_n 0.00140289f $X=-0.33 $Y=-0.265 $X2=0.84
+ $Y2=1.58
cc_2 N_VNB_M1001_b N_A_84_81#_c_37_n 0.0581956f $X=-0.33 $Y=-0.265 $X2=0.84
+ $Y2=1.58
cc_3 N_VNB_M1001_b N_A_84_81#_c_38_n 0.0121633f $X=-0.33 $Y=-0.265 $X2=1.975
+ $Y2=1.2
cc_4 N_VNB_M1001_b N_A_84_81#_c_39_n 0.0310211f $X=-0.33 $Y=-0.265 $X2=2.06
+ $Y2=0.745
cc_5 N_VNB_c_5_p N_A_84_81#_c_39_n 5.81195e-19 $X=0.24 $Y=0 $X2=2.06 $Y2=0.745
cc_6 N_VNB_M1001_b N_A_84_81#_c_41_n 0.030449f $X=-0.33 $Y=-0.265 $X2=2.06
+ $Y2=2.34
cc_7 N_VNB_M1001_b N_A_84_81#_c_42_n 0.00770964f $X=-0.33 $Y=-0.265 $X2=2.1
+ $Y2=1.2
cc_8 N_VNB_M1001_b N_A_84_81#_c_43_n 0.0441687f $X=-0.33 $Y=-0.265 $X2=0.722
+ $Y2=1.395
cc_9 N_VNB_c_5_p N_A_84_81#_c_43_n 5.86481e-19 $X=0.24 $Y=0 $X2=0.722 $Y2=1.395
cc_10 N_VNB_M1001_b N_A_M1002_g 0.128583f $X=-0.33 $Y=-0.265 $X2=0.775 $Y2=2.965
cc_11 N_VNB_c_5_p N_A_M1002_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.775 $Y2=2.965
cc_12 N_VNB_M1001_b N_X_c_104_n 0.0674551f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_13 N_VNB_c_5_p N_X_c_104_n 5.81195e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_14 N_VNB_M1001_b VGND 0.0658643f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_15 N_VNB_c_5_p VGND 0.256669f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_16 N_VNB_M1001_b N_VGND_c_140_n 0.0622807f $X=-0.33 $Y=-0.265 $X2=0.67
+ $Y2=1.395
cc_17 N_VNB_c_5_p N_VGND_c_140_n 0.0035518f $X=0.24 $Y=0 $X2=0.67 $Y2=1.395
cc_18 N_VPB_M1000_b N_A_84_81#_M1000_g 0.061601f $X=-0.33 $Y=1.885 $X2=0.775
+ $Y2=2.965
cc_19 VPB N_A_84_81#_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.775 $Y2=2.965
cc_20 N_VPB_c_20_p N_A_84_81#_M1000_g 0.0158814f $X=2.16 $Y=4.07 $X2=0.775
+ $Y2=2.965
cc_21 N_VPB_M1000_b N_A_84_81#_c_37_n 0.00408238f $X=-0.33 $Y=1.885 $X2=0.84
+ $Y2=1.58
cc_22 N_VPB_M1000_b N_A_84_81#_c_41_n 0.050803f $X=-0.33 $Y=1.885 $X2=2.06
+ $Y2=2.34
cc_23 N_VPB_M1000_b N_A_M1002_g 0.0652915f $X=-0.33 $Y=1.885 $X2=0.775 $Y2=2.965
cc_24 N_VPB_M1000_b N_A_c_86_n 0.0116704f $X=-0.33 $Y=1.885 $X2=0.84 $Y2=1.58
cc_25 N_VPB_M1000_b N_X_c_104_n 0.0158198f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_26 N_VPB_M1000_b X 0.0527822f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_27 VPB X 0.00136875f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_28 N_VPB_c_20_p X 0.0227858f $X=2.16 $Y=4.07 $X2=0 $Y2=0
cc_29 N_VPB_M1000_b N_X_c_110_n 0.0130587f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_30 N_VPB_M1000_b VPWR 0.0721634f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_31 VPB VPWR 0.255897f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_32 N_VPB_c_20_p VPWR 0.0142003f $X=2.16 $Y=4.07 $X2=0 $Y2=0
cc_33 N_VPB_M1000_b N_VPWR_c_125_n 0.0127017f $X=-0.33 $Y=1.885 $X2=0.67
+ $Y2=1.395
cc_34 VPB N_VPWR_c_125_n 0.00220475f $X=0 $Y=3.955 $X2=0.67 $Y2=1.395
cc_35 N_VPB_c_20_p N_VPWR_c_125_n 0.0280583f $X=2.16 $Y=4.07 $X2=0.67 $Y2=1.395
cc_36 N_A_84_81#_c_36_n N_A_M1002_g 0.00392032f $X=0.84 $Y=1.58 $X2=0 $Y2=0
cc_37 N_A_84_81#_c_37_n N_A_M1002_g 0.0408226f $X=0.84 $Y=1.58 $X2=0 $Y2=0
cc_38 N_A_84_81#_c_38_n N_A_M1002_g 0.034515f $X=1.975 $Y=1.2 $X2=0 $Y2=0
cc_39 N_A_84_81#_c_39_n N_A_M1002_g 0.0090774f $X=2.06 $Y=0.745 $X2=0 $Y2=0
cc_40 N_A_84_81#_c_41_n N_A_M1002_g 0.0335927f $X=2.06 $Y=2.34 $X2=0 $Y2=0
cc_41 N_A_84_81#_c_43_n N_A_M1002_g 0.0184277f $X=0.722 $Y=1.395 $X2=0 $Y2=0
cc_42 N_A_84_81#_M1000_g N_A_c_86_n 3.02269e-19 $X=0.775 $Y=2.965 $X2=2.16 $Y2=0
cc_43 N_A_84_81#_c_36_n N_A_c_86_n 0.00936991f $X=0.84 $Y=1.58 $X2=2.16 $Y2=0
cc_44 N_A_84_81#_c_37_n N_A_c_86_n 0.00392409f $X=0.84 $Y=1.58 $X2=2.16 $Y2=0
cc_45 N_A_84_81#_c_38_n N_A_c_86_n 0.0238596f $X=1.975 $Y=1.2 $X2=2.16 $Y2=0
cc_46 N_A_84_81#_c_41_n N_A_c_86_n 0.0853873f $X=2.06 $Y=2.34 $X2=2.16 $Y2=0
cc_47 N_A_84_81#_M1000_g N_X_c_104_n 0.0116165f $X=0.775 $Y=2.965 $X2=1.2
+ $Y2=0.058
cc_48 N_A_84_81#_c_36_n N_X_c_104_n 0.0226758f $X=0.84 $Y=1.58 $X2=1.2 $Y2=0.058
cc_49 N_A_84_81#_c_43_n N_X_c_104_n 0.0242663f $X=0.722 $Y=1.395 $X2=1.2
+ $Y2=0.058
cc_50 N_A_84_81#_M1000_g X 0.0235663f $X=0.775 $Y=2.965 $X2=0 $Y2=0
cc_51 N_A_84_81#_M1000_g N_X_c_110_n 0.00574889f $X=0.775 $Y=2.965 $X2=0 $Y2=0
cc_52 N_A_84_81#_c_37_n N_X_c_110_n 0.0045161f $X=0.84 $Y=1.58 $X2=0 $Y2=0
cc_53 N_A_84_81#_M1000_g VPWR 0.0112082f $X=0.775 $Y=2.965 $X2=0 $Y2=0
cc_54 N_A_84_81#_c_41_n VPWR 0.0109527f $X=2.06 $Y=2.34 $X2=0 $Y2=0
cc_55 N_A_84_81#_M1000_g N_VPWR_c_125_n 0.0763398f $X=0.775 $Y=2.965 $X2=0 $Y2=0
cc_56 N_A_84_81#_c_36_n N_VPWR_c_125_n 0.0107918f $X=0.84 $Y=1.58 $X2=0 $Y2=0
cc_57 N_A_84_81#_c_38_n N_VGND_M1001_d 0.00985042f $X=1.975 $Y=1.2 $X2=0 $Y2=0
cc_58 N_A_84_81#_c_72_p N_VGND_M1001_d 2.97932e-19 $X=1.005 $Y=1.2 $X2=0 $Y2=0
cc_59 N_A_84_81#_M1002_d VGND 6.76135e-19 $X=1.92 $Y=0.535 $X2=0 $Y2=0
cc_60 N_A_84_81#_c_38_n VGND 0.008626f $X=1.975 $Y=1.2 $X2=0 $Y2=0
cc_61 N_A_84_81#_c_72_p VGND 0.00135661f $X=1.005 $Y=1.2 $X2=0 $Y2=0
cc_62 N_A_84_81#_c_39_n VGND 0.0266128f $X=2.06 $Y=0.745 $X2=0 $Y2=0
cc_63 N_A_84_81#_c_43_n VGND 0.00869985f $X=0.722 $Y=1.395 $X2=0 $Y2=0
cc_64 N_A_84_81#_c_37_n N_VGND_c_140_n 3.04803e-19 $X=0.84 $Y=1.58 $X2=0 $Y2=0
cc_65 N_A_84_81#_c_38_n N_VGND_c_140_n 0.0543159f $X=1.975 $Y=1.2 $X2=0 $Y2=0
cc_66 N_A_84_81#_c_72_p N_VGND_c_140_n 0.0208495f $X=1.005 $Y=1.2 $X2=0 $Y2=0
cc_67 N_A_84_81#_c_39_n N_VGND_c_140_n 0.0192683f $X=2.06 $Y=0.745 $X2=0 $Y2=0
cc_68 N_A_84_81#_c_43_n N_VGND_c_140_n 0.0421821f $X=0.722 $Y=1.395 $X2=0 $Y2=0
cc_69 N_A_M1002_g VPWR 0.0048774f $X=1.67 $Y=0.745 $X2=0 $Y2=0
cc_70 N_A_c_86_n VPWR 0.0185236f $X=1.63 $Y=1.55 $X2=0 $Y2=0
cc_71 N_A_M1002_g N_VPWR_c_125_n 0.00883995f $X=1.67 $Y=0.745 $X2=0 $Y2=0
cc_72 N_A_c_86_n N_VPWR_c_125_n 0.0847009f $X=1.63 $Y=1.55 $X2=0 $Y2=0
cc_73 N_A_M1002_g VGND 0.00513207f $X=1.67 $Y=0.745 $X2=0 $Y2=0
cc_74 N_A_M1002_g N_VGND_c_140_n 0.0443101f $X=1.67 $Y=0.745 $X2=0 $Y2=0
cc_75 X VPWR 0.053097f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_76 N_X_c_110_n N_VPWR_c_125_n 0.115775f $X=0.385 $Y=2.34 $X2=0 $Y2=0
cc_77 N_X_M1001_s VGND 0.00221032f $X=0.155 $Y=0.535 $X2=0 $Y2=0
cc_78 N_X_c_104_n VGND 0.026283f $X=0.28 $Y=0.68 $X2=0 $Y2=0
cc_79 N_X_c_104_n N_VGND_c_140_n 0.0192683f $X=0.28 $Y=0.68 $X2=0 $Y2=0
