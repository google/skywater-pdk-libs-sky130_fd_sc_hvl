* File: sky130_fd_sc_hvl__mux4_1.pxi.spice
* Created: Fri Aug 28 09:37:49 2020
* 
x_PM_SKY130_FD_SC_HVL__MUX4_1%VNB N_VNB_M1020_b VNB N_VNB_c_3_p VNB
+ PM_SKY130_FD_SC_HVL__MUX4_1%VNB
x_PM_SKY130_FD_SC_HVL__MUX4_1%VPB N_VPB_M1013_b VPB N_VPB_c_95_p VPB
+ PM_SKY130_FD_SC_HVL__MUX4_1%VPB
x_PM_SKY130_FD_SC_HVL__MUX4_1%S0 N_S0_c_230_n N_S0_M1023_g N_S0_M1012_g
+ N_S0_c_217_n N_S0_M1018_g N_S0_M1025_g N_S0_c_237_n N_S0_c_238_n N_S0_c_252_p
+ N_S0_c_239_n N_S0_c_242_n N_S0_c_220_n N_S0_c_221_n N_S0_c_222_n N_S0_c_223_n
+ N_S0_c_265_p N_S0_c_253_p N_S0_c_246_n S0 S0 S0 N_S0_M1020_g N_S0_M1013_g
+ N_S0_c_227_n N_S0_c_228_n N_S0_c_229_n PM_SKY130_FD_SC_HVL__MUX4_1%S0
x_PM_SKY130_FD_SC_HVL__MUX4_1%A2 N_A2_c_390_n N_A2_M1006_g N_A2_M1000_g
+ N_A2_c_399_n A2 A2 N_A2_c_394_n PM_SKY130_FD_SC_HVL__MUX4_1%A2
x_PM_SKY130_FD_SC_HVL__MUX4_1%A_30_107# N_A_30_107#_M1020_s N_A_30_107#_M1013_s
+ N_A_30_107#_M1016_g N_A_30_107#_M1001_g N_A_30_107#_c_429_n
+ N_A_30_107#_c_431_n N_A_30_107#_c_465_n N_A_30_107#_c_445_n
+ N_A_30_107#_c_446_n N_A_30_107#_c_447_n N_A_30_107#_c_448_n
+ N_A_30_107#_c_432_n N_A_30_107#_c_433_n N_A_30_107#_c_450_n
+ N_A_30_107#_c_434_n N_A_30_107#_c_483_n N_A_30_107#_c_454_n
+ N_A_30_107#_M1007_g N_A_30_107#_M1021_g N_A_30_107#_c_438_n
+ PM_SKY130_FD_SC_HVL__MUX4_1%A_30_107#
x_PM_SKY130_FD_SC_HVL__MUX4_1%A3 N_A3_M1002_g N_A3_M1009_g N_A3_c_572_n A3 A3
+ N_A3_c_577_n N_A3_c_573_n PM_SKY130_FD_SC_HVL__MUX4_1%A3
x_PM_SKY130_FD_SC_HVL__MUX4_1%A1 N_A1_M1004_g N_A1_c_620_n A1 A1 A1 N_A1_c_621_n
+ N_A1_M1024_g PM_SKY130_FD_SC_HVL__MUX4_1%A1
x_PM_SKY130_FD_SC_HVL__MUX4_1%A0 N_A0_M1019_g N_A0_M1008_g N_A0_c_666_n
+ N_A0_c_662_n A0 A0 A0 N_A0_c_663_n PM_SKY130_FD_SC_HVL__MUX4_1%A0
x_PM_SKY130_FD_SC_HVL__MUX4_1%S1 N_S1_M1003_g N_S1_c_704_n N_S1_M1005_g
+ N_S1_c_706_n N_S1_c_707_n N_S1_M1010_g N_S1_M1014_g N_S1_c_708_n N_S1_c_716_n
+ N_S1_c_717_n N_S1_c_723_p N_S1_c_718_n N_S1_c_742_p S1 S1 S1 N_S1_c_720_n
+ PM_SKY130_FD_SC_HVL__MUX4_1%S1
x_PM_SKY130_FD_SC_HVL__MUX4_1%A_1681_89# N_A_1681_89#_M1010_s
+ N_A_1681_89#_M1014_s N_A_1681_89#_c_791_n N_A_1681_89#_M1017_g
+ N_A_1681_89#_M1011_g N_A_1681_89#_c_798_n N_A_1681_89#_c_794_n
+ N_A_1681_89#_c_800_n N_A_1681_89#_c_801_n
+ PM_SKY130_FD_SC_HVL__MUX4_1%A_1681_89#
x_PM_SKY130_FD_SC_HVL__MUX4_1%A_1669_615# N_A_1669_615#_M1011_d
+ N_A_1669_615#_M1003_d N_A_1669_615#_c_867_n N_A_1669_615#_c_868_n
+ N_A_1669_615#_c_871_n N_A_1669_615#_c_882_n N_A_1669_615#_c_859_n
+ N_A_1669_615#_c_861_n N_A_1669_615#_c_863_n N_A_1669_615#_c_874_n
+ N_A_1669_615#_c_864_n N_A_1669_615#_c_890_n N_A_1669_615#_M1022_g
+ N_A_1669_615#_M1015_g PM_SKY130_FD_SC_HVL__MUX4_1%A_1669_615#
x_PM_SKY130_FD_SC_HVL__MUX4_1%VPWR N_VPWR_M1013_d N_VPWR_M1009_d N_VPWR_M1019_d
+ N_VPWR_M1014_d VPWR N_VPWR_c_931_n N_VPWR_c_934_n N_VPWR_c_937_n
+ N_VPWR_c_940_n N_VPWR_c_943_n PM_SKY130_FD_SC_HVL__MUX4_1%VPWR
x_PM_SKY130_FD_SC_HVL__MUX4_1%A_481_107# N_A_481_107#_M1007_d
+ N_A_481_107#_M1005_d N_A_481_107#_M1023_d N_A_481_107#_M1017_d
+ N_A_481_107#_c_1027_n N_A_481_107#_c_1029_n N_A_481_107#_c_1030_n
+ N_A_481_107#_c_1031_n N_A_481_107#_c_1032_n N_A_481_107#_c_1034_n
+ N_A_481_107#_c_1087_n N_A_481_107#_c_1036_n N_A_481_107#_c_1105_n
+ N_A_481_107#_c_1037_n N_A_481_107#_c_1038_n N_A_481_107#_c_1040_n
+ N_A_481_107#_c_1108_n N_A_481_107#_c_1042_n N_A_481_107#_c_1043_n
+ N_A_481_107#_c_1044_n N_A_481_107#_c_1045_n N_A_481_107#_c_1046_n
+ N_A_481_107#_c_1071_n N_A_481_107#_c_1049_n
+ PM_SKY130_FD_SC_HVL__MUX4_1%A_481_107#
x_PM_SKY130_FD_SC_HVL__MUX4_1%A_1097_627# N_A_1097_627#_M1012_d
+ N_A_1097_627#_M1011_s N_A_1097_627#_M1001_d N_A_1097_627#_M1003_s
+ N_A_1097_627#_c_1190_n N_A_1097_627#_c_1191_n N_A_1097_627#_c_1209_n
+ N_A_1097_627#_c_1194_n N_A_1097_627#_c_1195_n N_A_1097_627#_c_1185_n
+ N_A_1097_627#_c_1197_n N_A_1097_627#_c_1186_n N_A_1097_627#_c_1199_n
+ N_A_1097_627#_c_1187_n N_A_1097_627#_c_1188_n N_A_1097_627#_c_1189_n
+ N_A_1097_627#_c_1200_n N_A_1097_627#_c_1201_n N_A_1097_627#_c_1202_n
+ N_A_1097_627#_c_1203_n PM_SKY130_FD_SC_HVL__MUX4_1%A_1097_627#
x_PM_SKY130_FD_SC_HVL__MUX4_1%X N_X_M1022_d N_X_M1015_d X X X X X X X
+ N_X_c_1296_n PM_SKY130_FD_SC_HVL__MUX4_1%X
x_PM_SKY130_FD_SC_HVL__MUX4_1%VGND N_VGND_M1020_d N_VGND_M1002_d N_VGND_M1008_d
+ N_VGND_M1010_d VGND N_VGND_c_1309_n N_VGND_c_1311_n N_VGND_c_1313_n
+ N_VGND_c_1315_n N_VGND_c_1317_n PM_SKY130_FD_SC_HVL__MUX4_1%VGND
cc_1 N_VNB_M1020_b N_S0_c_217_n 0.0493192f $X=-0.33 $Y=-0.265 $X2=5.41 $Y2=1.945
cc_2 N_VNB_M1020_b N_S0_M1025_g 0.0497677f $X=-0.33 $Y=-0.265 $X2=2.935
+ $Y2=0.745
cc_3 N_VNB_c_3_p N_S0_M1025_g 0.00232707f $X=0.24 $Y=0 $X2=2.935 $Y2=0.745
cc_4 N_VNB_M1020_b N_S0_c_220_n 0.00239223f $X=-0.33 $Y=-0.265 $X2=2.77 $Y2=2.8
cc_5 N_VNB_M1020_b N_S0_c_221_n 0.0140194f $X=-0.33 $Y=-0.265 $X2=4.925
+ $Y2=1.607
cc_6 N_VNB_M1020_b N_S0_c_222_n 0.00222112f $X=-0.33 $Y=-0.265 $X2=2.855
+ $Y2=1.607
cc_7 N_VNB_M1020_b N_S0_c_223_n 0.0531147f $X=-0.33 $Y=-0.265 $X2=2.87 $Y2=1.53
cc_8 N_VNB_M1020_b S0 0.00444456f $X=-0.33 $Y=-0.265 $X2=4.955 $Y2=0.84
cc_9 N_VNB_M1020_b N_S0_M1020_g 0.125986f $X=-0.33 $Y=-0.265 $X2=0.665 $Y2=0.745
cc_10 N_VNB_c_3_p N_S0_M1020_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=0.745
cc_11 N_VNB_M1020_b N_S0_c_227_n 0.02677f $X=-0.33 $Y=-0.265 $X2=5.31 $Y2=1.265
cc_12 N_VNB_M1020_b N_S0_c_228_n 0.0367878f $X=-0.33 $Y=-0.265 $X2=5.41 $Y2=1.08
cc_13 N_VNB_M1020_b N_S0_c_229_n 0.00162672f $X=-0.33 $Y=-0.265 $X2=5.172
+ $Y2=1.445
cc_14 N_VNB_M1020_b N_A2_c_390_n 0.0118295f $X=-0.33 $Y=-0.265 $X2=2.155
+ $Y2=3.345
cc_15 N_VNB_M1020_b N_A2_M1006_g 0.0742064f $X=-0.33 $Y=-0.265 $X2=5.375
+ $Y2=1.08
cc_16 N_VNB_c_3_p N_A2_M1006_g 5.86481e-19 $X=0.24 $Y=0 $X2=5.375 $Y2=1.08
cc_17 N_VNB_M1020_b A2 0.00462717f $X=-0.33 $Y=-0.265 $X2=6.015 $Y2=3.345
cc_18 N_VNB_M1020_b N_A2_c_394_n 0.0236216f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_19 N_VNB_M1020_b N_A_30_107#_c_429_n 0.0343513f $X=-0.33 $Y=-0.265 $X2=2.935
+ $Y2=1.085
cc_20 N_VNB_c_3_p N_A_30_107#_c_429_n 7.98897e-19 $X=0.24 $Y=0 $X2=2.935
+ $Y2=1.085
cc_21 N_VNB_M1020_b N_A_30_107#_c_431_n 0.0198941f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_22 N_VNB_M1020_b N_A_30_107#_c_432_n 0.00259179f $X=-0.33 $Y=-0.265 $X2=2.07
+ $Y2=2.47
cc_23 N_VNB_M1020_b N_A_30_107#_c_433_n 0.0132078f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_24 N_VNB_M1020_b N_A_30_107#_c_434_n 0.0264882f $X=-0.33 $Y=-0.265 $X2=4.955
+ $Y2=0.84
cc_25 N_VNB_M1020_b N_A_30_107#_M1007_g 0.0870979f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_26 N_VNB_c_3_p N_A_30_107#_M1007_g 0.0023273f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_27 N_VNB_M1020_b N_A_30_107#_M1021_g 0.106098f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_28 N_VNB_M1020_b N_A_30_107#_c_438_n 0.0356765f $X=-0.33 $Y=-0.265 $X2=5.41
+ $Y2=1.08
cc_29 N_VNB_M1020_b N_A3_M1002_g 0.0402114f $X=-0.33 $Y=-0.265 $X2=2.155
+ $Y2=3.345
cc_30 N_VNB_M1020_b N_A3_c_572_n 0.0540662f $X=-0.33 $Y=-0.265 $X2=6.015
+ $Y2=3.345
cc_31 N_VNB_M1020_b N_A3_c_573_n 0.028138f $X=-0.33 $Y=-0.265 $X2=6.015 $Y2=2.37
cc_32 N_VNB_M1020_b N_A1_M1004_g 0.0389975f $X=-0.33 $Y=-0.265 $X2=2.155
+ $Y2=3.345
cc_33 N_VNB_M1020_b N_A1_c_620_n 0.0580703f $X=-0.33 $Y=-0.265 $X2=5.375
+ $Y2=0.745
cc_34 N_VNB_M1020_b N_A1_c_621_n 0.0257569f $X=-0.33 $Y=-0.265 $X2=2.935
+ $Y2=0.745
cc_35 N_VNB_M1020_b N_A0_M1008_g 0.0480357f $X=-0.33 $Y=-0.265 $X2=5.375
+ $Y2=0.745
cc_36 N_VNB_c_3_p N_A0_M1008_g 8.30748e-19 $X=0.24 $Y=0 $X2=5.375 $Y2=0.745
cc_37 N_VNB_M1020_b N_A0_c_662_n 0.0285651f $X=-0.33 $Y=-0.265 $X2=6.015
+ $Y2=3.345
cc_38 N_VNB_M1020_b N_A0_c_663_n 0.0606272f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_39 N_VNB_M1020_b N_S1_c_704_n 0.053006f $X=-0.33 $Y=-0.265 $X2=5.375 $Y2=1.08
cc_40 N_VNB_M1020_b N_S1_M1005_g 0.0598177f $X=-0.33 $Y=-0.265 $X2=5.375
+ $Y2=0.745
cc_41 N_VNB_M1020_b N_S1_c_706_n 0.0653911f $X=-0.33 $Y=-0.265 $X2=5.41
+ $Y2=1.945
cc_42 N_VNB_M1020_b N_S1_c_707_n 0.0409344f $X=-0.33 $Y=-0.265 $X2=6.015
+ $Y2=3.345
cc_43 N_VNB_M1020_b N_S1_c_708_n 0.0300327f $X=-0.33 $Y=-0.265 $X2=2.935
+ $Y2=1.085
cc_44 N_VNB_M1020_b N_A_1681_89#_c_791_n 0.0584772f $X=-0.33 $Y=-0.265 $X2=5.41
+ $Y2=1.365
cc_45 N_VNB_M1020_b N_A_1681_89#_M1011_g 0.0550252f $X=-0.33 $Y=-0.265 $X2=2.945
+ $Y2=1.085
cc_46 N_VNB_c_3_p N_A_1681_89#_M1011_g 8.10183e-19 $X=0.24 $Y=0 $X2=2.945
+ $Y2=1.085
cc_47 N_VNB_M1020_b N_A_1681_89#_c_794_n 0.0107856f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_M1020_b N_A_1669_615#_c_859_n 0.138306f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_49 N_VNB_c_3_p N_A_1669_615#_c_859_n 0.00559603f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_50 N_VNB_M1020_b N_A_1669_615#_c_861_n 0.024013f $X=-0.33 $Y=-0.265 $X2=2.935
+ $Y2=1.085
cc_51 N_VNB_c_3_p N_A_1669_615#_c_861_n 0.00109845f $X=0.24 $Y=0 $X2=2.935
+ $Y2=1.085
cc_52 N_VNB_M1020_b N_A_1669_615#_c_863_n 0.0128533f $X=-0.33 $Y=-0.265
+ $X2=6.015 $Y2=2.37
cc_53 N_VNB_M1020_b N_A_1669_615#_c_864_n 0.00602302f $X=-0.33 $Y=-0.265
+ $X2=2.03 $Y2=2.5
cc_54 N_VNB_M1020_b N_A_1669_615#_M1022_g 0.0846381f $X=-0.33 $Y=-0.265 $X2=2.77
+ $Y2=2.8
cc_55 N_VNB_c_3_p N_A_1669_615#_M1022_g 5.29412e-19 $X=0.24 $Y=0 $X2=2.77
+ $Y2=2.8
cc_56 N_VNB_M1020_b N_A_481_107#_c_1027_n 0.0120645f $X=-0.33 $Y=-0.265
+ $X2=2.935 $Y2=0.745
cc_57 N_VNB_c_3_p N_A_481_107#_c_1027_n 0.00107308f $X=0.24 $Y=0 $X2=2.935
+ $Y2=0.745
cc_58 N_VNB_M1020_b N_A_481_107#_c_1029_n 0.00508042f $X=-0.33 $Y=-0.265
+ $X2=2.935 $Y2=1.085
cc_59 N_VNB_M1020_b N_A_481_107#_c_1030_n 0.00904915f $X=-0.33 $Y=-0.265
+ $X2=5.41 $Y2=1.945
cc_60 N_VNB_M1020_b N_A_481_107#_c_1031_n 0.00198331f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_61 N_VNB_M1020_b N_A_481_107#_c_1032_n 0.170895f $X=-0.33 $Y=-0.265 $X2=1.905
+ $Y2=2.415
cc_62 N_VNB_c_3_p N_A_481_107#_c_1032_n 0.0080622f $X=0.24 $Y=0 $X2=1.905
+ $Y2=2.415
cc_63 N_VNB_M1020_b N_A_481_107#_c_1034_n 0.0136651f $X=-0.33 $Y=-0.265
+ $X2=0.895 $Y2=2.415
cc_64 N_VNB_c_3_p N_A_481_107#_c_1034_n 5.63772e-19 $X=0.24 $Y=0 $X2=0.895
+ $Y2=2.415
cc_65 N_VNB_M1020_b N_A_481_107#_c_1036_n 0.0292845f $X=-0.33 $Y=-0.265 $X2=2.89
+ $Y2=3.72
cc_66 N_VNB_M1020_b N_A_481_107#_c_1037_n 0.0184968f $X=-0.33 $Y=-0.265 $X2=2.77
+ $Y2=2.8
cc_67 N_VNB_M1020_b N_A_481_107#_c_1038_n 0.0567952f $X=-0.33 $Y=-0.265
+ $X2=4.925 $Y2=1.607
cc_68 N_VNB_c_3_p N_A_481_107#_c_1038_n 0.00235285f $X=0.24 $Y=0 $X2=4.925
+ $Y2=1.607
cc_69 N_VNB_M1020_b N_A_481_107#_c_1040_n 0.014726f $X=-0.33 $Y=-0.265 $X2=2.855
+ $Y2=1.607
cc_70 N_VNB_c_3_p N_A_481_107#_c_1040_n 5.63772e-19 $X=0.24 $Y=0 $X2=2.855
+ $Y2=1.607
cc_71 N_VNB_M1020_b N_A_481_107#_c_1042_n 0.00766022f $X=-0.33 $Y=-0.265
+ $X2=2.87 $Y2=1.53
cc_72 N_VNB_M1020_b N_A_481_107#_c_1043_n 0.00396487f $X=-0.33 $Y=-0.265
+ $X2=2.975 $Y2=2.97
cc_73 N_VNB_M1020_b N_A_481_107#_c_1044_n 0.0174954f $X=-0.33 $Y=-0.265
+ $X2=2.975 $Y2=3.635
cc_74 N_VNB_M1020_b N_A_481_107#_c_1045_n 0.00530439f $X=-0.33 $Y=-0.265
+ $X2=0.73 $Y2=2.415
cc_75 N_VNB_M1020_b N_A_481_107#_c_1046_n 0.00323482f $X=-0.33 $Y=-0.265
+ $X2=0.73 $Y2=2.45
cc_76 N_VNB_M1020_b N_A_1097_627#_c_1185_n 0.0168821f $X=-0.33 $Y=-0.265
+ $X2=2.03 $Y2=3.635
cc_77 N_VNB_M1020_b N_A_1097_627#_c_1186_n 0.00705523f $X=-0.33 $Y=-0.265
+ $X2=2.77 $Y2=2.8
cc_78 N_VNB_M1020_b N_A_1097_627#_c_1187_n 0.0276624f $X=-0.33 $Y=-0.265
+ $X2=2.87 $Y2=1.607
cc_79 N_VNB_M1020_b N_A_1097_627#_c_1188_n 0.00430589f $X=-0.33 $Y=-0.265
+ $X2=2.87 $Y2=1.53
cc_80 N_VNB_M1020_b N_A_1097_627#_c_1189_n 0.0198854f $X=-0.33 $Y=-0.265
+ $X2=2.975 $Y2=3.635
cc_81 N_VNB_M1020_b N_X_c_1296_n 0.0624574f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_82 N_VNB_c_3_p N_X_c_1296_n 4.98928e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_83 N_VNB_M1020_b N_VGND_c_1309_n 0.0495712f $X=-0.33 $Y=-0.265 $X2=2.935
+ $Y2=0.745
cc_84 N_VNB_c_3_p N_VGND_c_1309_n 0.00269373f $X=0.24 $Y=0 $X2=2.935 $Y2=0.745
cc_85 N_VNB_M1020_b N_VGND_c_1311_n 0.0491776f $X=-0.33 $Y=-0.265 $X2=4.925
+ $Y2=1.607
cc_86 N_VNB_c_3_p N_VGND_c_1311_n 0.00270129f $X=0.24 $Y=0 $X2=4.925 $Y2=1.607
cc_87 N_VNB_M1020_b N_VGND_c_1313_n 0.0438232f $X=-0.33 $Y=-0.265 $X2=2.87
+ $Y2=1.53
cc_88 N_VNB_c_3_p N_VGND_c_1313_n 0.00150031f $X=0.24 $Y=0 $X2=2.87 $Y2=1.53
cc_89 N_VNB_M1020_b N_VGND_c_1315_n 0.0561597f $X=-0.33 $Y=-0.265 $X2=2.07
+ $Y2=2.47
cc_90 N_VNB_c_3_p N_VGND_c_1315_n 0.00252021f $X=0.24 $Y=0 $X2=2.07 $Y2=2.47
cc_91 N_VNB_M1020_b N_VGND_c_1317_n 0.171325f $X=-0.33 $Y=-0.265 $X2=2.975
+ $Y2=2.885
cc_92 N_VNB_c_3_p N_VGND_c_1317_n 1.33335f $X=0.24 $Y=0 $X2=2.975 $Y2=2.885
cc_93 N_VPB_M1013_b N_S0_c_230_n 0.0480505f $X=-0.33 $Y=1.885 $X2=2.155 $Y2=2.83
cc_94 N_VPB_M1013_b N_S0_M1023_g 0.0494778f $X=-0.33 $Y=1.885 $X2=2.155
+ $Y2=3.345
cc_95 N_VPB_c_95_p N_S0_M1023_g 0.00232682f $X=12.24 $Y=4.07 $X2=2.155 $Y2=3.345
cc_96 N_VPB_M1013_b N_S0_c_217_n 0.13854f $X=-0.33 $Y=1.885 $X2=5.41 $Y2=1.945
cc_97 N_VPB_M1013_b N_S0_M1018_g 0.0555231f $X=-0.33 $Y=1.885 $X2=6.015
+ $Y2=3.345
cc_98 VPB N_S0_M1018_g 0.0023833f $X=0 $Y=3.955 $X2=6.015 $Y2=3.345
cc_99 N_VPB_c_95_p N_S0_M1018_g 0.0117159f $X=12.24 $Y=4.07 $X2=6.015 $Y2=3.345
cc_100 N_VPB_M1013_b N_S0_c_237_n 0.0249226f $X=-0.33 $Y=1.885 $X2=1.905
+ $Y2=2.415
cc_101 N_VPB_M1013_b N_S0_c_238_n 0.00206759f $X=-0.33 $Y=1.885 $X2=2.03 $Y2=2.5
cc_102 N_VPB_M1013_b N_S0_c_239_n 0.00563378f $X=-0.33 $Y=1.885 $X2=2.89
+ $Y2=3.72
cc_103 VPB N_S0_c_239_n 0.00305249f $X=0 $Y=3.955 $X2=2.89 $Y2=3.72
cc_104 N_VPB_c_95_p N_S0_c_239_n 0.0597733f $X=12.24 $Y=4.07 $X2=2.89 $Y2=3.72
cc_105 N_VPB_M1013_b N_S0_c_242_n 0.00260995f $X=-0.33 $Y=1.885 $X2=2.155
+ $Y2=3.72
cc_106 VPB N_S0_c_242_n 8.36161e-19 $X=0 $Y=3.955 $X2=2.155 $Y2=3.72
cc_107 N_VPB_c_95_p N_S0_c_242_n 0.0169098f $X=12.24 $Y=4.07 $X2=2.155 $Y2=3.72
cc_108 N_VPB_M1013_b N_S0_c_220_n 4.1969e-19 $X=-0.33 $Y=1.885 $X2=2.77 $Y2=2.8
cc_109 N_VPB_M1013_b N_S0_c_246_n 0.00109946f $X=-0.33 $Y=1.885 $X2=2.975
+ $Y2=2.885
cc_110 N_VPB_M1013_b N_S0_M1020_g 0.148971f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=0.745
cc_111 VPB N_S0_M1020_g 9.8192e-19 $X=0 $Y=3.955 $X2=0.665 $Y2=0.745
cc_112 N_VPB_c_95_p N_S0_M1020_g 0.00625941f $X=12.24 $Y=4.07 $X2=0.665
+ $Y2=0.745
cc_113 N_VPB_M1013_b N_A2_c_390_n 0.0781288f $X=-0.33 $Y=1.885 $X2=2.155
+ $Y2=3.345
cc_114 N_VPB_M1013_b N_A2_M1000_g 0.0361993f $X=-0.33 $Y=1.885 $X2=5.41
+ $Y2=1.945
cc_115 VPB N_A2_M1000_g 6.00592e-19 $X=0 $Y=3.955 $X2=5.41 $Y2=1.945
cc_116 N_VPB_c_95_p N_A2_M1000_g 0.00496941f $X=12.24 $Y=4.07 $X2=5.41 $Y2=1.945
cc_117 N_VPB_M1013_b N_A2_c_399_n 0.0250397f $X=-0.33 $Y=1.885 $X2=6.015
+ $Y2=3.345
cc_118 N_VPB_M1013_b A2 0.00360544f $X=-0.33 $Y=1.885 $X2=6.015 $Y2=3.345
cc_119 N_VPB_M1013_b N_A_30_107#_M1016_g 0.0706357f $X=-0.33 $Y=1.885 $X2=5.41
+ $Y2=1.945
cc_120 VPB N_A_30_107#_M1016_g 6.12208e-19 $X=0 $Y=3.955 $X2=5.41 $Y2=1.945
cc_121 N_VPB_c_95_p N_A_30_107#_M1016_g 0.00472818f $X=12.24 $Y=4.07 $X2=5.41
+ $Y2=1.945
cc_122 N_VPB_M1013_b N_A_30_107#_M1001_g 0.046674f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_123 VPB N_A_30_107#_M1001_g 0.00238149f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_124 N_VPB_c_95_p N_A_30_107#_M1001_g 0.0117022f $X=12.24 $Y=4.07 $X2=0 $Y2=0
cc_125 N_VPB_M1013_b N_A_30_107#_c_445_n 0.0291488f $X=-0.33 $Y=1.885 $X2=4.925
+ $Y2=1.607
cc_126 N_VPB_M1013_b N_A_30_107#_c_446_n 0.00395841f $X=-0.33 $Y=1.885 $X2=2.87
+ $Y2=1.53
cc_127 N_VPB_M1013_b N_A_30_107#_c_447_n 0.0569946f $X=-0.33 $Y=1.885 $X2=2.975
+ $Y2=2.97
cc_128 N_VPB_M1013_b N_A_30_107#_c_448_n 0.00717989f $X=-0.33 $Y=1.885 $X2=0.73
+ $Y2=2.415
cc_129 N_VPB_M1013_b N_A_30_107#_c_432_n 0.00105996f $X=-0.33 $Y=1.885 $X2=2.07
+ $Y2=2.47
cc_130 N_VPB_M1013_b N_A_30_107#_c_450_n 0.0221168f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_131 VPB N_A_30_107#_c_450_n 8.17695e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_132 N_VPB_c_95_p N_A_30_107#_c_450_n 0.0090966f $X=12.24 $Y=4.07 $X2=0 $Y2=0
cc_133 N_VPB_M1013_b N_A_30_107#_c_434_n 0.0595727f $X=-0.33 $Y=1.885 $X2=4.955
+ $Y2=0.84
cc_134 N_VPB_M1013_b N_A_30_107#_c_454_n 0.00114685f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_135 N_VPB_M1013_b N_A_30_107#_c_438_n 0.143905f $X=-0.33 $Y=1.885 $X2=5.41
+ $Y2=1.08
cc_136 N_VPB_M1013_b N_A3_M1009_g 0.0362137f $X=-0.33 $Y=1.885 $X2=5.375
+ $Y2=0.745
cc_137 N_VPB_c_95_p N_A3_M1009_g 0.00263287f $X=12.24 $Y=4.07 $X2=5.375
+ $Y2=0.745
cc_138 N_VPB_M1013_b A3 0.00517285f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_139 N_VPB_M1013_b N_A3_c_577_n 0.0682347f $X=-0.33 $Y=1.885 $X2=2.935
+ $Y2=1.085
cc_140 N_VPB_M1013_b N_A3_c_573_n 0.0308135f $X=-0.33 $Y=1.885 $X2=6.015
+ $Y2=2.37
cc_141 N_VPB_M1013_b N_A1_c_621_n 0.138977f $X=-0.33 $Y=1.885 $X2=2.935
+ $Y2=0.745
cc_142 VPB N_A1_c_621_n 0.0023833f $X=0 $Y=3.955 $X2=2.935 $Y2=0.745
cc_143 N_VPB_c_95_p N_A1_c_621_n 0.0119141f $X=12.24 $Y=4.07 $X2=2.935 $Y2=0.745
cc_144 N_VPB_M1013_b N_A0_M1019_g 0.0888666f $X=-0.33 $Y=1.885 $X2=2.155
+ $Y2=3.345
cc_145 N_VPB_c_95_p N_A0_M1019_g 0.00263287f $X=12.24 $Y=4.07 $X2=2.155
+ $Y2=3.345
cc_146 N_VPB_M1013_b N_A0_c_666_n 0.0651272f $X=-0.33 $Y=1.885 $X2=6.015
+ $Y2=3.345
cc_147 N_VPB_M1013_b A0 0.00185361f $X=-0.33 $Y=1.885 $X2=2.945 $Y2=1.085
cc_148 N_VPB_M1013_b N_A0_c_663_n 0.00958111f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_149 N_VPB_M1013_b N_S1_M1003_g 0.0417086f $X=-0.33 $Y=1.885 $X2=2.155
+ $Y2=3.345
cc_150 VPB N_S1_M1003_g 0.00211427f $X=0 $Y=3.955 $X2=2.155 $Y2=3.345
cc_151 N_VPB_c_95_p N_S1_M1003_g 0.0101113f $X=12.24 $Y=4.07 $X2=2.155 $Y2=3.345
cc_152 N_VPB_M1013_b N_S1_c_704_n 0.0177101f $X=-0.33 $Y=1.885 $X2=5.375
+ $Y2=1.08
cc_153 N_VPB_M1013_b N_S1_c_706_n 0.0305581f $X=-0.33 $Y=1.885 $X2=5.41
+ $Y2=1.945
cc_154 N_VPB_M1013_b N_S1_M1014_g 0.058647f $X=-0.33 $Y=1.885 $X2=2.935
+ $Y2=0.745
cc_155 N_VPB_M1013_b N_S1_c_708_n 0.00775937f $X=-0.33 $Y=1.885 $X2=2.935
+ $Y2=1.085
cc_156 N_VPB_M1013_b N_S1_c_716_n 0.0154091f $X=-0.33 $Y=1.885 $X2=5.41
+ $Y2=1.945
cc_157 N_VPB_M1013_b N_S1_c_717_n 3.33139e-19 $X=-0.33 $Y=1.885 $X2=6.015
+ $Y2=2.37
cc_158 N_VPB_M1013_b N_S1_c_718_n 0.00454801f $X=-0.33 $Y=1.885 $X2=2.89
+ $Y2=3.72
cc_159 N_VPB_M1013_b S1 0.0180885f $X=-0.33 $Y=1.885 $X2=2.77 $Y2=2.8
cc_160 N_VPB_M1013_b N_S1_c_720_n 0.0900019f $X=-0.33 $Y=1.885 $X2=2.975
+ $Y2=3.635
cc_161 N_VPB_M1013_b N_A_1681_89#_c_791_n 0.0277009f $X=-0.33 $Y=1.885 $X2=5.41
+ $Y2=1.365
cc_162 N_VPB_M1013_b N_A_1681_89#_M1017_g 0.0422907f $X=-0.33 $Y=1.885 $X2=6.015
+ $Y2=3.345
cc_163 N_VPB_c_95_p N_A_1681_89#_M1017_g 6.36627e-19 $X=12.24 $Y=4.07 $X2=6.015
+ $Y2=3.345
cc_164 N_VPB_M1013_b N_A_1681_89#_c_798_n 0.0638821f $X=-0.33 $Y=1.885 $X2=2.935
+ $Y2=1.085
cc_165 N_VPB_M1013_b N_A_1681_89#_c_794_n 0.00267845f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_166 N_VPB_M1013_b N_A_1681_89#_c_800_n 0.145059f $X=-0.33 $Y=1.885 $X2=2.03
+ $Y2=2.5
cc_167 N_VPB_M1013_b N_A_1681_89#_c_801_n 0.0204114f $X=-0.33 $Y=1.885 $X2=2.89
+ $Y2=3.72
cc_168 N_VPB_M1013_b N_A_1669_615#_c_867_n 2.31702e-19 $X=-0.33 $Y=1.885
+ $X2=5.41 $Y2=1.945
cc_169 N_VPB_M1013_b N_A_1669_615#_c_868_n 0.0422592f $X=-0.33 $Y=1.885
+ $X2=6.015 $Y2=3.345
cc_170 VPB N_A_1669_615#_c_868_n 0.00749497f $X=0 $Y=3.955 $X2=6.015 $Y2=3.345
cc_171 N_VPB_c_95_p N_A_1669_615#_c_868_n 0.146261f $X=12.24 $Y=4.07 $X2=6.015
+ $Y2=3.345
cc_172 N_VPB_M1013_b N_A_1669_615#_c_871_n 0.00338087f $X=-0.33 $Y=1.885
+ $X2=6.015 $Y2=3.345
cc_173 VPB N_A_1669_615#_c_871_n 0.00110413f $X=0 $Y=3.955 $X2=6.015 $Y2=3.345
cc_174 N_VPB_c_95_p N_A_1669_615#_c_871_n 0.0222578f $X=12.24 $Y=4.07 $X2=6.015
+ $Y2=3.345
cc_175 N_VPB_M1013_b N_A_1669_615#_c_874_n 0.0320372f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_176 N_VPB_M1013_b N_A_1669_615#_c_864_n 0.0054287f $X=-0.33 $Y=1.885 $X2=2.03
+ $Y2=2.5
cc_177 N_VPB_M1013_b N_A_1669_615#_M1022_g 0.0632232f $X=-0.33 $Y=1.885 $X2=2.77
+ $Y2=2.8
cc_178 VPB N_A_1669_615#_M1022_g 0.00970178f $X=0 $Y=3.955 $X2=2.77 $Y2=2.8
cc_179 N_VPB_c_95_p N_A_1669_615#_M1022_g 0.0152133f $X=12.24 $Y=4.07 $X2=2.77
+ $Y2=2.8
cc_180 N_VPB_M1013_b N_VPWR_c_931_n 0.00970639f $X=-0.33 $Y=1.885 $X2=2.935
+ $Y2=0.745
cc_181 VPB N_VPWR_c_931_n 0.0026951f $X=0 $Y=3.955 $X2=2.935 $Y2=0.745
cc_182 N_VPB_c_95_p N_VPWR_c_931_n 0.0409241f $X=12.24 $Y=4.07 $X2=2.935
+ $Y2=0.745
cc_183 N_VPB_M1013_b N_VPWR_c_934_n 0.0250993f $X=-0.33 $Y=1.885 $X2=2.855
+ $Y2=1.607
cc_184 VPB N_VPWR_c_934_n 0.00269683f $X=0 $Y=3.955 $X2=2.855 $Y2=1.607
cc_185 N_VPB_c_95_p N_VPWR_c_934_n 0.0408562f $X=12.24 $Y=4.07 $X2=2.855
+ $Y2=1.607
cc_186 N_VPB_M1013_b N_VPWR_c_937_n 0.0174766f $X=-0.33 $Y=1.885 $X2=2.03
+ $Y2=2.402
cc_187 VPB N_VPWR_c_937_n 0.00269683f $X=0 $Y=3.955 $X2=2.03 $Y2=2.402
cc_188 N_VPB_c_95_p N_VPWR_c_937_n 0.0408562f $X=12.24 $Y=4.07 $X2=2.03
+ $Y2=2.402
cc_189 N_VPB_M1013_b N_VPWR_c_940_n 0.0197524f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_940_n 0.00337025f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_191 N_VPB_c_95_p N_VPWR_c_940_n 0.0454439f $X=12.24 $Y=4.07 $X2=0 $Y2=0
cc_192 N_VPB_M1013_b N_VPWR_c_943_n 0.120999f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=0.745
cc_193 VPB N_VPWR_c_943_n 1.333f $X=0 $Y=3.955 $X2=0.665 $Y2=0.745
cc_194 N_VPB_c_95_p N_VPWR_c_943_n 0.0604828f $X=12.24 $Y=4.07 $X2=0.665
+ $Y2=0.745
cc_195 N_VPB_M1013_b N_A_481_107#_c_1029_n 0.0098471f $X=-0.33 $Y=1.885
+ $X2=2.935 $Y2=1.085
cc_196 N_VPB_M1013_b N_A_481_107#_c_1045_n 0.0105244f $X=-0.33 $Y=1.885 $X2=0.73
+ $Y2=2.415
cc_197 N_VPB_M1013_b N_A_481_107#_c_1049_n 0.012926f $X=-0.33 $Y=1.885 $X2=2.975
+ $Y2=2.885
cc_198 N_VPB_M1013_b N_A_1097_627#_c_1190_n 0.00326637f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_199 N_VPB_M1013_b N_A_1097_627#_c_1191_n 0.00188589f $X=-0.33 $Y=1.885
+ $X2=2.935 $Y2=0.745
cc_200 VPB N_A_1097_627#_c_1191_n 8.90907e-19 $X=0 $Y=3.955 $X2=2.935 $Y2=0.745
cc_201 N_VPB_c_95_p N_A_1097_627#_c_1191_n 0.0095893f $X=12.24 $Y=4.07 $X2=2.935
+ $Y2=0.745
cc_202 N_VPB_M1013_b N_A_1097_627#_c_1194_n 0.0071263f $X=-0.33 $Y=1.885
+ $X2=1.905 $Y2=2.415
cc_203 N_VPB_M1013_b N_A_1097_627#_c_1195_n 9.3168e-19 $X=-0.33 $Y=1.885
+ $X2=0.895 $Y2=2.415
cc_204 N_VPB_M1013_b N_A_1097_627#_c_1185_n 0.00808116f $X=-0.33 $Y=1.885
+ $X2=2.03 $Y2=3.635
cc_205 N_VPB_M1013_b N_A_1097_627#_c_1197_n 0.0195903f $X=-0.33 $Y=1.885
+ $X2=2.89 $Y2=3.72
cc_206 N_VPB_M1013_b N_A_1097_627#_c_1186_n 0.0208156f $X=-0.33 $Y=1.885
+ $X2=2.77 $Y2=2.8
cc_207 N_VPB_M1013_b N_A_1097_627#_c_1199_n 0.00517222f $X=-0.33 $Y=1.885
+ $X2=2.855 $Y2=1.607
cc_208 N_VPB_M1013_b N_A_1097_627#_c_1200_n 0.00177216f $X=-0.33 $Y=1.885
+ $X2=0.73 $Y2=2.45
cc_209 N_VPB_M1013_b N_A_1097_627#_c_1201_n 4.83942e-19 $X=-0.33 $Y=1.885
+ $X2=0.73 $Y2=2.45
cc_210 N_VPB_M1013_b N_A_1097_627#_c_1202_n 0.00213799f $X=-0.33 $Y=1.885
+ $X2=2.03 $Y2=2.402
cc_211 N_VPB_M1013_b N_A_1097_627#_c_1203_n 0.00755711f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_212 VPB N_A_1097_627#_c_1203_n 9.62901e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_213 N_VPB_c_95_p N_A_1097_627#_c_1203_n 0.0100117f $X=12.24 $Y=4.07 $X2=0
+ $Y2=0
cc_214 N_VPB_M1013_b N_X_c_1296_n 0.0694102f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_215 VPB N_X_c_1296_n 7.36921e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_216 N_VPB_c_95_p N_X_c_1296_n 0.0120479f $X=12.24 $Y=4.07 $X2=0 $Y2=0
cc_217 N_S0_c_230_n N_A2_c_390_n 0.0478513f $X=2.155 $Y=2.83 $X2=0 $Y2=0
cc_218 N_S0_c_237_n N_A2_c_390_n 0.0411045f $X=1.905 $Y=2.415 $X2=0 $Y2=0
cc_219 N_S0_c_252_p N_A2_c_390_n 0.00665575f $X=2.03 $Y=3.635 $X2=0 $Y2=0
cc_220 N_S0_c_253_p N_A2_c_390_n 0.00288456f $X=0.73 $Y=2.45 $X2=0 $Y2=0
cc_221 N_S0_M1020_g N_A2_M1006_g 0.0360626f $X=0.665 $Y=0.745 $X2=-0.33
+ $Y2=-0.265
cc_222 N_S0_c_242_n N_A2_M1000_g 2.16406e-19 $X=2.155 $Y=3.72 $X2=0 $Y2=0
cc_223 N_S0_M1020_g N_A2_M1000_g 0.0145705f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_224 N_S0_M1023_g N_A2_c_399_n 0.0478513f $X=2.155 $Y=3.345 $X2=0.24 $Y2=0
cc_225 N_S0_c_237_n A2 0.0315708f $X=1.905 $Y=2.415 $X2=0 $Y2=0
cc_226 N_S0_M1020_g A2 0.0158951f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_227 N_S0_M1020_g N_A2_c_394_n 0.0876383f $X=0.665 $Y=0.745 $X2=12.24 $Y2=0
cc_228 N_S0_M1023_g N_A_30_107#_M1016_g 0.0168533f $X=2.155 $Y=3.345 $X2=0 $Y2=0
cc_229 N_S0_c_252_p N_A_30_107#_M1016_g 0.00103479f $X=2.03 $Y=3.635 $X2=0 $Y2=0
cc_230 N_S0_c_239_n N_A_30_107#_M1016_g 0.0126159f $X=2.89 $Y=3.72 $X2=0 $Y2=0
cc_231 N_S0_c_220_n N_A_30_107#_M1016_g 0.00719605f $X=2.77 $Y=2.8 $X2=0 $Y2=0
cc_232 N_S0_c_265_p N_A_30_107#_M1016_g 0.0274205f $X=2.975 $Y=3.635 $X2=0 $Y2=0
cc_233 N_S0_c_246_n N_A_30_107#_M1016_g 0.0230901f $X=2.975 $Y=2.885 $X2=0 $Y2=0
cc_234 N_S0_M1018_g N_A_30_107#_M1001_g 0.0136979f $X=6.015 $Y=3.345 $X2=0 $Y2=0
cc_235 N_S0_M1020_g N_A_30_107#_c_429_n 0.0213595f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_236 N_S0_M1020_g N_A_30_107#_c_431_n 0.0387426f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_237 N_S0_c_230_n N_A_30_107#_c_465_n 2.80812e-19 $X=2.155 $Y=2.83 $X2=0 $Y2=0
cc_238 N_S0_c_238_n N_A_30_107#_c_465_n 0.0144543f $X=2.03 $Y=2.5 $X2=0 $Y2=0
cc_239 N_S0_c_221_n N_A_30_107#_c_445_n 0.116733f $X=4.925 $Y=1.607 $X2=0 $Y2=0
cc_240 N_S0_c_229_n N_A_30_107#_c_445_n 0.0064521f $X=5.172 $Y=1.445 $X2=0 $Y2=0
cc_241 N_S0_c_217_n N_A_30_107#_c_446_n 0.0114377f $X=5.41 $Y=1.945 $X2=0 $Y2=0
cc_242 N_S0_c_217_n N_A_30_107#_c_447_n 0.0486172f $X=5.41 $Y=1.945 $X2=0 $Y2=0
cc_243 N_S0_M1018_g N_A_30_107#_c_447_n 0.00505697f $X=6.015 $Y=3.345 $X2=0
+ $Y2=0
cc_244 N_S0_c_229_n N_A_30_107#_c_447_n 5.91057e-19 $X=5.172 $Y=1.445 $X2=0
+ $Y2=0
cc_245 N_S0_c_217_n N_A_30_107#_c_448_n 0.0603921f $X=5.41 $Y=1.945 $X2=0 $Y2=0
cc_246 N_S0_c_229_n N_A_30_107#_c_448_n 0.00611037f $X=5.172 $Y=1.445 $X2=0
+ $Y2=0
cc_247 N_S0_c_217_n N_A_30_107#_c_432_n 0.0112723f $X=5.41 $Y=1.945 $X2=0 $Y2=0
cc_248 S0 N_A_30_107#_c_432_n 0.0114062f $X=4.955 $Y=0.84 $X2=0 $Y2=0
cc_249 N_S0_c_227_n N_A_30_107#_c_432_n 0.00287809f $X=5.31 $Y=1.265 $X2=0 $Y2=0
cc_250 N_S0_c_229_n N_A_30_107#_c_432_n 0.0110597f $X=5.172 $Y=1.445 $X2=0 $Y2=0
cc_251 N_S0_M1020_g N_A_30_107#_c_433_n 0.00513266f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_252 N_S0_M1020_g N_A_30_107#_c_450_n 0.00963741f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_253 N_S0_c_253_p N_A_30_107#_c_434_n 0.0303771f $X=0.73 $Y=2.45 $X2=0 $Y2=0
cc_254 N_S0_M1020_g N_A_30_107#_c_434_n 0.0603071f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_255 N_S0_c_220_n N_A_30_107#_c_483_n 0.045692f $X=2.77 $Y=2.8 $X2=0 $Y2=0
cc_256 N_S0_c_221_n N_A_30_107#_c_483_n 0.0200419f $X=4.925 $Y=1.607 $X2=0 $Y2=0
cc_257 N_S0_c_246_n N_A_30_107#_c_483_n 0.00174365f $X=2.975 $Y=2.885 $X2=0
+ $Y2=0
cc_258 N_S0_c_217_n N_A_30_107#_c_454_n 0.00999137f $X=5.41 $Y=1.945 $X2=0 $Y2=0
cc_259 N_S0_c_229_n N_A_30_107#_c_454_n 0.0277651f $X=5.172 $Y=1.445 $X2=0 $Y2=0
cc_260 N_S0_M1025_g N_A_30_107#_M1007_g 0.0138153f $X=2.935 $Y=0.745 $X2=0 $Y2=0
cc_261 N_S0_c_222_n N_A_30_107#_M1007_g 3.59453e-19 $X=2.855 $Y=1.607 $X2=0
+ $Y2=0
cc_262 N_S0_c_223_n N_A_30_107#_M1007_g 0.0193996f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_263 N_S0_c_217_n N_A_30_107#_M1021_g 0.0240924f $X=5.41 $Y=1.945 $X2=0 $Y2=0
cc_264 S0 N_A_30_107#_M1021_g 0.00162465f $X=4.955 $Y=0.84 $X2=0 $Y2=0
cc_265 N_S0_c_227_n N_A_30_107#_M1021_g 0.0451649f $X=5.31 $Y=1.265 $X2=0 $Y2=0
cc_266 N_S0_c_228_n N_A_30_107#_M1021_g 0.0153448f $X=5.41 $Y=1.08 $X2=0 $Y2=0
cc_267 N_S0_c_229_n N_A_30_107#_M1021_g 7.21105e-19 $X=5.172 $Y=1.445 $X2=0
+ $Y2=0
cc_268 N_S0_c_230_n N_A_30_107#_c_438_n 0.0540518f $X=2.155 $Y=2.83 $X2=0 $Y2=0
cc_269 N_S0_c_238_n N_A_30_107#_c_438_n 0.00111137f $X=2.03 $Y=2.5 $X2=0 $Y2=0
cc_270 N_S0_c_220_n N_A_30_107#_c_438_n 0.0326032f $X=2.77 $Y=2.8 $X2=0 $Y2=0
cc_271 N_S0_c_221_n N_A_30_107#_c_438_n 0.00827055f $X=4.925 $Y=1.607 $X2=0
+ $Y2=0
cc_272 N_S0_c_222_n N_A_30_107#_c_438_n 0.00109631f $X=2.855 $Y=1.607 $X2=0
+ $Y2=0
cc_273 N_S0_c_223_n N_A_30_107#_c_438_n 0.0408008f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_274 N_S0_M1025_g N_A3_M1002_g 0.0410449f $X=2.935 $Y=0.745 $X2=0 $Y2=0
cc_275 N_S0_c_265_p N_A3_M1009_g 4.83397e-19 $X=2.975 $Y=3.635 $X2=0 $Y2=0
cc_276 N_S0_c_221_n N_A3_c_572_n 0.0223967f $X=4.925 $Y=1.607 $X2=0 $Y2=0
cc_277 N_S0_c_223_n N_A3_c_572_n 0.0410449f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_278 N_S0_c_220_n A3 0.00506602f $X=2.77 $Y=2.8 $X2=0 $Y2=0
cc_279 N_S0_c_246_n A3 0.00463837f $X=2.975 $Y=2.885 $X2=0 $Y2=0
cc_280 N_S0_c_265_p N_A3_c_577_n 6.9993e-19 $X=2.975 $Y=3.635 $X2=0 $Y2=0
cc_281 N_S0_c_246_n N_A3_c_577_n 4.19745e-19 $X=2.975 $Y=2.885 $X2=0 $Y2=0
cc_282 N_S0_c_220_n N_A3_c_573_n 0.00341716f $X=2.77 $Y=2.8 $X2=0 $Y2=0
cc_283 N_S0_c_221_n N_A3_c_573_n 0.0211927f $X=4.925 $Y=1.607 $X2=0 $Y2=0
cc_284 N_S0_c_223_n N_A3_c_573_n 0.00386878f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_285 S0 N_A1_M1004_g 0.0102271f $X=4.955 $Y=0.84 $X2=0 $Y2=0
cc_286 N_S0_c_228_n N_A1_M1004_g 0.0396082f $X=5.41 $Y=1.08 $X2=0 $Y2=0
cc_287 N_S0_c_221_n N_A1_c_620_n 0.0350336f $X=4.925 $Y=1.607 $X2=0 $Y2=0
cc_288 N_S0_c_227_n N_A1_c_620_n 0.0396082f $X=5.31 $Y=1.265 $X2=0 $Y2=0
cc_289 N_S0_c_217_n N_A1_c_621_n 0.0202531f $X=5.41 $Y=1.945 $X2=0 $Y2=0
cc_290 N_S0_c_221_n N_A1_c_621_n 0.0204342f $X=4.925 $Y=1.607 $X2=0 $Y2=0
cc_291 N_S0_M1018_g N_A0_M1019_g 0.0573752f $X=6.015 $Y=3.345 $X2=0 $Y2=0
cc_292 N_S0_c_217_n N_A0_c_666_n 0.0573752f $X=5.41 $Y=1.945 $X2=0.24 $Y2=0
cc_293 N_S0_c_217_n N_A0_c_663_n 9.34053e-19 $X=5.41 $Y=1.945 $X2=6.24 $Y2=0
cc_294 N_S0_M1023_g N_VPWR_c_931_n 0.00177353f $X=2.155 $Y=3.345 $X2=12.24 $Y2=0
cc_295 N_S0_c_237_n N_VPWR_c_931_n 0.0201785f $X=1.905 $Y=2.415 $X2=12.24 $Y2=0
cc_296 N_S0_c_252_p N_VPWR_c_931_n 0.0213993f $X=2.03 $Y=3.635 $X2=12.24 $Y2=0
cc_297 N_S0_c_242_n N_VPWR_c_931_n 0.0022356f $X=2.155 $Y=3.72 $X2=12.24 $Y2=0
cc_298 N_S0_c_253_p N_VPWR_c_931_n 0.0208557f $X=0.73 $Y=2.45 $X2=12.24 $Y2=0
cc_299 N_S0_M1020_g N_VPWR_c_931_n 0.0366407f $X=0.665 $Y=0.745 $X2=12.24 $Y2=0
cc_300 N_S0_c_239_n N_VPWR_c_934_n 0.00396986f $X=2.89 $Y=3.72 $X2=0 $Y2=0
cc_301 N_S0_c_265_p N_VPWR_c_934_n 0.033899f $X=2.975 $Y=3.635 $X2=0 $Y2=0
cc_302 N_S0_M1018_g N_VPWR_c_937_n 0.00868788f $X=6.015 $Y=3.345 $X2=0 $Y2=0
cc_303 N_S0_M1023_g N_VPWR_c_943_n 0.0101339f $X=2.155 $Y=3.345 $X2=0 $Y2=0
cc_304 N_S0_M1018_g N_VPWR_c_943_n 0.0177046f $X=6.015 $Y=3.345 $X2=0 $Y2=0
cc_305 N_S0_c_252_p N_VPWR_c_943_n 0.0275599f $X=2.03 $Y=3.635 $X2=0 $Y2=0
cc_306 N_S0_c_239_n N_VPWR_c_943_n 0.0329953f $X=2.89 $Y=3.72 $X2=0 $Y2=0
cc_307 N_S0_c_242_n N_VPWR_c_943_n 0.00985244f $X=2.155 $Y=3.72 $X2=0 $Y2=0
cc_308 N_S0_c_265_p N_VPWR_c_943_n 0.0137273f $X=2.975 $Y=3.635 $X2=0 $Y2=0
cc_309 N_S0_c_253_p N_VPWR_c_943_n 0.0027992f $X=0.73 $Y=2.45 $X2=0 $Y2=0
cc_310 N_S0_c_246_n N_VPWR_c_943_n 0.0042576f $X=2.975 $Y=2.885 $X2=0 $Y2=0
cc_311 N_S0_M1020_g N_VPWR_c_943_n 0.010171f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_312 N_S0_M1025_g N_A_481_107#_c_1027_n 0.0166948f $X=2.935 $Y=0.745 $X2=0
+ $Y2=0
cc_313 N_S0_c_223_n N_A_481_107#_c_1027_n 2.79871e-19 $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_314 N_S0_c_230_n N_A_481_107#_c_1029_n 0.0101907f $X=2.155 $Y=2.83 $X2=0
+ $Y2=0
cc_315 N_S0_M1023_g N_A_481_107#_c_1029_n 0.00898738f $X=2.155 $Y=3.345 $X2=0
+ $Y2=0
cc_316 N_S0_c_238_n N_A_481_107#_c_1029_n 0.0147768f $X=2.03 $Y=2.5 $X2=0 $Y2=0
cc_317 N_S0_c_252_p N_A_481_107#_c_1029_n 0.0452365f $X=2.03 $Y=3.635 $X2=0
+ $Y2=0
cc_318 N_S0_c_220_n N_A_481_107#_c_1029_n 0.0692626f $X=2.77 $Y=2.8 $X2=0 $Y2=0
cc_319 N_S0_c_222_n N_A_481_107#_c_1029_n 0.0263504f $X=2.855 $Y=1.607 $X2=0
+ $Y2=0
cc_320 N_S0_c_223_n N_A_481_107#_c_1029_n 0.00452311f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_321 N_S0_c_265_p N_A_481_107#_c_1029_n 0.00791373f $X=2.975 $Y=3.635 $X2=0
+ $Y2=0
cc_322 N_S0_c_246_n N_A_481_107#_c_1029_n 0.0122694f $X=2.975 $Y=2.885 $X2=0
+ $Y2=0
cc_323 N_S0_c_221_n N_A_481_107#_c_1030_n 0.120343f $X=4.925 $Y=1.607 $X2=0
+ $Y2=0
cc_324 N_S0_c_222_n N_A_481_107#_c_1030_n 0.0105152f $X=2.855 $Y=1.607 $X2=0
+ $Y2=0
cc_325 N_S0_c_223_n N_A_481_107#_c_1030_n 0.025682f $X=2.87 $Y=1.53 $X2=0 $Y2=0
cc_326 S0 N_A_481_107#_c_1030_n 0.00812389f $X=4.955 $Y=0.84 $X2=0 $Y2=0
cc_327 S0 N_A_481_107#_c_1031_n 0.00862159f $X=4.955 $Y=0.84 $X2=0 $Y2=0
cc_328 N_S0_c_228_n N_A_481_107#_c_1031_n 0.00183915f $X=5.41 $Y=1.08 $X2=0
+ $Y2=0
cc_329 S0 N_A_481_107#_c_1032_n 0.0116646f $X=4.955 $Y=0.84 $X2=6.24 $Y2=0.057
cc_330 N_S0_c_228_n N_A_481_107#_c_1032_n 0.0194616f $X=5.41 $Y=1.08 $X2=6.24
+ $Y2=0.057
cc_331 N_S0_c_222_n N_A_481_107#_c_1046_n 0.00216263f $X=2.855 $Y=1.607 $X2=0
+ $Y2=0
cc_332 N_S0_c_223_n N_A_481_107#_c_1046_n 0.00221915f $X=2.87 $Y=1.53 $X2=0
+ $Y2=0
cc_333 N_S0_M1023_g N_A_481_107#_c_1071_n 0.0064386f $X=2.155 $Y=3.345 $X2=0
+ $Y2=0
cc_334 N_S0_c_252_p N_A_481_107#_c_1071_n 0.019719f $X=2.03 $Y=3.635 $X2=0 $Y2=0
cc_335 N_S0_c_239_n N_A_481_107#_c_1071_n 0.0225376f $X=2.89 $Y=3.72 $X2=0 $Y2=0
cc_336 N_S0_c_265_p N_A_481_107#_c_1071_n 0.0191841f $X=2.975 $Y=3.635 $X2=0
+ $Y2=0
cc_337 N_S0_c_246_n N_A_481_107#_c_1071_n 0.00137264f $X=2.975 $Y=2.885 $X2=0
+ $Y2=0
cc_338 N_S0_c_217_n N_A_1097_627#_c_1190_n 0.00303219f $X=5.41 $Y=1.945 $X2=0
+ $Y2=0
cc_339 N_S0_M1018_g N_A_1097_627#_c_1190_n 0.0046141f $X=6.015 $Y=3.345 $X2=0
+ $Y2=0
cc_340 N_S0_M1018_g N_A_1097_627#_c_1191_n 0.00825441f $X=6.015 $Y=3.345 $X2=0
+ $Y2=0
cc_341 S0 N_A_1097_627#_c_1209_n 0.00816719f $X=4.955 $Y=0.84 $X2=12.24 $Y2=0
cc_342 N_S0_c_227_n N_A_1097_627#_c_1209_n 0.00195912f $X=5.31 $Y=1.265
+ $X2=12.24 $Y2=0
cc_343 N_S0_c_228_n N_A_1097_627#_c_1209_n 0.00814982f $X=5.41 $Y=1.08 $X2=12.24
+ $Y2=0
cc_344 N_S0_c_217_n N_A_1097_627#_c_1194_n 0.0161954f $X=5.41 $Y=1.945 $X2=6.24
+ $Y2=0.057
cc_345 N_S0_M1018_g N_A_1097_627#_c_1194_n 0.0171196f $X=6.015 $Y=3.345 $X2=6.24
+ $Y2=0.057
cc_346 N_S0_c_217_n N_A_1097_627#_c_1195_n 0.00994378f $X=5.41 $Y=1.945 $X2=6.24
+ $Y2=0.058
cc_347 N_S0_M1018_g N_A_1097_627#_c_1195_n 0.00150732f $X=6.015 $Y=3.345
+ $X2=6.24 $Y2=0.058
cc_348 N_S0_c_217_n N_A_1097_627#_c_1185_n 0.0145101f $X=5.41 $Y=1.945 $X2=0
+ $Y2=0
cc_349 N_S0_M1018_g N_A_1097_627#_c_1200_n 0.00561412f $X=6.015 $Y=3.345 $X2=0
+ $Y2=0
cc_350 N_S0_M1020_g N_VGND_c_1309_n 0.0360692f $X=0.665 $Y=0.745 $X2=12.24 $Y2=0
cc_351 N_S0_M1025_g N_VGND_c_1311_n 0.00760888f $X=2.935 $Y=0.745 $X2=0 $Y2=0
cc_352 N_S0_M1025_g N_VGND_c_1317_n 0.0169955f $X=2.935 $Y=0.745 $X2=0 $Y2=0
cc_353 S0 N_VGND_c_1317_n 0.0153664f $X=4.955 $Y=0.84 $X2=0 $Y2=0
cc_354 N_S0_M1020_g N_VGND_c_1317_n 0.00647854f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_355 N_S0_c_228_n N_VGND_c_1317_n 0.014404f $X=5.41 $Y=1.08 $X2=0 $Y2=0
cc_356 S0 A_983_107# 0.00136176f $X=4.955 $Y=0.84 $X2=0 $Y2=0
cc_357 N_A2_M1006_g N_A_30_107#_c_431_n 0.0320819f $X=1.445 $Y=0.745 $X2=0 $Y2=0
cc_358 A2 N_A_30_107#_c_431_n 0.0316839f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_359 N_A2_c_394_n N_A_30_107#_c_431_n 8.27069e-19 $X=1.35 $Y=1.665 $X2=0 $Y2=0
cc_360 N_A2_M1006_g N_A_30_107#_c_465_n 0.00351414f $X=1.445 $Y=0.745 $X2=0
+ $Y2=0
cc_361 A2 N_A_30_107#_c_465_n 0.019571f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_362 N_A2_M1006_g N_A_30_107#_M1007_g 0.0595969f $X=1.445 $Y=0.745 $X2=0 $Y2=0
cc_363 A2 N_A_30_107#_M1007_g 0.00182455f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_364 N_A2_c_394_n N_A_30_107#_c_438_n 0.0595969f $X=1.35 $Y=1.665 $X2=0 $Y2=0
cc_365 N_A2_M1000_g N_VPWR_c_931_n 0.0450226f $X=1.445 $Y=3.345 $X2=12.24 $Y2=0
cc_366 N_A2_c_399_n N_VPWR_c_931_n 0.00109591f $X=1.43 $Y=3.005 $X2=12.24 $Y2=0
cc_367 N_A2_M1000_g N_VPWR_c_943_n 0.00843377f $X=1.445 $Y=3.345 $X2=0 $Y2=0
cc_368 N_A2_M1006_g N_A_481_107#_c_1027_n 0.00217364f $X=1.445 $Y=0.745 $X2=0
+ $Y2=0
cc_369 N_A2_c_390_n N_A_481_107#_c_1029_n 0.00515278f $X=1.43 $Y=2.74 $X2=0
+ $Y2=0
cc_370 N_A2_M1006_g N_A_481_107#_c_1029_n 3.48044e-19 $X=1.445 $Y=0.745 $X2=0
+ $Y2=0
cc_371 N_A2_M1006_g N_A_481_107#_c_1046_n 2.92858e-19 $X=1.445 $Y=0.745 $X2=0
+ $Y2=0
cc_372 N_A2_M1006_g N_VGND_c_1309_n 0.0445503f $X=1.445 $Y=0.745 $X2=12.24 $Y2=0
cc_373 N_A2_M1006_g N_VGND_c_1317_n 0.00461913f $X=1.445 $Y=0.745 $X2=0 $Y2=0
cc_374 N_A_30_107#_c_445_n N_A3_c_572_n 5.26927e-19 $X=5.005 $Y=2.035 $X2=0
+ $Y2=0
cc_375 N_A_30_107#_M1016_g A3 0.00259855f $X=2.935 $Y=3.345 $X2=0 $Y2=0
cc_376 N_A_30_107#_c_445_n A3 0.0260111f $X=5.005 $Y=2.035 $X2=0 $Y2=0
cc_377 N_A_30_107#_c_483_n A3 0.0221412f $X=3.12 $Y=2.115 $X2=0 $Y2=0
cc_378 N_A_30_107#_c_438_n A3 0.00220706f $X=2.935 $Y=2.097 $X2=0 $Y2=0
cc_379 N_A_30_107#_M1016_g N_A3_c_577_n 0.0436364f $X=2.935 $Y=3.345 $X2=0 $Y2=0
cc_380 N_A_30_107#_c_445_n N_A3_c_577_n 3.92599e-19 $X=5.005 $Y=2.035 $X2=0
+ $Y2=0
cc_381 N_A_30_107#_c_483_n N_A3_c_577_n 7.69712e-19 $X=3.12 $Y=2.115 $X2=0 $Y2=0
cc_382 N_A_30_107#_c_438_n N_A3_c_577_n 0.0261778f $X=2.935 $Y=2.097 $X2=0 $Y2=0
cc_383 N_A_30_107#_c_445_n N_A3_c_573_n 0.0309993f $X=5.005 $Y=2.035 $X2=0 $Y2=0
cc_384 N_A_30_107#_c_483_n N_A3_c_573_n 9.42932e-19 $X=3.12 $Y=2.115 $X2=0 $Y2=0
cc_385 N_A_30_107#_c_438_n N_A3_c_573_n 0.0208989f $X=2.935 $Y=2.097 $X2=0 $Y2=0
cc_386 N_A_30_107#_c_445_n N_A1_c_620_n 6.27545e-19 $X=5.005 $Y=2.035 $X2=0
+ $Y2=0
cc_387 N_A_30_107#_c_445_n A1 0.0238596f $X=5.005 $Y=2.035 $X2=0 $Y2=0
cc_388 N_A_30_107#_c_446_n A1 0.0314456f $X=5.17 $Y=2.47 $X2=0 $Y2=0
cc_389 N_A_30_107#_c_447_n A1 0.00431043f $X=5.17 $Y=2.47 $X2=0 $Y2=0
cc_390 N_A_30_107#_c_445_n N_A1_c_621_n 0.0316262f $X=5.005 $Y=2.035 $X2=0 $Y2=0
cc_391 N_A_30_107#_c_446_n N_A1_c_621_n 0.00956096f $X=5.17 $Y=2.47 $X2=0 $Y2=0
cc_392 N_A_30_107#_c_447_n N_A1_c_621_n 0.0949415f $X=5.17 $Y=2.47 $X2=0 $Y2=0
cc_393 N_A_30_107#_M1021_g N_A0_M1008_g 0.0851655f $X=6.155 $Y=0.745 $X2=0 $Y2=0
cc_394 N_A_30_107#_c_450_n N_VPWR_c_931_n 0.0330272f $X=0.275 $Y=3.345 $X2=12.24
+ $Y2=0
cc_395 N_A_30_107#_M1016_g N_VPWR_c_934_n 0.00529904f $X=2.935 $Y=3.345 $X2=0
+ $Y2=0
cc_396 N_A_30_107#_c_483_n N_VPWR_c_934_n 5.6898e-19 $X=3.12 $Y=2.115 $X2=0
+ $Y2=0
cc_397 N_A_30_107#_c_438_n N_VPWR_c_934_n 3.46935e-19 $X=2.935 $Y=2.097 $X2=0
+ $Y2=0
cc_398 N_A_30_107#_M1016_g N_VPWR_c_943_n 0.012085f $X=2.935 $Y=3.345 $X2=0
+ $Y2=0
cc_399 N_A_30_107#_M1001_g N_VPWR_c_943_n 0.0218609f $X=5.235 $Y=3.345 $X2=0
+ $Y2=0
cc_400 N_A_30_107#_c_446_n N_VPWR_c_943_n 0.0108221f $X=5.17 $Y=2.47 $X2=0 $Y2=0
cc_401 N_A_30_107#_c_450_n N_VPWR_c_943_n 0.0320429f $X=0.275 $Y=3.345 $X2=0
+ $Y2=0
cc_402 N_A_30_107#_M1007_g N_A_481_107#_c_1027_n 0.0198949f $X=2.155 $Y=0.745
+ $X2=0 $Y2=0
cc_403 N_A_30_107#_M1016_g N_A_481_107#_c_1029_n 0.00218005f $X=2.935 $Y=3.345
+ $X2=0 $Y2=0
cc_404 N_A_30_107#_c_431_n N_A_481_107#_c_1029_n 0.00578689f $X=1.905 $Y=1.26
+ $X2=0 $Y2=0
cc_405 N_A_30_107#_c_465_n N_A_481_107#_c_1029_n 0.0459359f $X=2.07 $Y=1.53
+ $X2=0 $Y2=0
cc_406 N_A_30_107#_M1007_g N_A_481_107#_c_1029_n 0.00767827f $X=2.155 $Y=0.745
+ $X2=0 $Y2=0
cc_407 N_A_30_107#_c_438_n N_A_481_107#_c_1029_n 0.0405144f $X=2.935 $Y=2.097
+ $X2=0 $Y2=0
cc_408 N_A_30_107#_M1021_g N_A_481_107#_c_1032_n 0.0145483f $X=6.155 $Y=0.745
+ $X2=6.24 $Y2=0.057
cc_409 N_A_30_107#_M1021_g N_A_481_107#_c_1087_n 0.00170055f $X=6.155 $Y=0.745
+ $X2=0 $Y2=0
cc_410 N_A_30_107#_c_431_n N_A_481_107#_c_1046_n 0.00727324f $X=1.905 $Y=1.26
+ $X2=0 $Y2=0
cc_411 N_A_30_107#_M1007_g N_A_481_107#_c_1046_n 0.00638567f $X=2.155 $Y=0.745
+ $X2=0 $Y2=0
cc_412 N_A_30_107#_c_438_n N_A_481_107#_c_1046_n 0.00518079f $X=2.935 $Y=2.097
+ $X2=0 $Y2=0
cc_413 N_A_30_107#_M1016_g N_A_481_107#_c_1071_n 0.005177f $X=2.935 $Y=3.345
+ $X2=0 $Y2=0
cc_414 N_A_30_107#_M1001_g N_A_1097_627#_c_1190_n 0.00568589f $X=5.235 $Y=3.345
+ $X2=0 $Y2=0
cc_415 N_A_30_107#_M1001_g N_A_1097_627#_c_1191_n 0.00904624f $X=5.235 $Y=3.345
+ $X2=0 $Y2=0
cc_416 N_A_30_107#_c_432_n N_A_1097_627#_c_1209_n 0.0236476f $X=6.075 $Y=1.23
+ $X2=12.24 $Y2=0
cc_417 N_A_30_107#_M1021_g N_A_1097_627#_c_1209_n 0.0327251f $X=6.155 $Y=0.745
+ $X2=12.24 $Y2=0
cc_418 N_A_30_107#_c_448_n N_A_1097_627#_c_1194_n 0.0112102f $X=5.91 $Y=2.035
+ $X2=6.24 $Y2=0.057
cc_419 N_A_30_107#_c_446_n N_A_1097_627#_c_1195_n 0.00952474f $X=5.17 $Y=2.47
+ $X2=6.24 $Y2=0.058
cc_420 N_A_30_107#_c_447_n N_A_1097_627#_c_1195_n 0.00119855f $X=5.17 $Y=2.47
+ $X2=6.24 $Y2=0.058
cc_421 N_A_30_107#_c_448_n N_A_1097_627#_c_1195_n 0.00437975f $X=5.91 $Y=2.035
+ $X2=6.24 $Y2=0.058
cc_422 N_A_30_107#_c_448_n N_A_1097_627#_c_1185_n 0.0130071f $X=5.91 $Y=2.035
+ $X2=0 $Y2=0
cc_423 N_A_30_107#_c_432_n N_A_1097_627#_c_1185_n 0.0623798f $X=6.075 $Y=1.23
+ $X2=0 $Y2=0
cc_424 N_A_30_107#_M1021_g N_A_1097_627#_c_1185_n 0.00871791f $X=6.155 $Y=0.745
+ $X2=0 $Y2=0
cc_425 N_A_30_107#_M1001_g N_A_1097_627#_c_1200_n 0.00202671f $X=5.235 $Y=3.345
+ $X2=0 $Y2=0
cc_426 N_A_30_107#_c_447_n N_A_1097_627#_c_1200_n 0.0017875f $X=5.17 $Y=2.47
+ $X2=0 $Y2=0
cc_427 N_A_30_107#_c_429_n N_VGND_c_1309_n 0.0348344f $X=0.275 $Y=0.745
+ $X2=12.24 $Y2=0
cc_428 N_A_30_107#_c_431_n N_VGND_c_1309_n 0.0686854f $X=1.905 $Y=1.26 $X2=12.24
+ $Y2=0
cc_429 N_A_30_107#_M1007_g N_VGND_c_1309_n 0.00407355f $X=2.155 $Y=0.745
+ $X2=12.24 $Y2=0
cc_430 N_A_30_107#_c_429_n N_VGND_c_1317_n 0.0319953f $X=0.275 $Y=0.745 $X2=0
+ $Y2=0
cc_431 N_A_30_107#_c_431_n N_VGND_c_1317_n 0.0270407f $X=1.905 $Y=1.26 $X2=0
+ $Y2=0
cc_432 N_A_30_107#_c_432_n N_VGND_c_1317_n 0.0013739f $X=6.075 $Y=1.23 $X2=0
+ $Y2=0
cc_433 N_A_30_107#_M1007_g N_VGND_c_1317_n 0.0221951f $X=2.155 $Y=0.745 $X2=0
+ $Y2=0
cc_434 N_A_30_107#_M1021_g N_VGND_c_1317_n 0.00176203f $X=6.155 $Y=0.745 $X2=0
+ $Y2=0
cc_435 N_A3_M1002_g N_A1_M1004_g 0.00898703f $X=3.645 $Y=0.745 $X2=0 $Y2=0
cc_436 N_A3_c_572_n N_A1_c_620_n 0.0563623f $X=3.71 $Y=1.585 $X2=0 $Y2=0
cc_437 N_A3_M1009_g A1 5.75519e-19 $X=3.745 $Y=3.345 $X2=0 $Y2=0
cc_438 A3 A1 0.0175662f $X=3.515 $Y=2.32 $X2=0 $Y2=0
cc_439 N_A3_c_577_n A1 0.00273283f $X=3.68 $Y=2.435 $X2=0 $Y2=0
cc_440 N_A3_M1009_g N_A1_c_621_n 0.0144085f $X=3.745 $Y=3.345 $X2=0 $Y2=0
cc_441 A3 N_A1_c_621_n 0.0019765f $X=3.515 $Y=2.32 $X2=0 $Y2=0
cc_442 N_A3_c_573_n N_A1_c_621_n 0.0563623f $X=3.76 $Y=2.25 $X2=0 $Y2=0
cc_443 N_A3_M1009_g N_VPWR_c_934_n 0.0552872f $X=3.745 $Y=3.345 $X2=0 $Y2=0
cc_444 A3 N_VPWR_c_934_n 0.0273827f $X=3.515 $Y=2.32 $X2=0 $Y2=0
cc_445 N_A3_c_577_n N_VPWR_c_934_n 0.00155189f $X=3.68 $Y=2.435 $X2=0 $Y2=0
cc_446 A3 N_VPWR_c_943_n 0.00134527f $X=3.515 $Y=2.32 $X2=0 $Y2=0
cc_447 N_A3_M1002_g N_A_481_107#_c_1027_n 8.64396e-19 $X=3.645 $Y=0.745 $X2=0
+ $Y2=0
cc_448 N_A3_c_572_n N_A_481_107#_c_1030_n 0.0298911f $X=3.71 $Y=1.585 $X2=0
+ $Y2=0
cc_449 N_A3_M1002_g N_A_481_107#_c_1031_n 0.00241201f $X=3.645 $Y=0.745 $X2=0
+ $Y2=0
cc_450 N_A3_M1002_g N_VGND_c_1311_n 0.0436842f $X=3.645 $Y=0.745 $X2=0 $Y2=0
cc_451 N_A3_c_572_n N_VGND_c_1311_n 0.00336273f $X=3.71 $Y=1.585 $X2=0 $Y2=0
cc_452 A1 N_VPWR_c_934_n 0.0076053f $X=4.475 $Y=2.32 $X2=0 $Y2=0
cc_453 N_A1_c_621_n N_VPWR_c_934_n 0.00475791f $X=4.565 $Y=2.47 $X2=0 $Y2=0
cc_454 A1 N_VPWR_c_943_n 0.0158931f $X=4.475 $Y=2.32 $X2=0 $Y2=0
cc_455 N_A1_c_621_n N_VPWR_c_943_n 0.0230935f $X=4.565 $Y=2.47 $X2=0 $Y2=0
cc_456 N_A1_c_620_n N_A_481_107#_c_1030_n 0.014932f $X=4.595 $Y=1.585 $X2=0
+ $Y2=0
cc_457 N_A1_M1004_g N_A_481_107#_c_1031_n 0.0260036f $X=4.665 $Y=0.745 $X2=0
+ $Y2=0
cc_458 N_A1_c_620_n N_A_481_107#_c_1031_n 0.00127977f $X=4.595 $Y=1.585 $X2=0
+ $Y2=0
cc_459 N_A1_M1004_g N_A_481_107#_c_1032_n 0.0162459f $X=4.665 $Y=0.745 $X2=6.24
+ $Y2=0.057
cc_460 N_A1_M1004_g N_A_481_107#_c_1034_n 0.00295244f $X=4.665 $Y=0.745 $X2=6.24
+ $Y2=0.058
cc_461 N_A1_c_621_n N_A_1097_627#_c_1190_n 0.00173957f $X=4.565 $Y=2.47 $X2=0
+ $Y2=0
cc_462 N_A1_M1004_g N_A_1097_627#_c_1209_n 6.17899e-19 $X=4.665 $Y=0.745
+ $X2=12.24 $Y2=0
cc_463 N_A1_M1004_g N_VGND_c_1311_n 0.00197129f $X=4.665 $Y=0.745 $X2=0 $Y2=0
cc_464 N_A1_M1004_g N_VGND_c_1317_n 0.0184926f $X=4.665 $Y=0.745 $X2=0 $Y2=0
cc_465 N_A1_c_620_n N_VGND_c_1317_n 0.00279482f $X=4.595 $Y=1.585 $X2=0 $Y2=0
cc_466 N_A0_c_666_n N_S1_c_720_n 0.0029509f $X=6.81 $Y=2.475 $X2=0 $Y2=0
cc_467 N_A0_M1019_g N_VPWR_c_937_n 0.0495004f $X=6.725 $Y=3.345 $X2=0 $Y2=0
cc_468 N_A0_M1008_g N_A_481_107#_c_1032_n 0.0106132f $X=6.865 $Y=0.745 $X2=6.24
+ $Y2=0.057
cc_469 N_A0_M1008_g N_A_481_107#_c_1087_n 0.0261993f $X=6.865 $Y=0.745 $X2=0
+ $Y2=0
cc_470 N_A0_c_662_n N_A_481_107#_c_1087_n 0.00566423f $X=6.88 $Y=1.35 $X2=0
+ $Y2=0
cc_471 N_A0_c_662_n N_A_481_107#_c_1036_n 0.0161608f $X=6.88 $Y=1.35 $X2=0 $Y2=0
cc_472 A0 N_A_481_107#_c_1036_n 0.0103889f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_473 N_A0_c_662_n N_A_481_107#_c_1105_n 0.00688643f $X=6.88 $Y=1.35 $X2=0
+ $Y2=0
cc_474 A0 N_A_481_107#_c_1105_n 0.0122587f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_475 N_A0_c_662_n N_A_481_107#_c_1037_n 0.00210249f $X=6.88 $Y=1.35 $X2=0
+ $Y2=0
cc_476 N_A0_M1019_g N_A_1097_627#_c_1190_n 3.73432e-19 $X=6.725 $Y=3.345 $X2=0
+ $Y2=0
cc_477 N_A0_M1008_g N_A_1097_627#_c_1209_n 0.0013771f $X=6.865 $Y=0.745
+ $X2=12.24 $Y2=0
cc_478 N_A0_M1019_g N_A_1097_627#_c_1185_n 0.0134366f $X=6.725 $Y=3.345 $X2=0
+ $Y2=0
cc_479 N_A0_M1008_g N_A_1097_627#_c_1185_n 0.0162291f $X=6.865 $Y=0.745 $X2=0
+ $Y2=0
cc_480 N_A0_c_666_n N_A_1097_627#_c_1185_n 0.0167581f $X=6.81 $Y=2.475 $X2=0
+ $Y2=0
cc_481 A0 N_A_1097_627#_c_1185_n 0.0676615f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_482 N_A0_M1019_g N_A_1097_627#_c_1197_n 0.0266156f $X=6.725 $Y=3.345 $X2=0
+ $Y2=0
cc_483 N_A0_c_666_n N_A_1097_627#_c_1197_n 0.00244755f $X=6.81 $Y=2.475 $X2=0
+ $Y2=0
cc_484 A0 N_A_1097_627#_c_1197_n 0.0210044f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_485 N_A0_M1019_g N_A_1097_627#_c_1186_n 0.00659605f $X=6.725 $Y=3.345 $X2=0
+ $Y2=0
cc_486 A0 N_A_1097_627#_c_1186_n 0.0336354f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_487 N_A0_c_663_n N_A_1097_627#_c_1186_n 0.0138973f $X=6.935 $Y=1.95 $X2=0
+ $Y2=0
cc_488 N_A0_M1019_g N_A_1097_627#_c_1199_n 0.00520195f $X=6.725 $Y=3.345 $X2=0
+ $Y2=0
cc_489 A0 N_A_1097_627#_c_1188_n 0.00820559f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_490 N_A0_c_663_n N_A_1097_627#_c_1188_n 0.0040616f $X=6.935 $Y=1.95 $X2=0
+ $Y2=0
cc_491 N_A0_M1019_g N_A_1097_627#_c_1200_n 5.53966e-19 $X=6.725 $Y=3.345 $X2=0
+ $Y2=0
cc_492 N_A0_M1019_g N_A_1097_627#_c_1201_n 0.00508655f $X=6.725 $Y=3.345 $X2=0
+ $Y2=0
cc_493 N_A0_M1019_g N_A_1097_627#_c_1203_n 6.75101e-19 $X=6.725 $Y=3.345 $X2=0
+ $Y2=0
cc_494 N_A0_M1008_g N_VGND_c_1313_n 0.00523047f $X=6.865 $Y=0.745 $X2=0 $Y2=0
cc_495 N_A0_c_662_n N_VGND_c_1313_n 7.21422e-19 $X=6.88 $Y=1.35 $X2=0 $Y2=0
cc_496 N_A0_M1008_g N_VGND_c_1317_n 0.0148881f $X=6.865 $Y=0.745 $X2=0 $Y2=0
cc_497 N_S1_c_704_n N_A_1681_89#_c_791_n 0.0505851f $X=9.435 $Y=1.295 $X2=0
+ $Y2=0
cc_498 N_S1_c_723_p N_A_1681_89#_c_791_n 0.00480283f $X=9.285 $Y=1.48 $X2=0
+ $Y2=0
cc_499 N_S1_c_718_n N_A_1681_89#_c_791_n 0.00769928f $X=9.205 $Y=2.885 $X2=0
+ $Y2=0
cc_500 S1 N_A_1681_89#_c_791_n 0.00966823f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_501 N_S1_M1003_g N_A_1681_89#_M1017_g 0.0283299f $X=8.095 $Y=3.285 $X2=0.24
+ $Y2=0
cc_502 N_S1_c_716_n N_A_1681_89#_M1017_g 0.0198257f $X=9.12 $Y=2.97 $X2=0.24
+ $Y2=0
cc_503 N_S1_M1005_g N_A_1681_89#_M1011_g 0.0260616f $X=9.435 $Y=0.785 $X2=0
+ $Y2=0
cc_504 N_S1_c_704_n N_A_1681_89#_c_798_n 0.0351814f $X=9.435 $Y=1.295 $X2=0
+ $Y2=0
cc_505 N_S1_c_716_n N_A_1681_89#_c_798_n 0.0250285f $X=9.12 $Y=2.97 $X2=0 $Y2=0
cc_506 N_S1_c_718_n N_A_1681_89#_c_798_n 0.0277513f $X=9.205 $Y=2.885 $X2=0
+ $Y2=0
cc_507 S1 N_A_1681_89#_c_798_n 0.00381936f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_508 N_S1_c_720_n N_A_1681_89#_c_798_n 0.0283299f $X=8.03 $Y=2.41 $X2=0 $Y2=0
cc_509 N_S1_M1005_g N_A_1681_89#_c_794_n 0.00268281f $X=9.435 $Y=0.785 $X2=6.24
+ $Y2=0
cc_510 N_S1_c_706_n N_A_1681_89#_c_794_n 0.0428751f $X=10.575 $Y=1.735 $X2=6.24
+ $Y2=0
cc_511 N_S1_c_707_n N_A_1681_89#_c_794_n 0.004986f $X=10.825 $Y=1.485 $X2=6.24
+ $Y2=0
cc_512 N_S1_M1014_g N_A_1681_89#_c_794_n 0.00366474f $X=10.825 $Y=2.425 $X2=6.24
+ $Y2=0
cc_513 N_S1_c_704_n N_A_1681_89#_c_800_n 0.0335234f $X=9.435 $Y=1.295 $X2=6.24
+ $Y2=0.058
cc_514 N_S1_M1014_g N_A_1681_89#_c_800_n 0.00985493f $X=10.825 $Y=2.425 $X2=6.24
+ $Y2=0.058
cc_515 N_S1_c_716_n N_A_1681_89#_c_800_n 0.00472238f $X=9.12 $Y=2.97 $X2=6.24
+ $Y2=0.058
cc_516 N_S1_c_718_n N_A_1681_89#_c_800_n 0.0230069f $X=9.205 $Y=2.885 $X2=6.24
+ $Y2=0.058
cc_517 N_S1_c_742_p N_A_1681_89#_c_800_n 5.71958e-19 $X=9.245 $Y=1.985 $X2=6.24
+ $Y2=0.058
cc_518 N_S1_c_706_n N_A_1681_89#_c_801_n 0.0126009f $X=10.575 $Y=1.735 $X2=0
+ $Y2=0
cc_519 N_S1_M1014_g N_A_1681_89#_c_801_n 0.00405101f $X=10.825 $Y=2.425 $X2=0
+ $Y2=0
cc_520 N_S1_M1003_g N_A_1669_615#_c_867_n 0.0117696f $X=8.095 $Y=3.285 $X2=0
+ $Y2=0
cc_521 N_S1_c_716_n N_A_1669_615#_c_867_n 0.0191209f $X=9.12 $Y=2.97 $X2=0 $Y2=0
cc_522 N_S1_c_716_n N_A_1669_615#_c_868_n 0.0102414f $X=9.12 $Y=2.97 $X2=0.24
+ $Y2=0
cc_523 N_S1_M1005_g N_A_1669_615#_c_882_n 0.0103569f $X=9.435 $Y=0.785 $X2=0
+ $Y2=0
cc_524 N_S1_M1005_g N_A_1669_615#_c_859_n 0.0130516f $X=9.435 $Y=0.785 $X2=12.24
+ $Y2=0
cc_525 N_S1_c_707_n N_A_1669_615#_c_859_n 0.00354091f $X=10.825 $Y=1.485
+ $X2=12.24 $Y2=0
cc_526 N_S1_c_707_n N_A_1669_615#_c_863_n 0.0321564f $X=10.825 $Y=1.485 $X2=0
+ $Y2=0
cc_527 N_S1_c_708_n N_A_1669_615#_c_863_n 0.00537439f $X=10.825 $Y=1.735 $X2=0
+ $Y2=0
cc_528 N_S1_M1014_g N_A_1669_615#_c_874_n 0.0357911f $X=10.825 $Y=2.425 $X2=0
+ $Y2=0
cc_529 N_S1_c_708_n N_A_1669_615#_c_874_n 0.00290907f $X=10.825 $Y=1.735 $X2=0
+ $Y2=0
cc_530 N_S1_c_708_n N_A_1669_615#_c_864_n 0.0300978f $X=10.825 $Y=1.735 $X2=6.24
+ $Y2=0.058
cc_531 N_S1_c_708_n N_A_1669_615#_c_890_n 0.0102103f $X=10.825 $Y=1.735 $X2=0
+ $Y2=0
cc_532 N_S1_c_707_n N_A_1669_615#_M1022_g 0.0396969f $X=10.825 $Y=1.485 $X2=0
+ $Y2=0
cc_533 N_S1_M1003_g N_VPWR_c_937_n 0.00214292f $X=8.095 $Y=3.285 $X2=0 $Y2=0
cc_534 N_S1_M1014_g N_VPWR_c_940_n 0.0216498f $X=10.825 $Y=2.425 $X2=0 $Y2=0
cc_535 N_S1_M1003_g N_VPWR_c_943_n 0.0149982f $X=8.095 $Y=3.285 $X2=0 $Y2=0
cc_536 N_S1_c_716_n N_VPWR_c_943_n 0.020471f $X=9.12 $Y=2.97 $X2=0 $Y2=0
cc_537 N_S1_c_717_n N_VPWR_c_943_n 0.0127062f $X=8.22 $Y=2.97 $X2=0 $Y2=0
cc_538 N_S1_M1005_g N_A_481_107#_c_1108_n 7.80701e-19 $X=9.435 $Y=0.785 $X2=0
+ $Y2=0
cc_539 N_S1_c_704_n N_A_481_107#_c_1042_n 0.00195999f $X=9.435 $Y=1.295 $X2=0
+ $Y2=0
cc_540 N_S1_M1005_g N_A_481_107#_c_1042_n 0.0261592f $X=9.435 $Y=0.785 $X2=0
+ $Y2=0
cc_541 N_S1_c_723_p N_A_481_107#_c_1042_n 0.0182743f $X=9.285 $Y=1.48 $X2=0
+ $Y2=0
cc_542 N_S1_M1005_g N_A_481_107#_c_1044_n 0.0172179f $X=9.435 $Y=0.785 $X2=0
+ $Y2=0
cc_543 N_S1_c_706_n N_A_481_107#_c_1044_n 0.00698756f $X=10.575 $Y=1.735 $X2=0
+ $Y2=0
cc_544 N_S1_c_707_n N_A_481_107#_c_1044_n 0.00282764f $X=10.825 $Y=1.485 $X2=0
+ $Y2=0
cc_545 N_S1_c_704_n N_A_481_107#_c_1045_n 0.0231817f $X=9.435 $Y=1.295 $X2=0
+ $Y2=0
cc_546 N_S1_M1005_g N_A_481_107#_c_1045_n 0.00737747f $X=9.435 $Y=0.785 $X2=0
+ $Y2=0
cc_547 N_S1_c_706_n N_A_481_107#_c_1045_n 0.0149324f $X=10.575 $Y=1.735 $X2=0
+ $Y2=0
cc_548 N_S1_c_716_n N_A_481_107#_c_1045_n 0.0101513f $X=9.12 $Y=2.97 $X2=0 $Y2=0
cc_549 N_S1_c_723_p N_A_481_107#_c_1045_n 0.0446682f $X=9.285 $Y=1.48 $X2=0
+ $Y2=0
cc_550 N_S1_c_718_n N_A_481_107#_c_1045_n 0.0451019f $X=9.205 $Y=2.885 $X2=0
+ $Y2=0
cc_551 S1 N_A_1097_627#_c_1186_n 0.0638838f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_552 N_S1_c_720_n N_A_1097_627#_c_1186_n 0.00286404f $X=8.03 $Y=2.41 $X2=0
+ $Y2=0
cc_553 N_S1_M1003_g N_A_1097_627#_c_1199_n 0.00453588f $X=8.095 $Y=3.285 $X2=0
+ $Y2=0
cc_554 N_S1_c_717_n N_A_1097_627#_c_1199_n 0.00560887f $X=8.22 $Y=2.97 $X2=0
+ $Y2=0
cc_555 N_S1_c_720_n N_A_1097_627#_c_1199_n 8.02962e-19 $X=8.03 $Y=2.41 $X2=0
+ $Y2=0
cc_556 S1 N_A_1097_627#_c_1187_n 0.0333993f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_557 N_S1_c_720_n N_A_1097_627#_c_1187_n 0.00584369f $X=8.03 $Y=2.41 $X2=0
+ $Y2=0
cc_558 N_S1_c_717_n N_A_1097_627#_c_1202_n 0.00269799f $X=8.22 $Y=2.97 $X2=0
+ $Y2=0
cc_559 S1 N_A_1097_627#_c_1202_n 0.0120359f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_560 N_S1_c_720_n N_A_1097_627#_c_1202_n 0.00132778f $X=8.03 $Y=2.41 $X2=0
+ $Y2=0
cc_561 N_S1_M1003_g N_A_1097_627#_c_1203_n 0.0147306f $X=8.095 $Y=3.285 $X2=0
+ $Y2=0
cc_562 N_S1_c_717_n N_A_1097_627#_c_1203_n 0.00285213f $X=8.22 $Y=2.97 $X2=0
+ $Y2=0
cc_563 N_S1_c_707_n N_VGND_c_1315_n 0.0215083f $X=10.825 $Y=1.485 $X2=0 $Y2=0
cc_564 N_S1_M1005_g N_VGND_c_1317_n 0.0123691f $X=9.435 $Y=0.785 $X2=0 $Y2=0
cc_565 N_S1_c_707_n N_VGND_c_1317_n 0.00953929f $X=10.825 $Y=1.485 $X2=0 $Y2=0
cc_566 N_A_1681_89#_M1017_g N_A_1669_615#_c_867_n 0.0166752f $X=8.875 $Y=3.285
+ $X2=0 $Y2=0
cc_567 N_A_1681_89#_M1017_g N_A_1669_615#_c_868_n 0.013865f $X=8.875 $Y=3.285
+ $X2=0.24 $Y2=0
cc_568 N_A_1681_89#_c_800_n N_A_1669_615#_c_868_n 0.0117988f $X=9.985 $Y=2.41
+ $X2=0.24 $Y2=0
cc_569 N_A_1681_89#_M1011_g N_A_1669_615#_c_882_n 0.00681521f $X=8.655 $Y=0.785
+ $X2=0 $Y2=0
cc_570 N_A_1681_89#_c_794_n N_A_1669_615#_c_859_n 0.00576468f $X=10.435 $Y=1.165
+ $X2=12.24 $Y2=0
cc_571 N_A_1681_89#_c_794_n N_A_1669_615#_c_863_n 0.031397f $X=10.435 $Y=1.165
+ $X2=0 $Y2=0
cc_572 N_A_1681_89#_c_794_n N_A_1669_615#_c_874_n 0.0130894f $X=10.435 $Y=1.165
+ $X2=0 $Y2=0
cc_573 N_A_1681_89#_c_800_n N_A_1669_615#_c_874_n 0.00456787f $X=9.985 $Y=2.41
+ $X2=0 $Y2=0
cc_574 N_A_1681_89#_c_801_n N_A_1669_615#_c_874_n 0.0302701f $X=10.435 $Y=2.425
+ $X2=0 $Y2=0
cc_575 N_A_1681_89#_c_794_n N_A_1669_615#_c_890_n 0.0246602f $X=10.435 $Y=1.165
+ $X2=0 $Y2=0
cc_576 N_A_1681_89#_M1017_g N_VPWR_c_943_n 0.015893f $X=8.875 $Y=3.285 $X2=0
+ $Y2=0
cc_577 N_A_1681_89#_c_800_n N_VPWR_c_943_n 0.0143692f $X=9.985 $Y=2.41 $X2=0
+ $Y2=0
cc_578 N_A_1681_89#_c_801_n N_VPWR_c_943_n 0.00918248f $X=10.435 $Y=2.425 $X2=0
+ $Y2=0
cc_579 N_A_1681_89#_M1011_g N_A_481_107#_c_1037_n 0.00294814f $X=8.655 $Y=0.785
+ $X2=0 $Y2=0
cc_580 N_A_1681_89#_M1011_g N_A_481_107#_c_1038_n 0.0049279f $X=8.655 $Y=0.785
+ $X2=0 $Y2=0
cc_581 N_A_1681_89#_M1011_g N_A_481_107#_c_1108_n 0.0226054f $X=8.655 $Y=0.785
+ $X2=0 $Y2=0
cc_582 N_A_1681_89#_c_791_n N_A_481_107#_c_1042_n 0.00927075f $X=8.765 $Y=2.225
+ $X2=0 $Y2=0
cc_583 N_A_1681_89#_M1011_g N_A_481_107#_c_1042_n 0.0084731f $X=8.655 $Y=0.785
+ $X2=0 $Y2=0
cc_584 N_A_1681_89#_c_791_n N_A_481_107#_c_1043_n 0.00410234f $X=8.765 $Y=2.225
+ $X2=0 $Y2=0
cc_585 N_A_1681_89#_M1011_g N_A_481_107#_c_1043_n 0.00528128f $X=8.655 $Y=0.785
+ $X2=0 $Y2=0
cc_586 N_A_1681_89#_M1011_g N_A_481_107#_c_1044_n 4.54677e-19 $X=8.655 $Y=0.785
+ $X2=0 $Y2=0
cc_587 N_A_1681_89#_c_794_n N_A_481_107#_c_1044_n 0.0110743f $X=10.435 $Y=1.165
+ $X2=0 $Y2=0
cc_588 N_A_1681_89#_c_791_n N_A_481_107#_c_1045_n 7.35739e-19 $X=8.765 $Y=2.225
+ $X2=0 $Y2=0
cc_589 N_A_1681_89#_M1017_g N_A_481_107#_c_1045_n 0.00230334f $X=8.875 $Y=3.285
+ $X2=0 $Y2=0
cc_590 N_A_1681_89#_c_794_n N_A_481_107#_c_1045_n 0.029778f $X=10.435 $Y=1.165
+ $X2=0 $Y2=0
cc_591 N_A_1681_89#_c_800_n N_A_481_107#_c_1045_n 0.0402007f $X=9.985 $Y=2.41
+ $X2=0 $Y2=0
cc_592 N_A_1681_89#_c_801_n N_A_481_107#_c_1045_n 0.0573273f $X=10.435 $Y=2.425
+ $X2=0 $Y2=0
cc_593 N_A_1681_89#_M1017_g N_A_481_107#_c_1049_n 0.0118481f $X=8.875 $Y=3.285
+ $X2=0 $Y2=0
cc_594 N_A_1681_89#_c_800_n N_A_481_107#_c_1049_n 0.00704358f $X=9.985 $Y=2.41
+ $X2=0 $Y2=0
cc_595 N_A_1681_89#_c_791_n N_A_1097_627#_c_1187_n 0.0066383f $X=8.765 $Y=2.225
+ $X2=0 $Y2=0
cc_596 N_A_1681_89#_c_791_n N_A_1097_627#_c_1189_n 0.0143501f $X=8.765 $Y=2.225
+ $X2=0 $Y2=0
cc_597 N_A_1681_89#_M1011_g N_A_1097_627#_c_1189_n 0.0039825f $X=8.655 $Y=0.785
+ $X2=0 $Y2=0
cc_598 N_A_1681_89#_M1011_g N_VGND_c_1317_n 0.013659f $X=8.655 $Y=0.785 $X2=0
+ $Y2=0
cc_599 N_A_1681_89#_c_794_n N_VGND_c_1317_n 0.00786189f $X=10.435 $Y=1.165 $X2=0
+ $Y2=0
cc_600 N_A_1669_615#_c_868_n N_VPWR_c_940_n 0.00839908f $X=10.7 $Y=3.72 $X2=0
+ $Y2=0
cc_601 N_A_1669_615#_c_874_n N_VPWR_c_940_n 0.110572f $X=10.785 $Y=3.635 $X2=0
+ $Y2=0
cc_602 N_A_1669_615#_c_864_n N_VPWR_c_940_n 0.0549914f $X=11.75 $Y=1.76 $X2=0
+ $Y2=0
cc_603 N_A_1669_615#_M1022_g N_VPWR_c_940_n 0.11059f $X=11.815 $Y=1 $X2=0 $Y2=0
cc_604 N_A_1669_615#_c_867_n N_VPWR_c_943_n 0.0218836f $X=8.485 $Y=3.345 $X2=0
+ $Y2=0
cc_605 N_A_1669_615#_c_868_n N_VPWR_c_943_n 0.0929115f $X=10.7 $Y=3.72 $X2=0
+ $Y2=0
cc_606 N_A_1669_615#_c_871_n N_VPWR_c_943_n 0.0128157f $X=8.65 $Y=3.72 $X2=0
+ $Y2=0
cc_607 N_A_1669_615#_c_874_n N_VPWR_c_943_n 0.0216909f $X=10.785 $Y=3.635 $X2=0
+ $Y2=0
cc_608 N_A_1669_615#_M1022_g N_VPWR_c_943_n 0.00914225f $X=11.815 $Y=1 $X2=0
+ $Y2=0
cc_609 N_A_1669_615#_c_861_n N_A_481_107#_c_1038_n 0.0119651f $X=9.21 $Y=0.35
+ $X2=0 $Y2=0
cc_610 N_A_1669_615#_c_882_n N_A_481_107#_c_1108_n 0.0225117f $X=9.045 $Y=0.7
+ $X2=0 $Y2=0
cc_611 N_A_1669_615#_M1011_d N_A_481_107#_c_1042_n 0.00171693f $X=8.905 $Y=0.575
+ $X2=0 $Y2=0
cc_612 N_A_1669_615#_c_882_n N_A_481_107#_c_1042_n 0.015004f $X=9.045 $Y=0.7
+ $X2=0 $Y2=0
cc_613 N_A_1669_615#_c_859_n N_A_481_107#_c_1042_n 0.00573334f $X=10.7 $Y=0.35
+ $X2=0 $Y2=0
cc_614 N_A_1669_615#_c_882_n N_A_481_107#_c_1044_n 0.00735258f $X=9.045 $Y=0.7
+ $X2=0 $Y2=0
cc_615 N_A_1669_615#_c_859_n N_A_481_107#_c_1044_n 0.0281924f $X=10.7 $Y=0.35
+ $X2=0 $Y2=0
cc_616 N_A_1669_615#_c_868_n N_A_481_107#_c_1049_n 0.0219235f $X=10.7 $Y=3.72
+ $X2=0 $Y2=0
cc_617 N_A_1669_615#_c_867_n N_A_1097_627#_c_1203_n 0.00897547f $X=8.485
+ $Y=3.345 $X2=0 $Y2=0
cc_618 N_A_1669_615#_c_864_n N_X_c_1296_n 0.0233946f $X=11.75 $Y=1.76 $X2=0
+ $Y2=0
cc_619 N_A_1669_615#_M1022_g N_X_c_1296_n 0.0358732f $X=11.815 $Y=1 $X2=0 $Y2=0
cc_620 N_A_1669_615#_c_859_n N_VGND_c_1315_n 0.00489946f $X=10.7 $Y=0.35 $X2=0
+ $Y2=0
cc_621 N_A_1669_615#_c_863_n N_VGND_c_1315_n 0.0717942f $X=10.785 $Y=1.595 $X2=0
+ $Y2=0
cc_622 N_A_1669_615#_c_864_n N_VGND_c_1315_n 0.0701333f $X=11.75 $Y=1.76 $X2=0
+ $Y2=0
cc_623 N_A_1669_615#_M1022_g N_VGND_c_1315_n 0.059832f $X=11.815 $Y=1 $X2=0
+ $Y2=0
cc_624 N_A_1669_615#_c_882_n N_VGND_c_1317_n 0.0187582f $X=9.045 $Y=0.7 $X2=0
+ $Y2=0
cc_625 N_A_1669_615#_c_859_n N_VGND_c_1317_n 0.0649911f $X=10.7 $Y=0.35 $X2=0
+ $Y2=0
cc_626 N_A_1669_615#_c_861_n N_VGND_c_1317_n 0.00868351f $X=9.21 $Y=0.35 $X2=0
+ $Y2=0
cc_627 N_A_1669_615#_c_863_n N_VGND_c_1317_n 0.0167622f $X=10.785 $Y=1.595 $X2=0
+ $Y2=0
cc_628 N_A_1669_615#_M1022_g N_VGND_c_1317_n 0.00886025f $X=11.815 $Y=1 $X2=0
+ $Y2=0
cc_629 N_VPWR_c_943_n A_339_627# 0.00871617f $X=11.855 $Y=3.59 $X2=0 $Y2=3.985
cc_630 N_VPWR_c_943_n N_A_481_107#_M1017_d 0.00543808f $X=11.855 $Y=3.59
+ $X2=-0.33 $Y2=1.885
cc_631 N_VPWR_c_943_n N_A_481_107#_c_1029_n 5.69188e-19 $X=11.855 $Y=3.59
+ $X2=6.24 $Y2=4.012
cc_632 N_VPWR_c_943_n N_A_481_107#_c_1071_n 0.0161284f $X=11.855 $Y=3.59 $X2=0
+ $Y2=0
cc_633 N_VPWR_c_943_n N_A_481_107#_c_1049_n 0.0137798f $X=11.855 $Y=3.59 $X2=0
+ $Y2=0
cc_634 N_VPWR_c_934_n A_637_627# 0.00455105f $X=4.135 $Y=3.345 $X2=0 $Y2=3.985
cc_635 N_VPWR_c_943_n A_637_627# 0.00354485f $X=11.855 $Y=3.59 $X2=0 $Y2=3.985
cc_636 N_VPWR_c_943_n A_955_627# 0.00875788f $X=11.855 $Y=3.59 $X2=0 $Y2=3.985
cc_637 N_VPWR_c_937_n N_A_1097_627#_c_1190_n 0.014128f $X=7.165 $Y=3.59
+ $X2=12.24 $Y2=4.07
cc_638 N_VPWR_c_943_n N_A_1097_627#_c_1191_n 0.0352842f $X=11.855 $Y=3.59
+ $X2=12.24 $Y2=4.07
cc_639 N_VPWR_c_937_n N_A_1097_627#_c_1194_n 0.00693017f $X=7.165 $Y=3.59 $X2=0
+ $Y2=0
cc_640 N_VPWR_c_943_n N_A_1097_627#_c_1194_n 0.0160931f $X=11.855 $Y=3.59 $X2=0
+ $Y2=0
cc_641 N_VPWR_c_937_n N_A_1097_627#_c_1197_n 0.0502699f $X=7.165 $Y=3.59 $X2=0
+ $Y2=0
cc_642 N_VPWR_c_943_n N_A_1097_627#_c_1197_n 0.0087779f $X=11.855 $Y=3.59 $X2=0
+ $Y2=0
cc_643 N_VPWR_c_937_n N_A_1097_627#_c_1199_n 0.00154098f $X=7.165 $Y=3.59 $X2=0
+ $Y2=0
cc_644 N_VPWR_c_943_n N_A_1097_627#_c_1199_n 4.93401e-19 $X=11.855 $Y=3.59 $X2=0
+ $Y2=0
cc_645 N_VPWR_c_937_n N_A_1097_627#_c_1201_n 0.0134642f $X=7.165 $Y=3.59 $X2=0
+ $Y2=0
cc_646 N_VPWR_c_943_n N_A_1097_627#_c_1201_n 6.61476e-19 $X=11.855 $Y=3.59 $X2=0
+ $Y2=0
cc_647 N_VPWR_c_937_n N_A_1097_627#_c_1203_n 0.0347251f $X=7.165 $Y=3.59 $X2=0
+ $Y2=0
cc_648 N_VPWR_c_943_n N_A_1097_627#_c_1203_n 0.0266379f $X=11.855 $Y=3.59 $X2=0
+ $Y2=0
cc_649 N_VPWR_c_937_n A_1253_627# 0.00557635f $X=7.165 $Y=3.59 $X2=0 $Y2=3.985
cc_650 N_VPWR_c_943_n A_1253_627# 8.67137e-19 $X=11.855 $Y=3.59 $X2=0 $Y2=3.985
cc_651 N_VPWR_c_943_n N_X_M1015_d 0.00221032f $X=11.855 $Y=3.59 $X2=0 $Y2=0
cc_652 N_VPWR_c_940_n N_X_c_1296_n 0.0664963f $X=11.33 $Y=2.34 $X2=6.24 $Y2=4.07
cc_653 N_VPWR_c_943_n N_X_c_1296_n 0.0341921f $X=11.855 $Y=3.59 $X2=6.24
+ $Y2=4.07
cc_654 N_A_481_107#_c_1032_n N_A_1097_627#_c_1209_n 0.0597316f $X=6.77 $Y=0.35
+ $X2=12.24 $Y2=0
cc_655 N_A_481_107#_c_1087_n N_A_1097_627#_c_1209_n 0.00991117f $X=6.855
+ $Y=1.175 $X2=12.24 $Y2=0
cc_656 N_A_481_107#_c_1087_n N_A_1097_627#_c_1185_n 0.0162652f $X=6.855 $Y=1.175
+ $X2=0 $Y2=0
cc_657 N_A_481_107#_c_1105_n N_A_1097_627#_c_1185_n 0.0130053f $X=6.94 $Y=1.26
+ $X2=0 $Y2=0
cc_658 N_A_481_107#_c_1036_n N_A_1097_627#_c_1187_n 0.0241093f $X=7.83 $Y=1.26
+ $X2=0 $Y2=0
cc_659 N_A_481_107#_c_1036_n N_A_1097_627#_c_1188_n 0.0117907f $X=7.83 $Y=1.26
+ $X2=0 $Y2=0
cc_660 N_A_481_107#_c_1036_n N_A_1097_627#_c_1189_n 0.0137879f $X=7.83 $Y=1.26
+ $X2=0 $Y2=0
cc_661 N_A_481_107#_c_1037_n N_A_1097_627#_c_1189_n 0.0398982f $X=7.915 $Y=1.175
+ $X2=0 $Y2=0
cc_662 N_A_481_107#_c_1038_n N_A_1097_627#_c_1189_n 0.0112524f $X=8.53 $Y=0.35
+ $X2=0 $Y2=0
cc_663 N_A_481_107#_c_1108_n N_A_1097_627#_c_1189_n 0.0114451f $X=8.615 $Y=0.965
+ $X2=0 $Y2=0
cc_664 N_A_481_107#_c_1043_n N_A_1097_627#_c_1189_n 0.0119269f $X=8.7 $Y=1.05
+ $X2=0 $Y2=0
cc_665 N_A_481_107#_c_1027_n N_VGND_c_1311_n 0.0118393f $X=2.545 $Y=0.745 $X2=0
+ $Y2=0
cc_666 N_A_481_107#_c_1030_n N_VGND_c_1311_n 0.0623437f $X=4.38 $Y=1.18 $X2=0
+ $Y2=0
cc_667 N_A_481_107#_c_1031_n N_VGND_c_1311_n 0.0237468f $X=4.465 $Y=1.095 $X2=0
+ $Y2=0
cc_668 N_A_481_107#_c_1034_n N_VGND_c_1311_n 0.00485641f $X=4.55 $Y=0.35 $X2=0
+ $Y2=0
cc_669 N_A_481_107#_c_1032_n N_VGND_c_1313_n 0.00476005f $X=6.77 $Y=0.35 $X2=0
+ $Y2=0
cc_670 N_A_481_107#_c_1087_n N_VGND_c_1313_n 0.0243957f $X=6.855 $Y=1.175 $X2=0
+ $Y2=0
cc_671 N_A_481_107#_c_1036_n N_VGND_c_1313_n 0.041168f $X=7.83 $Y=1.26 $X2=0
+ $Y2=0
cc_672 N_A_481_107#_c_1037_n N_VGND_c_1313_n 0.0421329f $X=7.915 $Y=1.175 $X2=0
+ $Y2=0
cc_673 N_A_481_107#_c_1040_n N_VGND_c_1313_n 0.00488019f $X=8 $Y=0.35 $X2=0
+ $Y2=0
cc_674 N_A_481_107#_c_1027_n N_VGND_c_1317_n 0.0388338f $X=2.545 $Y=0.745 $X2=0
+ $Y2=0
cc_675 N_A_481_107#_c_1030_n N_VGND_c_1317_n 0.0267461f $X=4.38 $Y=1.18 $X2=0
+ $Y2=0
cc_676 N_A_481_107#_c_1031_n N_VGND_c_1317_n 0.0193536f $X=4.465 $Y=1.095 $X2=0
+ $Y2=0
cc_677 N_A_481_107#_c_1032_n N_VGND_c_1317_n 0.0830365f $X=6.77 $Y=0.35 $X2=0
+ $Y2=0
cc_678 N_A_481_107#_c_1034_n N_VGND_c_1317_n 0.0077932f $X=4.55 $Y=0.35 $X2=0
+ $Y2=0
cc_679 N_A_481_107#_c_1087_n N_VGND_c_1317_n 0.0199529f $X=6.855 $Y=1.175 $X2=0
+ $Y2=0
cc_680 N_A_481_107#_c_1036_n N_VGND_c_1317_n 0.013131f $X=7.83 $Y=1.26 $X2=0
+ $Y2=0
cc_681 N_A_481_107#_c_1037_n N_VGND_c_1317_n 0.0194693f $X=7.915 $Y=1.175 $X2=0
+ $Y2=0
cc_682 N_A_481_107#_c_1038_n N_VGND_c_1317_n 0.0280262f $X=8.53 $Y=0.35 $X2=0
+ $Y2=0
cc_683 N_A_481_107#_c_1040_n N_VGND_c_1317_n 0.00777234f $X=8 $Y=0.35 $X2=0
+ $Y2=0
cc_684 N_A_481_107#_c_1108_n N_VGND_c_1317_n 0.0182656f $X=8.615 $Y=0.965 $X2=0
+ $Y2=0
cc_685 N_A_481_107#_c_1042_n N_VGND_c_1317_n 0.0160506f $X=9.55 $Y=1.05 $X2=0
+ $Y2=0
cc_686 N_A_481_107#_c_1044_n N_VGND_c_1317_n 0.0291924f $X=9.635 $Y=1.135 $X2=0
+ $Y2=0
cc_687 N_A_1097_627#_M1011_s N_VGND_c_1317_n 0.00479598f $X=8.12 $Y=0.575 $X2=0
+ $Y2=0
cc_688 N_A_1097_627#_c_1209_n N_VGND_c_1317_n 0.0498389f $X=6.42 $Y=0.765 $X2=0
+ $Y2=0
cc_689 N_A_1097_627#_c_1189_n N_VGND_c_1317_n 0.0117486f $X=8.265 $Y=0.825 $X2=0
+ $Y2=0
cc_690 N_A_1097_627#_c_1209_n A_1281_107# 4.80934e-19 $X=6.42 $Y=0.765 $X2=0
+ $Y2=0
cc_691 N_X_c_1296_n N_VGND_c_1315_n 0.0344049f $X=12.205 $Y=0.77 $X2=0 $Y2=0
cc_692 N_X_M1022_d N_VGND_c_1317_n 0.00221032f $X=12.065 $Y=0.625 $X2=0 $Y2=0
cc_693 N_X_c_1296_n N_VGND_c_1317_n 0.0204166f $X=12.205 $Y=0.77 $X2=0 $Y2=0
cc_694 N_VGND_c_1317_n A_339_107# 0.00286287f $X=11.855 $Y=0.48 $X2=0 $Y2=0
cc_695 N_VGND_c_1311_n A_637_107# 0.00604574f $X=4.085 $Y=0.48 $X2=0 $Y2=0
cc_696 N_VGND_c_1317_n A_637_107# 8.10341e-19 $X=11.855 $Y=0.48 $X2=0 $Y2=0
cc_697 N_VGND_c_1317_n A_983_107# 0.00220765f $X=11.855 $Y=0.48 $X2=0 $Y2=0
cc_698 N_VGND_c_1317_n A_1281_107# 0.0010009f $X=11.855 $Y=0.48 $X2=0 $Y2=0
