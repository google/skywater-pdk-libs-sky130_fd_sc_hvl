# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__dfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__dfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.00000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595000 1.555000 2.470000 1.750000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.560000 2.185000 11.890000 3.735000 ;
        RECT 11.640000 0.685000 11.890000 2.185000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.540000 1.905000 0.870000 2.575000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.560000 0.365000  1.510000 1.095000 ;
        RECT  2.200000 0.365000  2.765000 1.025000 ;
        RECT  5.255000 0.365000  6.205000 0.995000 ;
        RECT  8.780000 0.365000  9.730000 1.245000 ;
        RECT 10.690000 0.365000 11.280000 1.495000 ;
      LAYER mcon ;
        RECT  0.590000 0.395000  0.760000 0.565000 ;
        RECT  0.950000 0.395000  1.120000 0.565000 ;
        RECT  1.310000 0.395000  1.480000 0.565000 ;
        RECT  2.215000 0.395000  2.385000 0.565000 ;
        RECT  2.575000 0.395000  2.745000 0.565000 ;
        RECT  5.285000 0.395000  5.455000 0.565000 ;
        RECT  5.645000 0.395000  5.815000 0.565000 ;
        RECT  6.005000 0.395000  6.175000 0.565000 ;
        RECT  8.810000 0.395000  8.980000 0.565000 ;
        RECT  9.170000 0.395000  9.340000 0.565000 ;
        RECT  9.530000 0.395000  9.700000 0.565000 ;
        RECT 10.720000 0.395000 10.890000 0.565000 ;
        RECT 11.080000 0.395000 11.250000 0.565000 ;
      LAYER met1 ;
        RECT 0.000000 0.255000 12.000000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 12.000000 0.085000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.115000 12.000000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 12.000000 4.155000 ;
      LAYER mcon ;
        RECT  0.155000 3.985000  0.325000 4.155000 ;
        RECT  0.635000 3.985000  0.805000 4.155000 ;
        RECT  1.115000 3.985000  1.285000 4.155000 ;
        RECT  1.595000 3.985000  1.765000 4.155000 ;
        RECT  2.075000 3.985000  2.245000 4.155000 ;
        RECT  2.555000 3.985000  2.725000 4.155000 ;
        RECT  3.035000 3.985000  3.205000 4.155000 ;
        RECT  3.515000 3.985000  3.685000 4.155000 ;
        RECT  3.995000 3.985000  4.165000 4.155000 ;
        RECT  4.475000 3.985000  4.645000 4.155000 ;
        RECT  4.955000 3.985000  5.125000 4.155000 ;
        RECT  5.435000 3.985000  5.605000 4.155000 ;
        RECT  5.915000 3.985000  6.085000 4.155000 ;
        RECT  6.395000 3.985000  6.565000 4.155000 ;
        RECT  6.875000 3.985000  7.045000 4.155000 ;
        RECT  7.355000 3.985000  7.525000 4.155000 ;
        RECT  7.835000 3.985000  8.005000 4.155000 ;
        RECT  8.315000 3.985000  8.485000 4.155000 ;
        RECT  8.795000 3.985000  8.965000 4.155000 ;
        RECT  9.275000 3.985000  9.445000 4.155000 ;
        RECT  9.755000 3.985000  9.925000 4.155000 ;
        RECT 10.235000 3.985000 10.405000 4.155000 ;
        RECT 10.715000 3.985000 10.885000 4.155000 ;
        RECT 11.195000 3.985000 11.365000 4.155000 ;
        RECT 11.675000 3.985000 11.845000 4.155000 ;
      LAYER met1 ;
        RECT 0.000000 3.955000 12.000000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.540000 2.755000  1.490000 3.705000 ;
        RECT  2.220000 2.795000  2.470000 3.705000 ;
        RECT  5.070000 3.485000  6.020000 3.735000 ;
        RECT  8.815000 2.695000  9.765000 3.735000 ;
        RECT 10.725000 2.195000 11.315000 3.735000 ;
      LAYER mcon ;
        RECT  0.570000 3.505000  0.740000 3.675000 ;
        RECT  0.930000 3.505000  1.100000 3.675000 ;
        RECT  1.290000 3.505000  1.460000 3.675000 ;
        RECT  2.250000 3.505000  2.420000 3.675000 ;
        RECT  5.100000 3.515000  5.270000 3.685000 ;
        RECT  5.460000 3.515000  5.630000 3.685000 ;
        RECT  5.820000 3.515000  5.990000 3.685000 ;
        RECT  8.845000 3.505000  9.015000 3.675000 ;
        RECT  9.205000 3.505000  9.375000 3.675000 ;
        RECT  9.565000 3.505000  9.735000 3.675000 ;
        RECT 10.755000 3.505000 10.925000 3.675000 ;
        RECT 11.115000 3.505000 11.285000 3.675000 ;
      LAYER met1 ;
        RECT 0.000000 3.445000 12.000000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.110000 0.595000  0.380000 1.555000 ;
      RECT  0.110000 1.555000  1.415000 1.725000 ;
      RECT  0.110000 1.725000  0.360000 3.565000 ;
      RECT  1.165000 1.725000  1.415000 1.930000 ;
      RECT  1.165000 1.930000  2.820000 2.225000 ;
      RECT  1.670000 2.445000  2.820000 2.615000 ;
      RECT  1.670000 2.615000  2.000000 3.565000 ;
      RECT  1.690000 0.595000  2.020000 1.205000 ;
      RECT  1.690000 1.205000  3.115000 1.375000 ;
      RECT  2.650000 1.760000  3.685000 1.930000 ;
      RECT  2.650000 2.615000  2.820000 3.305000 ;
      RECT  2.650000 3.305000  3.680000 3.475000 ;
      RECT  2.945000 0.265000  5.055000 0.435000 ;
      RECT  2.945000 0.435000  3.115000 1.205000 ;
      RECT  3.000000 2.110000  4.035000 2.280000 ;
      RECT  3.000000 2.280000  3.330000 3.125000 ;
      RECT  3.295000 0.615000  4.035000 1.025000 ;
      RECT  3.430000 1.205000  3.685000 1.760000 ;
      RECT  3.510000 2.460000  3.840000 3.135000 ;
      RECT  3.510000 3.135000  7.655000 3.305000 ;
      RECT  3.865000 1.025000  4.035000 2.110000 ;
      RECT  4.055000 2.675000  4.385000 2.955000 ;
      RECT  4.215000 0.615000  4.545000 1.525000 ;
      RECT  4.215000 1.525000  6.345000 1.695000 ;
      RECT  4.215000 1.695000  4.385000 2.675000 ;
      RECT  4.565000 1.885000  4.890000 2.385000 ;
      RECT  4.565000 2.385000  6.955000 2.555000 ;
      RECT  4.725000 0.435000  5.055000 1.175000 ;
      RECT  4.725000 1.175000  6.555000 1.345000 ;
      RECT  5.435000 1.875000  7.305000 2.045000 ;
      RECT  5.435000 2.045000  5.765000 2.205000 ;
      RECT  6.385000 0.265000  7.450000 0.435000 ;
      RECT  6.385000 0.435000  6.555000 1.175000 ;
      RECT  6.470000 2.755000  7.305000 2.955000 ;
      RECT  6.705000 2.225000  6.955000 2.385000 ;
      RECT  6.735000 0.615000  7.065000 1.875000 ;
      RECT  7.135000 2.045000  7.305000 2.755000 ;
      RECT  7.280000 0.435000  7.450000 1.125000 ;
      RECT  7.280000 1.125000  7.655000 1.445000 ;
      RECT  7.485000 1.445000  7.655000 2.225000 ;
      RECT  7.485000 2.225000  8.250000 2.515000 ;
      RECT  7.485000 2.515000  7.655000 3.135000 ;
      RECT  7.630000 0.525000  8.005000 0.855000 ;
      RECT  7.630000 0.855000  8.600000 0.945000 ;
      RECT  7.835000 0.945000  8.600000 1.025000 ;
      RECT  7.835000 2.695000  8.600000 2.865000 ;
      RECT  7.835000 2.865000  8.085000 3.735000 ;
      RECT  8.430000 1.025000  8.600000 2.275000 ;
      RECT  8.430000 2.275000 10.035000 2.445000 ;
      RECT  8.430000 2.445000  8.600000 2.695000 ;
      RECT  9.000000 1.425000 10.510000 1.595000 ;
      RECT  9.000000 1.595000  9.330000 2.015000 ;
      RECT  9.705000 1.775000 10.035000 2.275000 ;
      RECT 10.180000 0.525000 10.510000 1.425000 ;
      RECT 10.215000 1.595000 10.510000 1.675000 ;
      RECT 10.215000 1.675000 11.460000 2.005000 ;
      RECT 10.215000 2.005000 10.545000 3.735000 ;
  END
END sky130_fd_sc_hvl__dfxtp_1
