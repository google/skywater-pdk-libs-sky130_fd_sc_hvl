# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__dfstp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__dfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.88000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.525000 2.835000 2.095000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.478750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.420000 0.645000 14.770000 3.615000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.165000 1.555000  8.100000 1.795000 ;
        RECT  7.930000 0.840000 11.160000 1.010000 ;
        RECT  7.930000 1.010000  8.100000 1.555000 ;
        RECT  8.285000 0.555000 11.160000 0.840000 ;
        RECT 10.885000 1.010000 11.160000 1.040000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.545000 2.075000 0.875000 2.745000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.570000 0.365000  1.160000 1.115000 ;
        RECT  2.470000 0.365000  3.005000 0.995000 ;
        RECT  4.855000 0.365000  5.805000 0.785000 ;
        RECT  6.800000 0.365000  7.750000 1.375000 ;
        RECT 11.340000 0.365000 11.930000 1.475000 ;
        RECT 13.255000 0.365000 14.205000 1.475000 ;
      LAYER mcon ;
        RECT  0.600000 0.395000  0.770000 0.565000 ;
        RECT  0.960000 0.395000  1.130000 0.565000 ;
        RECT  2.470000 0.395000  2.640000 0.565000 ;
        RECT  2.830000 0.395000  3.000000 0.565000 ;
        RECT  4.885000 0.395000  5.055000 0.565000 ;
        RECT  5.245000 0.395000  5.415000 0.565000 ;
        RECT  5.605000 0.395000  5.775000 0.565000 ;
        RECT  6.830000 0.395000  7.000000 0.565000 ;
        RECT  7.190000 0.395000  7.360000 0.565000 ;
        RECT  7.550000 0.395000  7.720000 0.565000 ;
        RECT 11.370000 0.395000 11.540000 0.565000 ;
        RECT 11.730000 0.395000 11.900000 0.565000 ;
        RECT 13.285000 0.395000 13.455000 0.565000 ;
        RECT 13.645000 0.395000 13.815000 0.565000 ;
        RECT 14.005000 0.395000 14.175000 0.565000 ;
      LAYER met1 ;
        RECT 0.000000 0.255000 14.880000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 14.880000 0.085000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.115000 14.880000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 14.880000 4.155000 ;
      LAYER mcon ;
        RECT  0.155000 3.985000  0.325000 4.155000 ;
        RECT  0.635000 3.985000  0.805000 4.155000 ;
        RECT  1.115000 3.985000  1.285000 4.155000 ;
        RECT  1.595000 3.985000  1.765000 4.155000 ;
        RECT  2.075000 3.985000  2.245000 4.155000 ;
        RECT  2.555000 3.985000  2.725000 4.155000 ;
        RECT  3.035000 3.985000  3.205000 4.155000 ;
        RECT  3.515000 3.985000  3.685000 4.155000 ;
        RECT  3.995000 3.985000  4.165000 4.155000 ;
        RECT  4.475000 3.985000  4.645000 4.155000 ;
        RECT  4.955000 3.985000  5.125000 4.155000 ;
        RECT  5.435000 3.985000  5.605000 4.155000 ;
        RECT  5.915000 3.985000  6.085000 4.155000 ;
        RECT  6.395000 3.985000  6.565000 4.155000 ;
        RECT  6.875000 3.985000  7.045000 4.155000 ;
        RECT  7.355000 3.985000  7.525000 4.155000 ;
        RECT  7.835000 3.985000  8.005000 4.155000 ;
        RECT  8.315000 3.985000  8.485000 4.155000 ;
        RECT  8.795000 3.985000  8.965000 4.155000 ;
        RECT  9.275000 3.985000  9.445000 4.155000 ;
        RECT  9.755000 3.985000  9.925000 4.155000 ;
        RECT 10.235000 3.985000 10.405000 4.155000 ;
        RECT 10.715000 3.985000 10.885000 4.155000 ;
        RECT 11.195000 3.985000 11.365000 4.155000 ;
        RECT 11.675000 3.985000 11.845000 4.155000 ;
        RECT 12.155000 3.985000 12.325000 4.155000 ;
        RECT 12.635000 3.985000 12.805000 4.155000 ;
        RECT 13.115000 3.985000 13.285000 4.155000 ;
        RECT 13.595000 3.985000 13.765000 4.155000 ;
        RECT 14.075000 3.985000 14.245000 4.155000 ;
        RECT 14.555000 3.985000 14.725000 4.155000 ;
      LAYER met1 ;
        RECT 0.000000 3.955000 14.880000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.545000 2.925000  1.495000 3.755000 ;
        RECT  2.235000 2.625000  2.485000 3.705000 ;
        RECT  5.605000 2.855000  5.935000 3.705000 ;
        RECT  7.075000 2.675000  8.025000 3.705000 ;
        RECT 10.010000 2.665000 10.960000 3.705000 ;
        RECT 11.730000 3.355000 12.680000 3.735000 ;
        RECT 13.295000 2.575000 14.240000 3.705000 ;
      LAYER mcon ;
        RECT  0.575000 3.505000  0.745000 3.675000 ;
        RECT  0.935000 3.505000  1.105000 3.675000 ;
        RECT  1.295000 3.505000  1.465000 3.675000 ;
        RECT  2.265000 3.505000  2.435000 3.675000 ;
        RECT  5.635000 3.505000  5.805000 3.675000 ;
        RECT  7.105000 3.505000  7.275000 3.675000 ;
        RECT  7.465000 3.505000  7.635000 3.675000 ;
        RECT  7.825000 3.505000  7.995000 3.675000 ;
        RECT 10.040000 3.505000 10.210000 3.675000 ;
        RECT 10.400000 3.505000 10.570000 3.675000 ;
        RECT 10.760000 3.505000 10.930000 3.675000 ;
        RECT 11.760000 3.505000 11.930000 3.675000 ;
        RECT 12.120000 3.505000 12.290000 3.675000 ;
        RECT 12.480000 3.505000 12.650000 3.675000 ;
        RECT 13.320000 3.505000 13.490000 3.675000 ;
        RECT 13.680000 3.505000 13.850000 3.675000 ;
        RECT 14.040000 3.505000 14.210000 3.675000 ;
      LAYER met1 ;
        RECT 0.000000 3.445000 14.880000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.615000  0.380000 1.295000 ;
      RECT  0.115000 1.295000  1.510000 1.465000 ;
      RECT  0.115000 1.465000  0.365000 3.735000 ;
      RECT  1.180000 1.465000  1.510000 1.895000 ;
      RECT  1.340000 0.265000  2.290000 0.435000 ;
      RECT  1.340000 0.435000  1.510000 1.295000 ;
      RECT  1.675000 2.945000  2.005000 3.735000 ;
      RECT  1.690000 0.615000  1.940000 2.275000 ;
      RECT  1.690000 2.275000  2.835000 2.445000 ;
      RECT  1.690000 2.445000  2.005000 2.945000 ;
      RECT  2.120000 0.435000  2.290000 1.175000 ;
      RECT  2.120000 1.175000  3.185000 1.345000 ;
      RECT  2.665000 2.445000  2.835000 3.755000 ;
      RECT  3.015000 1.345000  3.185000 3.285000 ;
      RECT  3.015000 3.285000  5.005000 3.615000 ;
      RECT  3.185000 0.495000  3.535000 0.995000 ;
      RECT  3.365000 0.995000  3.535000 3.105000 ;
      RECT  3.715000 1.085000  3.885000 3.285000 ;
      RECT  4.065000 0.495000  4.315000 0.965000 ;
      RECT  4.065000 0.965000  6.315000 1.135000 ;
      RECT  4.065000 1.135000  4.235000 2.605000 ;
      RECT  4.065000 2.605000  4.395000 3.105000 ;
      RECT  4.415000 1.495000  4.655000 1.805000 ;
      RECT  4.415000 1.805000  6.985000 1.975000 ;
      RECT  4.415000 1.975000  4.655000 2.165000 ;
      RECT  4.835000 2.155000  6.635000 2.325000 ;
      RECT  4.835000 2.325000  5.005000 3.285000 ;
      RECT  5.135000 1.315000  5.865000 1.625000 ;
      RECT  5.185000 2.505000  6.285000 2.675000 ;
      RECT  5.185000 2.675000  5.425000 3.555000 ;
      RECT  5.985000 0.265000  6.315000 0.965000 ;
      RECT  6.115000 2.675000  6.895000 2.845000 ;
      RECT  6.465000 2.325000  8.960000 2.495000 ;
      RECT  6.565000 2.845000  6.895000 3.105000 ;
      RECT  6.815000 1.975000  8.450000 2.145000 ;
      RECT  8.280000 1.545000  8.785000 1.705000 ;
      RECT  8.280000 1.705000  9.310000 1.875000 ;
      RECT  8.280000 1.875000  8.450000 1.975000 ;
      RECT  8.630000 2.085000  8.960000 2.325000 ;
      RECT  8.695000 2.675000  9.310000 2.845000 ;
      RECT  8.695000 2.845000  8.865000 3.595000 ;
      RECT  8.695000 3.595000  9.825000 3.805000 ;
      RECT  9.025000 1.190000  9.660000 1.475000 ;
      RECT  9.045000 3.025000  9.660000 3.415000 ;
      RECT  9.140000 1.875000  9.310000 2.675000 ;
      RECT  9.490000 1.475000  9.660000 2.315000 ;
      RECT  9.490000 2.315000 12.210000 2.485000 ;
      RECT  9.490000 2.485000  9.660000 3.025000 ;
      RECT 10.305000 1.545000 10.635000 1.655000 ;
      RECT 10.305000 1.655000 12.560000 1.825000 ;
      RECT 10.305000 1.825000 10.635000 2.135000 ;
      RECT 11.300000 3.255000 11.550000 3.755000 ;
      RECT 11.380000 3.005000 12.560000 3.175000 ;
      RECT 11.380000 3.175000 11.550000 3.255000 ;
      RECT 11.410000 2.485000 12.210000 2.675000 ;
      RECT 11.410000 2.675000 11.740000 2.825000 ;
      RECT 11.880000 2.005000 12.210000 2.315000 ;
      RECT 12.120000 0.975000 12.450000 1.655000 ;
      RECT 12.390000 1.825000 12.560000 3.005000 ;
      RECT 12.745000 0.975000 13.075000 1.475000 ;
      RECT 12.865000 1.475000 13.075000 2.225000 ;
      RECT 12.865000 2.225000 14.240000 2.395000 ;
      RECT 12.865000 2.395000 13.115000 3.365000 ;
      RECT 13.910000 1.725000 14.240000 2.225000 ;
  END
END sky130_fd_sc_hvl__dfstp_1
