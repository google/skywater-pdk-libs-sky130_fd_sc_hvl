* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_4 A VGND VNB VPB VPWR X
M1000 VGND a_149_81# X VNB nhv w=750000u l=500000u
+  ad=6.3375e+11p pd=6.19e+06u as=4.2e+11p ps=4.12e+06u
M1001 a_149_81# A VPWR VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=1.2675e+12p ps=1.069e+07u
M1002 VGND a_149_81# X VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_149_81# VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_149_81# X VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=8.4e+11p ps=7.12e+06u
M1005 X a_149_81# VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_149_81# X VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_149_81# A VGND VNB nhv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
M1008 X a_149_81# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_149_81# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
