# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__lsbufhv2lv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbufhv2lv_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  8.140000 ;
  SYMMETRY X Y R90 ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.630000 4.870000 1.300000 5.200000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.492900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 0.735000 3.960000 3.245000 ;
    END
  END X
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 8.090000 3.305000 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 8.160000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 8.160000 8.255000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 8.160000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 8.160000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.985000 0.885000 4.155000 ;
      RECT 0.000000  8.055000 8.160000 8.225000 ;
      RECT 0.130000  2.260000 0.460000 3.445000 ;
      RECT 0.130000  3.445000 0.720000 3.675000 ;
      RECT 0.130000  4.465000 0.720000 4.695000 ;
      RECT 0.130000  4.695000 0.460000 5.880000 ;
      RECT 0.170000  1.080000 0.420000 1.565000 ;
      RECT 0.170000  1.565000 1.750000 1.895000 ;
      RECT 0.170000  6.220000 1.750000 6.575000 ;
      RECT 0.170000  6.575000 0.420000 7.060000 ;
      RECT 0.630000  2.835000 1.750000 3.085000 ;
      RECT 0.895000  0.395000 1.485000 1.395000 ;
      RECT 0.895000  6.745000 1.485000 7.745000 ;
      RECT 0.950000  1.895000 1.200000 2.590000 ;
      RECT 0.950000  5.550000 1.750000 6.220000 ;
      RECT 1.445000  1.895000 1.750000 2.235000 ;
      RECT 1.470000  3.085000 1.750000 5.550000 ;
      RECT 1.920000  0.685000 2.250000 4.255000 ;
      RECT 1.920000  4.255000 3.960000 4.595000 ;
      RECT 1.920000  5.195000 3.540000 5.445000 ;
      RECT 1.920000  5.445000 2.250000 7.455000 ;
      RECT 2.530000  5.615000 3.120000 7.745000 ;
      RECT 2.570000  0.395000 3.160000 3.910000 ;
      RECT 3.290000  5.445000 3.540000 5.595000 ;
      RECT 3.290000  5.595000 5.170000 5.845000 ;
      RECT 3.480000  5.845000 3.810000 7.455000 ;
      RECT 3.710000  4.595000 3.960000 5.415000 ;
      RECT 3.780000  3.415000 4.750000 4.085000 ;
      RECT 4.130000  0.395000 4.720000 1.515000 ;
      RECT 4.130000  2.085000 4.400000 3.075000 ;
      RECT 4.130000  3.075000 4.750000 3.415000 ;
      RECT 4.130000  4.085000 4.400000 5.415000 ;
      RECT 4.570000  2.085000 4.820000 2.655000 ;
      RECT 4.570000  2.655000 5.170000 2.905000 ;
      RECT 4.920000  2.905000 5.170000 5.595000 ;
      RECT 7.275000  3.985000 8.160000 4.155000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.155000  8.055000 0.325000 8.225000 ;
      RECT 0.160000  3.475000 0.330000 3.645000 ;
      RECT 0.160000  4.495000 0.330000 4.665000 ;
      RECT 0.520000  3.475000 0.690000 3.645000 ;
      RECT 0.520000  4.495000 0.690000 4.665000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.635000  8.055000 0.805000 8.225000 ;
      RECT 0.925000  0.425000 1.095000 0.595000 ;
      RECT 0.925000  7.545000 1.095000 7.715000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  8.055000 1.285000 8.225000 ;
      RECT 1.285000  0.425000 1.455000 0.595000 ;
      RECT 1.285000  7.545000 1.455000 7.715000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  8.055000 1.765000 8.225000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  8.055000 2.245000 8.225000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  8.055000 2.725000 8.225000 ;
      RECT 2.560000  7.545000 2.730000 7.715000 ;
      RECT 2.600000  0.425000 2.770000 0.595000 ;
      RECT 2.920000  7.545000 3.090000 7.715000 ;
      RECT 2.960000  0.425000 3.130000 0.595000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  8.055000 3.205000 8.225000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  8.055000 3.685000 8.225000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  8.055000 4.165000 8.225000 ;
      RECT 4.160000  0.425000 4.330000 0.595000 ;
      RECT 4.160000  3.105000 4.330000 3.275000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  8.055000 4.645000 8.225000 ;
      RECT 4.520000  0.425000 4.690000 0.595000 ;
      RECT 4.520000  3.105000 4.690000 3.275000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  8.055000 5.125000 8.225000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  8.055000 5.605000 8.225000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  8.055000 6.085000 8.225000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  8.055000 6.565000 8.225000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  8.055000 7.045000 8.225000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.355000  8.055000 7.525000 8.225000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 7.835000  8.055000 8.005000 8.225000 ;
    LAYER met1 ;
      RECT 0.000000 -0.115000 8.160000 0.115000 ;
      RECT 0.000000  0.255000 8.160000 0.625000 ;
      RECT 0.000000  3.445000 8.160000 3.815000 ;
  END
END sky130_fd_sc_hvl__lsbufhv2lv_1
END LIBRARY
