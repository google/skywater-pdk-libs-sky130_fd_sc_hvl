* File: sky130_fd_sc_hvl__inv_8.pxi.spice
* Created: Wed Sep  2 09:07:07 2020
* 
x_PM_SKY130_FD_SC_HVL__INV_8%VNB N_VNB_M1000_b VNB N_VNB_c_14_p VNB
+ PM_SKY130_FD_SC_HVL__INV_8%VNB
x_PM_SKY130_FD_SC_HVL__INV_8%VPB N_VPB_M1003_b VPB N_VPB_c_30_p VPB
+ PM_SKY130_FD_SC_HVL__INV_8%VPB
x_PM_SKY130_FD_SC_HVL__INV_8%A N_A_c_86_n N_A_M1000_g N_A_M1003_g N_A_c_87_n
+ N_A_M1001_g N_A_M1004_g N_A_c_88_n N_A_M1002_g N_A_M1007_g N_A_c_89_n
+ N_A_M1005_g N_A_M1009_g N_A_c_90_n N_A_M1006_g N_A_M1011_g N_A_c_91_n
+ N_A_M1008_g N_A_M1012_g N_A_c_92_n N_A_M1010_g N_A_M1014_g N_A_c_93_n
+ N_A_M1013_g N_A_M1015_g A A A A A A A N_A_c_94_n N_A_c_95_n
+ PM_SKY130_FD_SC_HVL__INV_8%A
x_PM_SKY130_FD_SC_HVL__INV_8%VPWR N_VPWR_M1003_s N_VPWR_M1004_s N_VPWR_M1009_s
+ N_VPWR_M1012_s N_VPWR_M1015_s N_VPWR_c_264_n N_VPWR_c_267_n N_VPWR_c_270_n
+ N_VPWR_c_273_n N_VPWR_c_276_n N_VPWR_c_279_n N_VPWR_c_282_n N_VPWR_c_285_n
+ VPWR N_VPWR_c_288_n N_VPWR_c_311_n N_VPWR_c_316_n N_VPWR_c_321_n
+ N_VPWR_c_326_n N_VPWR_c_289_n PM_SKY130_FD_SC_HVL__INV_8%VPWR
x_PM_SKY130_FD_SC_HVL__INV_8%Y N_Y_M1000_d N_Y_M1002_d N_Y_M1006_d N_Y_M1010_d
+ N_Y_M1003_d N_Y_M1007_d N_Y_M1011_d N_Y_M1014_d N_Y_c_466_p N_Y_c_367_n
+ N_Y_c_369_n N_Y_c_373_n N_Y_c_362_n N_Y_c_379_n N_Y_c_468_p N_Y_c_383_n
+ N_Y_c_385_n N_Y_c_363_n N_Y_c_470_p N_Y_c_393_n N_Y_c_395_n N_Y_c_364_n
+ N_Y_c_403_n N_Y_c_365_n N_Y_c_360_n N_Y_c_361_n N_Y_c_413_n N_Y_c_415_n
+ N_Y_c_419_n N_Y_c_421_n N_Y_c_425_n Y N_Y_c_429_n PM_SKY130_FD_SC_HVL__INV_8%Y
x_PM_SKY130_FD_SC_HVL__INV_8%VGND N_VGND_M1000_s N_VGND_M1001_s N_VGND_M1005_s
+ N_VGND_M1008_s N_VGND_M1013_s N_VGND_c_481_n N_VGND_c_483_n VGND
+ N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_487_n N_VGND_c_489_n N_VGND_c_490_n
+ N_VGND_c_491_n N_VGND_c_492_n N_VGND_c_493_n N_VGND_c_494_n
+ PM_SKY130_FD_SC_HVL__INV_8%VGND
cc_1 N_VNB_M1000_b N_A_c_86_n 0.0426879f $X=-0.33 $Y=-0.265 $X2=0.91 $Y2=1.565
cc_2 N_VNB_M1000_b N_A_c_87_n 0.0365315f $X=-0.33 $Y=-0.265 $X2=1.69 $Y2=1.565
cc_3 N_VNB_M1000_b N_A_c_88_n 0.0371653f $X=-0.33 $Y=-0.265 $X2=2.47 $Y2=1.565
cc_4 N_VNB_M1000_b N_A_c_89_n 0.0371653f $X=-0.33 $Y=-0.265 $X2=3.25 $Y2=1.565
cc_5 N_VNB_M1000_b N_A_c_90_n 0.0371653f $X=-0.33 $Y=-0.265 $X2=4.03 $Y2=1.565
cc_6 N_VNB_M1000_b N_A_c_91_n 0.0383712f $X=-0.33 $Y=-0.265 $X2=4.81 $Y2=1.565
cc_7 N_VNB_M1000_b N_A_c_92_n 0.0379462f $X=-0.33 $Y=-0.265 $X2=5.73 $Y2=1.565
cc_8 N_VNB_M1000_b N_A_c_93_n 0.0406388f $X=-0.33 $Y=-0.265 $X2=6.51 $Y2=1.565
cc_9 N_VNB_M1000_b N_A_c_94_n 0.270046f $X=-0.33 $Y=-0.265 $X2=6.595 $Y2=1.73
cc_10 N_VNB_M1000_b N_A_c_95_n 0.0117206f $X=-0.33 $Y=-0.265 $X2=6.595 $Y2=1.73
cc_11 N_VNB_M1000_b N_Y_c_360_n 0.00814524f $X=-0.33 $Y=-0.265 $X2=0.91
+ $Y2=1.815
cc_12 N_VNB_M1000_b N_Y_c_361_n 0.0229642f $X=-0.33 $Y=-0.265 $X2=1.83 $Y2=1.815
cc_13 N_VNB_M1000_b N_VGND_c_481_n 0.0205089f $X=-0.33 $Y=-0.265 $X2=2.61
+ $Y2=2.065
cc_14 N_VNB_c_14_p N_VGND_c_481_n 0.00102686f $X=0.24 $Y=0 $X2=2.61 $Y2=2.065
cc_15 N_VNB_M1000_b N_VGND_c_483_n 0.0195973f $X=-0.33 $Y=-0.265 $X2=2.61
+ $Y2=2.965
cc_16 N_VNB_M1000_b N_VGND_c_484_n 0.0155621f $X=-0.33 $Y=-0.265 $X2=4.17
+ $Y2=2.965
cc_17 N_VNB_M1000_b N_VGND_c_485_n 0.0972358f $X=-0.33 $Y=-0.265 $X2=5.73
+ $Y2=1.565
cc_18 N_VNB_c_14_p N_VGND_c_485_n 0.0024636f $X=0.24 $Y=0 $X2=5.73 $Y2=1.565
cc_19 N_VNB_M1000_b N_VGND_c_487_n 0.242552f $X=-0.33 $Y=-0.265 $X2=6.51
+ $Y2=2.965
cc_20 N_VNB_c_14_p N_VGND_c_487_n 0.0160888f $X=0.24 $Y=0 $X2=6.51 $Y2=2.965
cc_21 N_VNB_M1000_b N_VGND_c_489_n 0.00648994f $X=-0.33 $Y=-0.265 $X2=3.035
+ $Y2=1.58
cc_22 N_VNB_M1000_b N_VGND_c_490_n 0.00820065f $X=-0.33 $Y=-0.265 $X2=4.475
+ $Y2=1.58
cc_23 N_VNB_M1000_b N_VGND_c_491_n 0.00648092f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_24 N_VNB_M1000_b N_VGND_c_492_n 0.00820065f $X=-0.33 $Y=-0.265 $X2=0.475
+ $Y2=1.815
cc_25 N_VNB_M1000_b N_VGND_c_493_n 0.00752522f $X=-0.33 $Y=-0.265 $X2=1.69
+ $Y2=1.815
cc_26 N_VNB_M1000_b N_VGND_c_494_n 0.105347f $X=-0.33 $Y=-0.265 $X2=2.61
+ $Y2=1.815
cc_27 N_VNB_c_14_p N_VGND_c_494_n 0.769619f $X=0.24 $Y=0 $X2=2.61 $Y2=1.815
cc_28 N_VPB_M1003_b N_A_M1003_g 0.0438905f $X=-0.33 $Y=1.885 $X2=1.05 $Y2=2.965
cc_29 VPB N_A_M1003_g 0.00970178f $X=0 $Y=3.955 $X2=1.05 $Y2=2.965
cc_30 N_VPB_c_30_p N_A_M1003_g 0.0135168f $X=6.96 $Y=4.07 $X2=1.05 $Y2=2.965
cc_31 N_VPB_M1003_b N_A_M1004_g 0.035291f $X=-0.33 $Y=1.885 $X2=1.83 $Y2=2.965
cc_32 VPB N_A_M1004_g 0.00970178f $X=0 $Y=3.955 $X2=1.83 $Y2=2.965
cc_33 N_VPB_c_30_p N_A_M1004_g 0.0135156f $X=6.96 $Y=4.07 $X2=1.83 $Y2=2.965
cc_34 N_VPB_M1003_b N_A_M1007_g 0.035291f $X=-0.33 $Y=1.885 $X2=2.61 $Y2=2.965
cc_35 VPB N_A_M1007_g 0.00970178f $X=0 $Y=3.955 $X2=2.61 $Y2=2.965
cc_36 N_VPB_c_30_p N_A_M1007_g 0.0135156f $X=6.96 $Y=4.07 $X2=2.61 $Y2=2.965
cc_37 N_VPB_M1003_b N_A_M1009_g 0.035291f $X=-0.33 $Y=1.885 $X2=3.39 $Y2=2.965
cc_38 VPB N_A_M1009_g 0.00970178f $X=0 $Y=3.955 $X2=3.39 $Y2=2.965
cc_39 N_VPB_c_30_p N_A_M1009_g 0.0135156f $X=6.96 $Y=4.07 $X2=3.39 $Y2=2.965
cc_40 N_VPB_M1003_b N_A_M1011_g 0.035291f $X=-0.33 $Y=1.885 $X2=4.17 $Y2=2.965
cc_41 VPB N_A_M1011_g 0.00970178f $X=0 $Y=3.955 $X2=4.17 $Y2=2.965
cc_42 N_VPB_c_30_p N_A_M1011_g 0.0135156f $X=6.96 $Y=4.07 $X2=4.17 $Y2=2.965
cc_43 N_VPB_M1003_b N_A_M1012_g 0.035291f $X=-0.33 $Y=1.885 $X2=4.95 $Y2=2.965
cc_44 VPB N_A_M1012_g 0.00970178f $X=0 $Y=3.955 $X2=4.95 $Y2=2.965
cc_45 N_VPB_c_30_p N_A_M1012_g 0.0135156f $X=6.96 $Y=4.07 $X2=4.95 $Y2=2.965
cc_46 N_VPB_M1003_b N_A_M1014_g 0.035291f $X=-0.33 $Y=1.885 $X2=5.73 $Y2=2.965
cc_47 VPB N_A_M1014_g 0.00970178f $X=0 $Y=3.955 $X2=5.73 $Y2=2.965
cc_48 N_VPB_c_30_p N_A_M1014_g 0.0135156f $X=6.96 $Y=4.07 $X2=5.73 $Y2=2.965
cc_49 N_VPB_M1003_b N_A_M1015_g 0.0404836f $X=-0.33 $Y=1.885 $X2=6.51 $Y2=2.965
cc_50 VPB N_A_M1015_g 0.00970178f $X=0 $Y=3.955 $X2=6.51 $Y2=2.965
cc_51 N_VPB_c_30_p N_A_M1015_g 0.0135156f $X=6.96 $Y=4.07 $X2=6.51 $Y2=2.965
cc_52 N_VPB_M1003_b N_A_c_94_n 0.172395f $X=-0.33 $Y=1.885 $X2=6.595 $Y2=1.73
cc_53 N_VPB_M1003_b N_VPWR_c_264_n 0.0010569f $X=-0.33 $Y=1.885 $X2=2.47
+ $Y2=1.08
cc_54 VPB N_VPWR_c_264_n 0.00314862f $X=0 $Y=3.955 $X2=2.47 $Y2=1.08
cc_55 N_VPB_c_30_p N_VPWR_c_264_n 0.0476561f $X=6.96 $Y=4.07 $X2=2.47 $Y2=1.08
cc_56 N_VPB_M1003_b N_VPWR_c_267_n 0.00788f $X=-0.33 $Y=1.885 $X2=2.47 $Y2=1.08
cc_57 VPB N_VPWR_c_267_n 0.00319302f $X=0 $Y=3.955 $X2=2.47 $Y2=1.08
cc_58 N_VPB_c_30_p N_VPWR_c_267_n 0.0562134f $X=6.96 $Y=4.07 $X2=2.47 $Y2=1.08
cc_59 N_VPB_M1003_b N_VPWR_c_270_n 0.0010569f $X=-0.33 $Y=1.885 $X2=2.61
+ $Y2=2.065
cc_60 VPB N_VPWR_c_270_n 0.00262607f $X=0 $Y=3.955 $X2=2.61 $Y2=2.065
cc_61 N_VPB_c_30_p N_VPWR_c_270_n 0.0405322f $X=6.96 $Y=4.07 $X2=2.61 $Y2=2.065
cc_62 N_VPB_M1003_b N_VPWR_c_273_n 0.0010569f $X=-0.33 $Y=1.885 $X2=2.61
+ $Y2=2.965
cc_63 VPB N_VPWR_c_273_n 0.00262607f $X=0 $Y=3.955 $X2=2.61 $Y2=2.965
cc_64 N_VPB_c_30_p N_VPWR_c_273_n 0.0405322f $X=6.96 $Y=4.07 $X2=2.61 $Y2=2.965
cc_65 N_VPB_M1003_b N_VPWR_c_276_n 0.00450725f $X=-0.33 $Y=1.885 $X2=3.25
+ $Y2=1.565
cc_66 VPB N_VPWR_c_276_n 0.00496432f $X=0 $Y=3.955 $X2=3.25 $Y2=1.565
cc_67 N_VPB_c_30_p N_VPWR_c_276_n 0.0758096f $X=6.96 $Y=4.07 $X2=3.25 $Y2=1.565
cc_68 N_VPB_M1003_b N_VPWR_c_279_n 0.00105831f $X=-0.33 $Y=1.885 $X2=3.39
+ $Y2=2.965
cc_69 VPB N_VPWR_c_279_n 0.00385318f $X=0 $Y=3.955 $X2=3.39 $Y2=2.965
cc_70 N_VPB_c_30_p N_VPWR_c_279_n 0.0545489f $X=6.96 $Y=4.07 $X2=3.39 $Y2=2.965
cc_71 N_VPB_M1003_b N_VPWR_c_282_n 0.00105831f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_282_n 0.00385318f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_73 N_VPB_c_30_p N_VPWR_c_282_n 0.0545489f $X=6.96 $Y=4.07 $X2=0 $Y2=0
cc_74 N_VPB_M1003_b N_VPWR_c_285_n 0.00105831f $X=-0.33 $Y=1.885 $X2=4.03
+ $Y2=1.08
cc_75 VPB N_VPWR_c_285_n 0.00385318f $X=0 $Y=3.955 $X2=4.03 $Y2=1.08
cc_76 N_VPB_c_30_p N_VPWR_c_285_n 0.0545489f $X=6.96 $Y=4.07 $X2=4.03 $Y2=1.08
cc_77 N_VPB_M1003_b N_VPWR_c_288_n 0.0734495f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_78 N_VPB_M1003_b N_VPWR_c_289_n 0.0523846f $X=-0.33 $Y=1.885 $X2=5.73
+ $Y2=1.815
cc_79 VPB N_VPWR_c_289_n 0.76217f $X=0 $Y=3.955 $X2=5.73 $Y2=1.815
cc_80 N_VPB_c_30_p N_VPWR_c_289_n 0.024597f $X=6.96 $Y=4.07 $X2=5.73 $Y2=1.815
cc_81 N_VPB_M1003_b N_Y_c_362_n 0.00261732f $X=-0.33 $Y=1.885 $X2=4.81 $Y2=1.08
cc_82 N_VPB_M1003_b N_Y_c_363_n 0.00261732f $X=-0.33 $Y=1.885 $X2=6.51 $Y2=1.08
cc_83 N_VPB_M1003_b N_Y_c_364_n 0.00261732f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_84 N_VPB_M1003_b N_Y_c_365_n 0.0165641f $X=-0.33 $Y=1.885 $X2=0.475 $Y2=1.73
cc_85 N_VPB_M1003_b N_Y_c_361_n 0.00748448f $X=-0.33 $Y=1.885 $X2=1.83 $Y2=1.815
cc_86 N_A_M1003_g N_VPWR_c_264_n 0.0149041f $X=1.05 $Y=2.965 $X2=6.96 $Y2=0
cc_87 N_A_M1004_g N_VPWR_c_264_n 0.00984257f $X=1.83 $Y=2.965 $X2=6.96 $Y2=0
cc_88 N_A_M1003_g N_VPWR_c_267_n 0.00528717f $X=1.05 $Y=2.965 $X2=6.96 $Y2=0
cc_89 N_A_M1007_g N_VPWR_c_270_n 0.00984257f $X=2.61 $Y=2.965 $X2=0 $Y2=0
cc_90 N_A_M1009_g N_VPWR_c_270_n 0.00984257f $X=3.39 $Y=2.965 $X2=0 $Y2=0
cc_91 N_A_M1011_g N_VPWR_c_273_n 0.00984257f $X=4.17 $Y=2.965 $X2=0 $Y2=0
cc_92 N_A_M1012_g N_VPWR_c_273_n 0.00984257f $X=4.95 $Y=2.965 $X2=0 $Y2=0
cc_93 N_A_M1014_g N_VPWR_c_276_n 0.00984257f $X=5.73 $Y=2.965 $X2=0 $Y2=0
cc_94 N_A_M1015_g N_VPWR_c_276_n 0.0170097f $X=6.51 $Y=2.965 $X2=0 $Y2=0
cc_95 N_A_M1004_g N_VPWR_c_279_n 0.00656544f $X=1.83 $Y=2.965 $X2=0 $Y2=0
cc_96 N_A_M1007_g N_VPWR_c_279_n 0.00656544f $X=2.61 $Y=2.965 $X2=0 $Y2=0
cc_97 N_A_M1009_g N_VPWR_c_282_n 0.00656544f $X=3.39 $Y=2.965 $X2=0 $Y2=0
cc_98 N_A_M1011_g N_VPWR_c_282_n 0.00656544f $X=4.17 $Y=2.965 $X2=0 $Y2=0
cc_99 N_A_M1012_g N_VPWR_c_285_n 0.00656544f $X=4.95 $Y=2.965 $X2=0 $Y2=0
cc_100 N_A_M1014_g N_VPWR_c_285_n 0.00656544f $X=5.73 $Y=2.965 $X2=0 $Y2=0
cc_101 N_A_M1003_g N_VPWR_c_288_n 0.0482271f $X=1.05 $Y=2.965 $X2=0 $Y2=0
cc_102 N_A_M1004_g N_VPWR_c_288_n 9.35642e-19 $X=1.83 $Y=2.965 $X2=0 $Y2=0
cc_103 N_A_c_94_n N_VPWR_c_288_n 0.0117776f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_104 N_A_c_95_n N_VPWR_c_288_n 0.0183431f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_105 N_A_M1003_g N_VPWR_c_311_n 0.0011619f $X=1.05 $Y=2.965 $X2=0 $Y2=0
cc_106 N_A_M1004_g N_VPWR_c_311_n 0.0581477f $X=1.83 $Y=2.965 $X2=0 $Y2=0
cc_107 N_A_M1007_g N_VPWR_c_311_n 0.0570434f $X=2.61 $Y=2.965 $X2=0 $Y2=0
cc_108 N_A_M1009_g N_VPWR_c_311_n 4.54877e-19 $X=3.39 $Y=2.965 $X2=0 $Y2=0
cc_109 N_A_c_94_n N_VPWR_c_311_n 5.59492e-19 $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_110 N_A_M1007_g N_VPWR_c_316_n 4.54877e-19 $X=2.61 $Y=2.965 $X2=0 $Y2=0
cc_111 N_A_M1009_g N_VPWR_c_316_n 0.0570434f $X=3.39 $Y=2.965 $X2=0 $Y2=0
cc_112 N_A_M1011_g N_VPWR_c_316_n 0.0570434f $X=4.17 $Y=2.965 $X2=0 $Y2=0
cc_113 N_A_M1012_g N_VPWR_c_316_n 4.54877e-19 $X=4.95 $Y=2.965 $X2=0 $Y2=0
cc_114 N_A_c_94_n N_VPWR_c_316_n 5.59492e-19 $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_115 N_A_M1011_g N_VPWR_c_321_n 4.54877e-19 $X=4.17 $Y=2.965 $X2=0 $Y2=0
cc_116 N_A_M1012_g N_VPWR_c_321_n 0.0570434f $X=4.95 $Y=2.965 $X2=0 $Y2=0
cc_117 N_A_M1014_g N_VPWR_c_321_n 0.0570434f $X=5.73 $Y=2.965 $X2=0 $Y2=0
cc_118 N_A_M1015_g N_VPWR_c_321_n 4.54877e-19 $X=6.51 $Y=2.965 $X2=0 $Y2=0
cc_119 N_A_c_94_n N_VPWR_c_321_n 5.62414e-19 $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_120 N_A_M1014_g N_VPWR_c_326_n 4.47096e-19 $X=5.73 $Y=2.965 $X2=0 $Y2=0
cc_121 N_A_M1015_g N_VPWR_c_326_n 0.0569302f $X=6.51 $Y=2.965 $X2=0 $Y2=0
cc_122 N_A_M1003_g N_VPWR_c_289_n 0.0159798f $X=1.05 $Y=2.965 $X2=0 $Y2=0
cc_123 N_A_M1004_g N_VPWR_c_289_n 0.00994001f $X=1.83 $Y=2.965 $X2=0 $Y2=0
cc_124 N_A_M1007_g N_VPWR_c_289_n 0.00994001f $X=2.61 $Y=2.965 $X2=0 $Y2=0
cc_125 N_A_M1009_g N_VPWR_c_289_n 0.00994001f $X=3.39 $Y=2.965 $X2=0 $Y2=0
cc_126 N_A_M1011_g N_VPWR_c_289_n 0.00994001f $X=4.17 $Y=2.965 $X2=0 $Y2=0
cc_127 N_A_M1012_g N_VPWR_c_289_n 0.00994001f $X=4.95 $Y=2.965 $X2=0 $Y2=0
cc_128 N_A_M1014_g N_VPWR_c_289_n 0.00994001f $X=5.73 $Y=2.965 $X2=0 $Y2=0
cc_129 N_A_M1015_g N_VPWR_c_289_n 0.010089f $X=6.51 $Y=2.965 $X2=0 $Y2=0
cc_130 N_A_M1003_g N_Y_c_367_n 0.0324785f $X=1.05 $Y=2.965 $X2=0 $Y2=0
cc_131 N_A_M1004_g N_Y_c_367_n 0.0259143f $X=1.83 $Y=2.965 $X2=0 $Y2=0
cc_132 N_A_c_87_n N_Y_c_369_n 0.0252852f $X=1.69 $Y=1.565 $X2=0 $Y2=0
cc_133 N_A_c_88_n N_Y_c_369_n 0.0252852f $X=2.47 $Y=1.565 $X2=0 $Y2=0
cc_134 N_A_c_94_n N_Y_c_369_n 0.00266332f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_135 N_A_c_95_n N_Y_c_369_n 0.0840169f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_136 N_A_c_94_n N_Y_c_373_n 0.00275161f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_137 N_A_c_95_n N_Y_c_373_n 0.0142996f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_138 N_A_M1004_g N_Y_c_362_n 0.0195999f $X=1.83 $Y=2.965 $X2=0 $Y2=0
cc_139 N_A_M1007_g N_Y_c_362_n 0.0195999f $X=2.61 $Y=2.965 $X2=0 $Y2=0
cc_140 N_A_c_94_n N_Y_c_362_n 0.0243226f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_141 N_A_c_95_n N_Y_c_362_n 0.0695158f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_142 N_A_M1003_g N_Y_c_379_n 0.00874394f $X=1.05 $Y=2.965 $X2=0 $Y2=0
cc_143 N_A_M1004_g N_Y_c_379_n 0.00198744f $X=1.83 $Y=2.965 $X2=0 $Y2=0
cc_144 N_A_c_94_n N_Y_c_379_n 0.0104892f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_145 N_A_c_95_n N_Y_c_379_n 0.0208988f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_146 N_A_M1007_g N_Y_c_383_n 0.0259143f $X=2.61 $Y=2.965 $X2=0 $Y2=0
cc_147 N_A_M1009_g N_Y_c_383_n 0.0259143f $X=3.39 $Y=2.965 $X2=0 $Y2=0
cc_148 N_A_c_89_n N_Y_c_385_n 0.0252852f $X=3.25 $Y=1.565 $X2=0 $Y2=0
cc_149 N_A_c_90_n N_Y_c_385_n 0.0252852f $X=4.03 $Y=1.565 $X2=0 $Y2=0
cc_150 N_A_c_94_n N_Y_c_385_n 0.00266332f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_151 N_A_c_95_n N_Y_c_385_n 0.0840169f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_152 N_A_M1009_g N_Y_c_363_n 0.0195999f $X=3.39 $Y=2.965 $X2=0 $Y2=0
cc_153 N_A_M1011_g N_Y_c_363_n 0.0195999f $X=4.17 $Y=2.965 $X2=0 $Y2=0
cc_154 N_A_c_94_n N_Y_c_363_n 0.0243226f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_155 N_A_c_95_n N_Y_c_363_n 0.0695158f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_156 N_A_M1011_g N_Y_c_393_n 0.0259143f $X=4.17 $Y=2.965 $X2=0 $Y2=0
cc_157 N_A_M1012_g N_Y_c_393_n 0.0259143f $X=4.95 $Y=2.965 $X2=0 $Y2=0
cc_158 N_A_c_91_n N_Y_c_395_n 0.0260043f $X=4.81 $Y=1.565 $X2=0 $Y2=0
cc_159 N_A_c_92_n N_Y_c_395_n 0.0234556f $X=5.73 $Y=1.565 $X2=0 $Y2=0
cc_160 N_A_c_94_n N_Y_c_395_n 0.00619804f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_161 N_A_c_95_n N_Y_c_395_n 0.0881462f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_162 N_A_M1012_g N_Y_c_364_n 0.0195999f $X=4.95 $Y=2.965 $X2=0 $Y2=0
cc_163 N_A_M1014_g N_Y_c_364_n 0.0195999f $X=5.73 $Y=2.965 $X2=0 $Y2=0
cc_164 N_A_c_94_n N_Y_c_364_n 0.0243226f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_165 N_A_c_95_n N_Y_c_364_n 0.0695158f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_166 N_A_M1014_g N_Y_c_403_n 0.0259143f $X=5.73 $Y=2.965 $X2=0 $Y2=0
cc_167 N_A_M1015_g N_Y_c_403_n 0.0259143f $X=6.51 $Y=2.965 $X2=0 $Y2=0
cc_168 N_A_M1015_g N_Y_c_365_n 0.0208295f $X=6.51 $Y=2.965 $X2=0 $Y2=0
cc_169 N_A_c_94_n N_Y_c_365_n 0.00933213f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_170 N_A_c_95_n N_Y_c_365_n 0.0268393f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_171 N_A_c_93_n N_Y_c_360_n 0.0141558f $X=6.51 $Y=1.565 $X2=0 $Y2=0
cc_172 N_A_c_95_n N_Y_c_360_n 0.0126346f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_173 N_A_c_93_n N_Y_c_361_n 0.00727371f $X=6.51 $Y=1.565 $X2=0 $Y2=0
cc_174 N_A_c_94_n N_Y_c_361_n 0.0106582f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_175 N_A_c_95_n N_Y_c_361_n 0.017828f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_176 N_A_c_94_n N_Y_c_413_n 0.00275161f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_177 N_A_c_95_n N_Y_c_413_n 0.0142996f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_178 N_A_M1007_g N_Y_c_415_n 0.00198744f $X=2.61 $Y=2.965 $X2=0 $Y2=0
cc_179 N_A_M1009_g N_Y_c_415_n 0.00198744f $X=3.39 $Y=2.965 $X2=0 $Y2=0
cc_180 N_A_c_94_n N_Y_c_415_n 0.00893179f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_181 N_A_c_95_n N_Y_c_415_n 0.0208988f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_182 N_A_c_94_n N_Y_c_419_n 0.00275161f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_183 N_A_c_95_n N_Y_c_419_n 0.0142996f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_184 N_A_M1011_g N_Y_c_421_n 0.00198744f $X=4.17 $Y=2.965 $X2=0 $Y2=0
cc_185 N_A_M1012_g N_Y_c_421_n 0.00198744f $X=4.95 $Y=2.965 $X2=0 $Y2=0
cc_186 N_A_c_94_n N_Y_c_421_n 0.00893179f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_187 N_A_c_95_n N_Y_c_421_n 0.0208988f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_188 N_A_M1014_g N_Y_c_425_n 0.00198744f $X=5.73 $Y=2.965 $X2=0 $Y2=0
cc_189 N_A_M1015_g N_Y_c_425_n 0.00198744f $X=6.51 $Y=2.965 $X2=0 $Y2=0
cc_190 N_A_c_94_n N_Y_c_425_n 0.00890704f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_191 N_A_c_95_n N_Y_c_425_n 0.0208988f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_192 N_A_c_92_n N_Y_c_429_n 0.0190294f $X=5.73 $Y=1.565 $X2=0 $Y2=0
cc_193 N_A_c_93_n N_Y_c_429_n 0.0391113f $X=6.51 $Y=1.565 $X2=0 $Y2=0
cc_194 N_A_c_94_n N_Y_c_429_n 0.00255747f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_195 N_A_c_95_n N_Y_c_429_n 0.0435735f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_196 N_A_c_93_n N_VGND_c_483_n 0.0156984f $X=6.51 $Y=1.565 $X2=0 $Y2=0
cc_197 N_A_c_92_n N_VGND_c_484_n 0.0081029f $X=5.73 $Y=1.565 $X2=0 $Y2=0
cc_198 N_A_c_93_n N_VGND_c_484_n 0.0122041f $X=6.51 $Y=1.565 $X2=0 $Y2=0
cc_199 N_A_c_86_n N_VGND_c_485_n 0.0485944f $X=0.91 $Y=1.565 $X2=0 $Y2=0
cc_200 N_A_c_87_n N_VGND_c_485_n 6.02822e-19 $X=1.69 $Y=1.565 $X2=0 $Y2=0
cc_201 N_A_c_94_n N_VGND_c_485_n 0.00870161f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_202 N_A_c_95_n N_VGND_c_485_n 0.0458048f $X=6.595 $Y=1.73 $X2=0 $Y2=0
cc_203 N_A_c_86_n N_VGND_c_487_n 0.00676958f $X=0.91 $Y=1.565 $X2=0 $Y2=0
cc_204 N_A_c_87_n N_VGND_c_487_n 0.00520463f $X=1.69 $Y=1.565 $X2=0 $Y2=0
cc_205 N_A_c_86_n N_VGND_c_489_n 5.80624e-19 $X=0.91 $Y=1.565 $X2=0 $Y2=0
cc_206 N_A_c_87_n N_VGND_c_489_n 0.0351936f $X=1.69 $Y=1.565 $X2=0 $Y2=0
cc_207 N_A_c_88_n N_VGND_c_489_n 0.035096f $X=2.47 $Y=1.565 $X2=0 $Y2=0
cc_208 N_A_c_89_n N_VGND_c_489_n 5.69649e-19 $X=3.25 $Y=1.565 $X2=0 $Y2=0
cc_209 N_A_c_88_n N_VGND_c_490_n 0.00328808f $X=2.47 $Y=1.565 $X2=0 $Y2=0
cc_210 N_A_c_89_n N_VGND_c_490_n 0.00328808f $X=3.25 $Y=1.565 $X2=0 $Y2=0
cc_211 N_A_c_88_n N_VGND_c_491_n 5.69649e-19 $X=2.47 $Y=1.565 $X2=0 $Y2=0
cc_212 N_A_c_89_n N_VGND_c_491_n 0.035096f $X=3.25 $Y=1.565 $X2=0 $Y2=0
cc_213 N_A_c_90_n N_VGND_c_491_n 0.035096f $X=4.03 $Y=1.565 $X2=0 $Y2=0
cc_214 N_A_c_91_n N_VGND_c_491_n 5.69649e-19 $X=4.81 $Y=1.565 $X2=0 $Y2=0
cc_215 N_A_c_90_n N_VGND_c_492_n 0.00328808f $X=4.03 $Y=1.565 $X2=0 $Y2=0
cc_216 N_A_c_91_n N_VGND_c_492_n 0.00328808f $X=4.81 $Y=1.565 $X2=0 $Y2=0
cc_217 N_A_c_90_n N_VGND_c_493_n 5.69649e-19 $X=4.03 $Y=1.565 $X2=0 $Y2=0
cc_218 N_A_c_91_n N_VGND_c_493_n 0.0358237f $X=4.81 $Y=1.565 $X2=0 $Y2=0
cc_219 N_A_c_92_n N_VGND_c_493_n 0.0356436f $X=5.73 $Y=1.565 $X2=0 $Y2=0
cc_220 N_A_c_93_n N_VGND_c_493_n 7.59266e-19 $X=6.51 $Y=1.565 $X2=0 $Y2=0
cc_221 N_A_c_86_n N_VGND_c_494_n 0.0104303f $X=0.91 $Y=1.565 $X2=0 $Y2=0
cc_222 N_A_c_87_n N_VGND_c_494_n 0.00420368f $X=1.69 $Y=1.565 $X2=0 $Y2=0
cc_223 N_A_c_88_n N_VGND_c_494_n 0.00420368f $X=2.47 $Y=1.565 $X2=0 $Y2=0
cc_224 N_A_c_89_n N_VGND_c_494_n 0.00420368f $X=3.25 $Y=1.565 $X2=0 $Y2=0
cc_225 N_A_c_90_n N_VGND_c_494_n 0.00420368f $X=4.03 $Y=1.565 $X2=0 $Y2=0
cc_226 N_A_c_91_n N_VGND_c_494_n 0.00420368f $X=4.81 $Y=1.565 $X2=0 $Y2=0
cc_227 N_A_c_92_n N_VGND_c_494_n 0.00663464f $X=5.73 $Y=1.565 $X2=0 $Y2=0
cc_228 N_A_c_93_n N_VGND_c_494_n 0.0118818f $X=6.51 $Y=1.565 $X2=0 $Y2=0
cc_229 N_VPWR_c_264_n N_Y_M1003_d 8.28689e-19 $X=1.775 $Y=3.71 $X2=0 $Y2=0
cc_230 N_VPWR_c_270_n N_Y_M1007_d 8.28689e-19 $X=3.335 $Y=3.71 $X2=0 $Y2=3.955
cc_231 N_VPWR_c_273_n N_Y_M1011_d 8.28689e-19 $X=4.895 $Y=3.71 $X2=0 $Y2=0
cc_232 N_VPWR_c_276_n N_Y_M1014_d 8.28689e-19 $X=6.455 $Y=3.71 $X2=0.24 $Y2=4.07
cc_233 N_VPWR_c_264_n N_Y_c_367_n 0.0178796f $X=1.775 $Y=3.71 $X2=0 $Y2=0
cc_234 N_VPWR_c_288_n N_Y_c_367_n 0.0518399f $X=0.66 $Y=2.55 $X2=0 $Y2=0
cc_235 N_VPWR_c_311_n N_Y_c_367_n 0.0842143f $X=2.22 $Y=2.55 $X2=0 $Y2=0
cc_236 N_VPWR_c_289_n N_Y_c_367_n 0.01238f $X=6.94 $Y=3.56 $X2=0 $Y2=0
cc_237 N_VPWR_c_311_n N_Y_c_362_n 0.0614512f $X=2.22 $Y=2.55 $X2=0 $Y2=0
cc_238 N_VPWR_c_270_n N_Y_c_383_n 0.0178796f $X=3.335 $Y=3.71 $X2=0 $Y2=0
cc_239 N_VPWR_c_311_n N_Y_c_383_n 0.0842143f $X=2.22 $Y=2.55 $X2=0 $Y2=0
cc_240 N_VPWR_c_316_n N_Y_c_383_n 0.0842143f $X=3.78 $Y=2.55 $X2=0 $Y2=0
cc_241 N_VPWR_c_289_n N_Y_c_383_n 0.01238f $X=6.94 $Y=3.56 $X2=0 $Y2=0
cc_242 N_VPWR_c_316_n N_Y_c_363_n 0.0614512f $X=3.78 $Y=2.55 $X2=0 $Y2=0
cc_243 N_VPWR_c_273_n N_Y_c_393_n 0.0178796f $X=4.895 $Y=3.71 $X2=0 $Y2=0
cc_244 N_VPWR_c_316_n N_Y_c_393_n 0.0842143f $X=3.78 $Y=2.55 $X2=0 $Y2=0
cc_245 N_VPWR_c_321_n N_Y_c_393_n 0.0842143f $X=5.34 $Y=2.55 $X2=0 $Y2=0
cc_246 N_VPWR_c_289_n N_Y_c_393_n 0.01238f $X=6.94 $Y=3.56 $X2=0 $Y2=0
cc_247 N_VPWR_c_321_n N_Y_c_364_n 0.0614512f $X=5.34 $Y=2.55 $X2=0 $Y2=0
cc_248 N_VPWR_c_276_n N_Y_c_403_n 0.0178796f $X=6.455 $Y=3.71 $X2=0 $Y2=0
cc_249 N_VPWR_c_321_n N_Y_c_403_n 0.0842143f $X=5.34 $Y=2.55 $X2=0 $Y2=0
cc_250 N_VPWR_c_326_n N_Y_c_403_n 0.0830137f $X=6.9 $Y=2.55 $X2=0 $Y2=0
cc_251 N_VPWR_c_289_n N_Y_c_403_n 0.01238f $X=6.94 $Y=3.56 $X2=0 $Y2=0
cc_252 N_VPWR_c_326_n N_Y_c_365_n 0.0412221f $X=6.9 $Y=2.55 $X2=0 $Y2=0
cc_253 N_Y_c_369_n N_VGND_M1001_s 0.00338216f $X=2.755 $Y=1.315 $X2=0 $Y2=0
cc_254 N_Y_c_385_n N_VGND_M1005_s 0.00338216f $X=4.315 $Y=1.315 $X2=0 $Y2=0
cc_255 N_Y_c_395_n N_VGND_M1008_s 0.00666022f $X=5.915 $Y=1.315 $X2=0 $Y2=0
cc_256 N_Y_c_360_n N_VGND_M1013_s 0.00564286f $X=6.94 $Y=1.31 $X2=-0.33
+ $Y2=-0.265
cc_257 N_Y_c_361_n N_VGND_M1013_s 9.95917e-19 $X=7.025 $Y=2.035 $X2=-0.33
+ $Y2=-0.265
cc_258 N_Y_c_360_n N_VGND_c_483_n 0.0249362f $X=6.94 $Y=1.31 $X2=0 $Y2=0
cc_259 N_Y_c_429_n N_VGND_c_483_n 0.0252638f $X=6.24 $Y=1.31 $X2=0 $Y2=0
cc_260 N_Y_c_360_n N_VGND_c_484_n 0.00216751f $X=6.94 $Y=1.31 $X2=0 $Y2=0
cc_261 N_Y_c_429_n N_VGND_c_484_n 0.0386695f $X=6.24 $Y=1.31 $X2=0 $Y2=0
cc_262 N_Y_c_466_p N_VGND_c_487_n 0.0124682f $X=1.3 $Y=0.895 $X2=0 $Y2=0
cc_263 N_Y_c_369_n N_VGND_c_489_n 0.0623739f $X=2.755 $Y=1.315 $X2=0 $Y2=0
cc_264 N_Y_c_468_p N_VGND_c_490_n 0.0124682f $X=2.86 $Y=0.895 $X2=0 $Y2=0
cc_265 N_Y_c_385_n N_VGND_c_491_n 0.0623739f $X=4.315 $Y=1.315 $X2=0 $Y2=0
cc_266 N_Y_c_470_p N_VGND_c_492_n 0.0124682f $X=4.42 $Y=0.895 $X2=0 $Y2=0
cc_267 N_Y_c_395_n N_VGND_c_493_n 0.0658729f $X=5.915 $Y=1.315 $X2=0 $Y2=0
cc_268 N_Y_c_429_n N_VGND_c_493_n 0.0264894f $X=6.24 $Y=1.31 $X2=0 $Y2=0
cc_269 N_Y_c_466_p N_VGND_c_494_n 0.00694322f $X=1.3 $Y=0.895 $X2=0 $Y2=0
cc_270 N_Y_c_369_n N_VGND_c_494_n 0.0124291f $X=2.755 $Y=1.315 $X2=0 $Y2=0
cc_271 N_Y_c_468_p N_VGND_c_494_n 0.00694322f $X=2.86 $Y=0.895 $X2=0 $Y2=0
cc_272 N_Y_c_385_n N_VGND_c_494_n 0.0124291f $X=4.315 $Y=1.315 $X2=0 $Y2=0
cc_273 N_Y_c_470_p N_VGND_c_494_n 0.00694322f $X=4.42 $Y=0.895 $X2=0 $Y2=0
cc_274 N_Y_c_395_n N_VGND_c_494_n 0.0123792f $X=5.915 $Y=1.315 $X2=0 $Y2=0
cc_275 N_Y_c_360_n N_VGND_c_494_n 0.00460189f $X=6.94 $Y=1.31 $X2=0 $Y2=0
cc_276 N_Y_c_429_n N_VGND_c_494_n 0.020002f $X=6.24 $Y=1.31 $X2=0 $Y2=0
