* File: sky130_fd_sc_hvl__dfrbp_1.pxi.spice
* Created: Wed Sep  2 09:04:58 2020
* 
x_PM_SKY130_FD_SC_HVL__DFRBP_1%VNB N_VNB_M1020_b VNB N_VNB_c_2_p
+ PM_SKY130_FD_SC_HVL__DFRBP_1%VNB
x_PM_SKY130_FD_SC_HVL__DFRBP_1%VPB N_VPB_M1004_b VPB N_VPB_c_117_p
+ PM_SKY130_FD_SC_HVL__DFRBP_1%VPB
x_PM_SKY130_FD_SC_HVL__DFRBP_1%CLK CLK N_CLK_M1020_g N_CLK_M1004_g
+ PM_SKY130_FD_SC_HVL__DFRBP_1%CLK
x_PM_SKY130_FD_SC_HVL__DFRBP_1%A_37_107# N_A_37_107#_M1020_s N_A_37_107#_M1004_s
+ N_A_37_107#_M1003_g N_A_37_107#_M1026_g N_A_37_107#_M1006_g
+ N_A_37_107#_c_290_n N_A_37_107#_c_304_n N_A_37_107#_c_305_n
+ N_A_37_107#_c_291_n N_A_37_107#_c_293_n N_A_37_107#_c_307_n
+ N_A_37_107#_c_310_n N_A_37_107#_c_353_n N_A_37_107#_c_294_n
+ N_A_37_107#_c_312_n N_A_37_107#_c_313_n N_A_37_107#_c_316_n
+ N_A_37_107#_c_319_n N_A_37_107#_c_320_n N_A_37_107#_c_359_p
+ N_A_37_107#_c_360_p N_A_37_107#_c_321_n N_A_37_107#_c_324_n
+ N_A_37_107#_c_430_p N_A_37_107#_c_327_n N_A_37_107#_c_381_p
+ N_A_37_107#_c_330_n N_A_37_107#_c_331_n N_A_37_107#_c_332_n
+ N_A_37_107#_c_335_n N_A_37_107#_c_338_n N_A_37_107#_c_339_n
+ N_A_37_107#_c_340_n N_A_37_107#_c_295_n N_A_37_107#_c_296_n
+ N_A_37_107#_c_297_n N_A_37_107#_c_383_p N_A_37_107#_c_298_n
+ N_A_37_107#_c_343_n N_A_37_107#_c_395_p N_A_37_107#_c_469_p
+ N_A_37_107#_c_384_p N_A_37_107#_M1019_g N_A_37_107#_M1002_g
+ N_A_37_107#_M1005_g PM_SKY130_FD_SC_HVL__DFRBP_1%A_37_107#
x_PM_SKY130_FD_SC_HVL__DFRBP_1%RESET_B N_RESET_B_M1018_g N_RESET_B_c_552_n
+ N_RESET_B_M1013_g N_RESET_B_c_575_n N_RESET_B_M1011_g N_RESET_B_M1025_g
+ N_RESET_B_M1000_g N_RESET_B_c_579_n N_RESET_B_c_554_n N_RESET_B_c_555_n
+ N_RESET_B_c_557_n N_RESET_B_c_559_n N_RESET_B_c_560_n N_RESET_B_c_618_p
+ N_RESET_B_c_561_n N_RESET_B_c_611_p N_RESET_B_c_620_p N_RESET_B_c_562_n
+ N_RESET_B_c_564_n N_RESET_B_c_598_n N_RESET_B_c_566_n N_RESET_B_c_681_p
+ N_RESET_B_c_647_p N_RESET_B_c_567_n N_RESET_B_c_568_n RESET_B
+ N_RESET_B_M1029_g N_RESET_B_c_570_n N_RESET_B_c_571_n
+ PM_SKY130_FD_SC_HVL__DFRBP_1%RESET_B
x_PM_SKY130_FD_SC_HVL__DFRBP_1%D N_D_M1008_g N_D_c_751_n N_D_c_752_n N_D_c_746_n
+ D D N_D_M1014_g PM_SKY130_FD_SC_HVL__DFRBP_1%D
x_PM_SKY130_FD_SC_HVL__DFRBP_1%A_350_107# N_A_350_107#_M1003_d
+ N_A_350_107#_M1026_d N_A_350_107#_M1030_g N_A_350_107#_c_796_n
+ N_A_350_107#_M1016_g N_A_350_107#_c_797_n N_A_350_107#_c_798_n
+ N_A_350_107#_M1015_g N_A_350_107#_c_799_n N_A_350_107#_c_815_n
+ N_A_350_107#_c_816_n N_A_350_107#_c_800_n N_A_350_107#_c_843_n
+ N_A_350_107#_c_844_n N_A_350_107#_c_802_n N_A_350_107#_c_803_n
+ N_A_350_107#_c_804_n N_A_350_107#_c_805_n N_A_350_107#_c_851_n
+ N_A_350_107#_c_806_n N_A_350_107#_c_807_n N_A_350_107#_c_808_n
+ N_A_350_107#_M1028_g N_A_350_107#_c_810_n N_A_350_107#_c_811_n
+ N_A_350_107#_c_819_n N_A_350_107#_c_812_n
+ PM_SKY130_FD_SC_HVL__DFRBP_1%A_350_107#
x_PM_SKY130_FD_SC_HVL__DFRBP_1%A_1176_466# N_A_1176_466#_M1032_d
+ N_A_1176_466#_M1009_d N_A_1176_466#_c_987_n N_A_1176_466#_M1022_g
+ N_A_1176_466#_M1031_g N_A_1176_466#_c_984_n N_A_1176_466#_c_1018_n
+ N_A_1176_466#_c_985_n N_A_1176_466#_c_991_n N_A_1176_466#_c_1049_p
+ N_A_1176_466#_c_986_n N_A_1176_466#_c_1006_n
+ PM_SKY130_FD_SC_HVL__DFRBP_1%A_1176_466#
x_PM_SKY130_FD_SC_HVL__DFRBP_1%A_978_608# N_A_978_608#_M1006_d
+ N_A_978_608#_M1030_d N_A_978_608#_M1011_d N_A_978_608#_c_1073_n
+ N_A_978_608#_M1032_g N_A_978_608#_M1009_g N_A_978_608#_c_1084_n
+ N_A_978_608#_c_1085_n N_A_978_608#_c_1075_n N_A_978_608#_c_1076_n
+ N_A_978_608#_c_1077_n N_A_978_608#_c_1102_n N_A_978_608#_c_1078_n
+ N_A_978_608#_c_1087_n N_A_978_608#_c_1104_n N_A_978_608#_c_1088_n
+ N_A_978_608#_c_1089_n N_A_978_608#_c_1090_n N_A_978_608#_c_1079_n
+ N_A_978_608#_c_1080_n N_A_978_608#_c_1091_n N_A_978_608#_c_1081_n
+ PM_SKY130_FD_SC_HVL__DFRBP_1%A_978_608#
x_PM_SKY130_FD_SC_HVL__DFRBP_1%A_2122_348# N_A_2122_348#_M1001_d
+ N_A_2122_348#_M1025_d N_A_2122_348#_M1027_g N_A_2122_348#_c_1217_n
+ N_A_2122_348#_c_1218_n N_A_2122_348#_c_1256_p N_A_2122_348#_c_1219_n
+ N_A_2122_348#_c_1226_n N_A_2122_348#_c_1235_n N_A_2122_348#_c_1227_n
+ N_A_2122_348#_c_1220_n N_A_2122_348#_c_1222_n N_A_2122_348#_M1007_g
+ PM_SKY130_FD_SC_HVL__DFRBP_1%A_2122_348#
x_PM_SKY130_FD_SC_HVL__DFRBP_1%A_1900_107# N_A_1900_107#_M1016_d
+ N_A_1900_107#_M1002_d N_A_1900_107#_M1001_g N_A_1900_107#_c_1305_n
+ N_A_1900_107#_M1012_g N_A_1900_107#_c_1295_n N_A_1900_107#_M1023_g
+ N_A_1900_107#_M1017_g N_A_1900_107#_c_1298_n N_A_1900_107#_M1033_g
+ N_A_1900_107#_M1024_g N_A_1900_107#_c_1300_n N_A_1900_107#_c_1301_n
+ N_A_1900_107#_c_1314_n N_A_1900_107#_c_1315_n N_A_1900_107#_c_1317_n
+ N_A_1900_107#_c_1326_n N_A_1900_107#_c_1302_n N_A_1900_107#_c_1319_n
+ N_A_1900_107#_c_1320_n N_A_1900_107#_c_1303_n N_A_1900_107#_c_1345_n
+ N_A_1900_107#_c_1304_n PM_SKY130_FD_SC_HVL__DFRBP_1%A_1900_107#
x_PM_SKY130_FD_SC_HVL__DFRBP_1%A_2937_443# N_A_2937_443#_M1024_s
+ N_A_2937_443#_M1033_s N_A_2937_443#_M1010_g N_A_2937_443#_M1021_g
+ N_A_2937_443#_c_1446_n N_A_2937_443#_c_1453_n N_A_2937_443#_c_1447_n
+ N_A_2937_443#_c_1448_n N_A_2937_443#_c_1449_n
+ PM_SKY130_FD_SC_HVL__DFRBP_1%A_2937_443#
x_PM_SKY130_FD_SC_HVL__DFRBP_1%VPWR N_VPWR_M1004_d N_VPWR_M1018_d N_VPWR_M1022_d
+ N_VPWR_M1009_s N_VPWR_M1027_d N_VPWR_M1012_d N_VPWR_M1033_d VPWR
+ N_VPWR_c_1490_n N_VPWR_c_1493_n N_VPWR_c_1496_n N_VPWR_c_1499_n
+ N_VPWR_c_1502_n N_VPWR_c_1505_n N_VPWR_c_1508_n N_VPWR_c_1511_n
+ PM_SKY130_FD_SC_HVL__DFRBP_1%VPWR
x_PM_SKY130_FD_SC_HVL__DFRBP_1%A_509_608# N_A_509_608#_M1014_d
+ N_A_509_608#_M1018_s N_A_509_608#_M1008_d N_A_509_608#_c_1619_n
+ N_A_509_608#_c_1620_n N_A_509_608#_c_1621_n N_A_509_608#_c_1616_n
+ N_A_509_608#_c_1617_n N_A_509_608#_c_1623_n N_A_509_608#_c_1624_n
+ N_A_509_608#_c_1618_n N_A_509_608#_c_1670_n
+ PM_SKY130_FD_SC_HVL__DFRBP_1%A_509_608#
x_PM_SKY130_FD_SC_HVL__DFRBP_1%Q_N N_Q_N_M1017_d N_Q_N_M1023_d N_Q_N_c_1683_n
+ N_Q_N_c_1685_n Q_N Q_N Q_N N_Q_N_c_1684_n Q_N PM_SKY130_FD_SC_HVL__DFRBP_1%Q_N
x_PM_SKY130_FD_SC_HVL__DFRBP_1%Q N_Q_M1021_d N_Q_M1010_d Q Q Q Q Q Q Q
+ N_Q_c_1709_n PM_SKY130_FD_SC_HVL__DFRBP_1%Q
x_PM_SKY130_FD_SC_HVL__DFRBP_1%VGND N_VGND_M1020_d N_VGND_M1013_s N_VGND_M1029_d
+ N_VGND_M1007_d N_VGND_M1017_s N_VGND_M1024_d VGND N_VGND_c_1722_n
+ N_VGND_c_1724_n N_VGND_c_1726_n N_VGND_c_1728_n N_VGND_c_1730_n
+ N_VGND_c_1732_n N_VGND_c_1734_n PM_SKY130_FD_SC_HVL__DFRBP_1%VGND
cc_1 N_VNB_M1020_b N_CLK_M1020_g 0.124197f $X=-0.33 $Y=-0.265 $X2=0.72 $Y2=0.745
cc_2 N_VNB_c_2_p N_CLK_M1020_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.72 $Y2=0.745
cc_3 N_VNB_M1020_b N_A_37_107#_M1003_g 0.11788f $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=3.04
cc_4 N_VNB_c_2_p N_A_37_107#_M1003_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.72 $Y2=3.04
cc_5 N_VNB_M1020_b N_A_37_107#_M1006_g 0.0375635f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_M1020_b N_A_37_107#_c_290_n 0.0613139f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_7 N_VNB_M1020_b N_A_37_107#_c_291_n 0.0209007f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_8 N_VNB_c_2_p N_A_37_107#_c_291_n 8.17109e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_9 N_VNB_M1020_b N_A_37_107#_c_293_n 0.0458629f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_10 N_VNB_M1020_b N_A_37_107#_c_294_n 0.0200303f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1020_b N_A_37_107#_c_295_n 0.0024039f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1020_b N_A_37_107#_c_296_n 0.0142647f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1020_b N_A_37_107#_c_297_n 0.00488464f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_M1020_b N_A_37_107#_c_298_n 0.00857833f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_15 N_VNB_M1020_b N_A_37_107#_M1005_g 0.088947f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_16 N_VNB_M1020_b N_RESET_B_c_552_n 0.0438121f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_17 N_VNB_M1020_b N_RESET_B_M1025_g 0.0295649f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_18 N_VNB_M1020_b N_RESET_B_c_554_n 0.00911751f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_19 N_VNB_M1020_b N_RESET_B_c_555_n 0.16234f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_20 N_VNB_c_2_p N_RESET_B_c_555_n 0.00745873f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_21 N_VNB_M1020_b N_RESET_B_c_557_n 0.0076791f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_22 N_VNB_c_2_p N_RESET_B_c_557_n 4.18973e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_23 N_VNB_M1020_b N_RESET_B_c_559_n 0.00520894f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_24 N_VNB_M1020_b N_RESET_B_c_560_n 0.00647334f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_25 N_VNB_M1020_b N_RESET_B_c_561_n 0.00220419f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_26 N_VNB_M1020_b N_RESET_B_c_562_n 0.185623f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_27 N_VNB_c_2_p N_RESET_B_c_562_n 0.00863651f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_28 N_VNB_M1020_b N_RESET_B_c_564_n 0.0135577f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_29 N_VNB_c_2_p N_RESET_B_c_564_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_30 N_VNB_M1020_b N_RESET_B_c_566_n 0.00481238f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_31 N_VNB_M1020_b N_RESET_B_c_567_n 6.1416e-19 $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_32 N_VNB_M1020_b N_RESET_B_c_568_n 0.0467f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_33 N_VNB_M1020_b N_RESET_B_M1029_g 0.0848743f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_34 N_VNB_M1020_b N_RESET_B_c_570_n 0.0719739f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_35 N_VNB_M1020_b N_RESET_B_c_571_n 0.0357531f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_36 N_VNB_M1020_b N_D_c_746_n 0.0178776f $X=-0.33 $Y=-0.265 $X2=0.72 $Y2=3.04
cc_37 N_VNB_M1020_b N_D_M1014_g 0.0550252f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_38 N_VNB_M1020_b N_A_350_107#_c_796_n 0.0375799f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_39 N_VNB_M1020_b N_A_350_107#_c_797_n 0.0287947f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_M1020_b N_A_350_107#_c_798_n 0.0201578f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_41 N_VNB_M1020_b N_A_350_107#_c_799_n 0.00703171f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_42 N_VNB_M1020_b N_A_350_107#_c_800_n 0.029728f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_c_2_p N_A_350_107#_c_800_n 8.94283e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_44 N_VNB_M1020_b N_A_350_107#_c_802_n 0.00423199f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_45 N_VNB_M1020_b N_A_350_107#_c_803_n 0.0290394f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_M1020_b N_A_350_107#_c_804_n 0.0107717f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_47 N_VNB_M1020_b N_A_350_107#_c_805_n 0.0176161f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_M1020_b N_A_350_107#_c_806_n 0.00573325f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_49 N_VNB_M1020_b N_A_350_107#_c_807_n 0.00183994f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_M1020_b N_A_350_107#_c_808_n 0.00349603f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_51 N_VNB_M1020_b N_A_350_107#_M1028_g 0.0746712f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_52 N_VNB_M1020_b N_A_350_107#_c_810_n 0.0279405f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_53 N_VNB_M1020_b N_A_350_107#_c_811_n 0.0113251f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_54 N_VNB_M1020_b N_A_350_107#_c_812_n 0.0173397f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_55 N_VNB_M1020_b N_A_1176_466#_M1031_g 0.0415436f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_56 N_VNB_M1020_b N_A_1176_466#_c_984_n 0.0209602f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_57 N_VNB_M1020_b N_A_1176_466#_c_985_n 0.0178583f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_58 N_VNB_M1020_b N_A_1176_466#_c_986_n 0.00106385f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_59 N_VNB_M1020_b N_A_978_608#_c_1073_n 0.0432147f $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=3.04
cc_60 N_VNB_c_2_p N_A_978_608#_c_1073_n 5.98017e-19 $X=0.24 $Y=0 $X2=0.72
+ $Y2=3.04
cc_61 N_VNB_M1020_b N_A_978_608#_c_1075_n 7.19138e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_62 N_VNB_M1020_b N_A_978_608#_c_1076_n 0.00267229f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_63 N_VNB_M1020_b N_A_978_608#_c_1077_n 0.00388216f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_64 N_VNB_M1020_b N_A_978_608#_c_1078_n 0.00799773f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_65 N_VNB_M1020_b N_A_978_608#_c_1079_n 0.00575428f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_66 N_VNB_M1020_b N_A_978_608#_c_1080_n 0.00103536f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_67 N_VNB_M1020_b N_A_978_608#_c_1081_n 0.0747696f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_68 N_VNB_M1020_b N_A_2122_348#_c_1217_n 0.0206419f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_69 N_VNB_M1020_b N_A_2122_348#_c_1218_n 0.0157782f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_70 N_VNB_M1020_b N_A_2122_348#_c_1219_n 0.00771876f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_71 N_VNB_M1020_b N_A_2122_348#_c_1220_n 0.0184452f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_72 N_VNB_c_2_p N_A_2122_348#_c_1220_n 9.57246e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_73 N_VNB_M1020_b N_A_2122_348#_c_1222_n 0.00224001f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_74 N_VNB_M1020_b N_A_2122_348#_M1007_g 0.0983185f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_75 N_VNB_c_2_p N_A_2122_348#_M1007_g 8.54021e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_76 N_VNB_M1020_b N_A_1900_107#_M1001_g 0.102339f $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=3.04
cc_77 N_VNB_c_2_p N_A_1900_107#_M1001_g 0.0023273f $X=0.24 $Y=0 $X2=0.72
+ $Y2=3.04
cc_78 N_VNB_M1020_b N_A_1900_107#_c_1295_n 0.049186f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_79 N_VNB_M1020_b N_A_1900_107#_M1017_g 0.0526762f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_80 N_VNB_c_2_p N_A_1900_107#_M1017_g 0.00106379f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_81 N_VNB_M1020_b N_A_1900_107#_c_1298_n 0.0569497f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_82 N_VNB_M1020_b N_A_1900_107#_M1024_g 0.0474248f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_83 N_VNB_M1020_b N_A_1900_107#_c_1300_n 0.0173521f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_84 N_VNB_M1020_b N_A_1900_107#_c_1301_n 0.0392618f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_85 N_VNB_M1020_b N_A_1900_107#_c_1302_n 0.0087482f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_86 N_VNB_M1020_b N_A_1900_107#_c_1303_n 0.00184547f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_87 N_VNB_M1020_b N_A_1900_107#_c_1304_n 0.0235034f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_88 N_VNB_M1020_b N_A_2937_443#_M1021_g 0.0502106f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_89 N_VNB_c_2_p N_A_2937_443#_M1021_g 0.00112176f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_90 N_VNB_M1020_b N_A_2937_443#_c_1446_n 0.0113731f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_91 N_VNB_M1020_b N_A_2937_443#_c_1447_n 0.00693298f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_92 N_VNB_M1020_b N_A_2937_443#_c_1448_n 0.0518684f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_93 N_VNB_M1020_b N_A_2937_443#_c_1449_n 7.15764e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_94 N_VNB_M1020_b N_A_509_608#_c_1616_n 0.00225276f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_95 N_VNB_M1020_b N_A_509_608#_c_1617_n 0.00353466f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_96 N_VNB_M1020_b N_A_509_608#_c_1618_n 0.00160812f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_97 N_VNB_M1020_b N_Q_N_c_1683_n 0.00296361f $X=-0.33 $Y=-0.265 $X2=0.76
+ $Y2=1.28
cc_98 N_VNB_M1020_b N_Q_N_c_1684_n 0.0175611f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_99 N_VNB_M1020_b N_Q_c_1709_n 0.0638623f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_100 N_VNB_c_2_p N_Q_c_1709_n 8.87563e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_101 N_VNB_M1020_b N_VGND_c_1722_n 0.058257f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_102 N_VNB_c_2_p N_VGND_c_1722_n 0.00269373f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_103 N_VNB_M1020_b N_VGND_c_1724_n 0.086594f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_104 N_VNB_c_2_p N_VGND_c_1724_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_105 N_VNB_M1020_b N_VGND_c_1726_n 0.0591196f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_106 N_VNB_c_2_p N_VGND_c_1726_n 0.002699f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_107 N_VNB_M1020_b N_VGND_c_1728_n 0.0478209f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_108 N_VNB_c_2_p N_VGND_c_1728_n 0.00271358f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_109 N_VNB_M1020_b N_VGND_c_1730_n 0.0507186f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_110 N_VNB_c_2_p N_VGND_c_1730_n 0.00166879f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_111 N_VNB_M1020_b N_VGND_c_1732_n 0.0614104f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_112 N_VNB_c_2_p N_VGND_c_1732_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_113 N_VNB_M1020_b N_VGND_c_1734_n 0.24828f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_114 N_VNB_c_2_p N_VGND_c_1734_n 1.79618f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_115 N_VPB_M1004_b N_CLK_M1020_g 0.104299f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=0.745
cc_116 VPB N_CLK_M1020_g 5.12332e-19 $X=0 $Y=3.955 $X2=0.72 $Y2=0.745
cc_117 N_VPB_c_117_p N_CLK_M1020_g 0.00378627f $X=16.56 $Y=4.07 $X2=0.72
+ $Y2=0.745
cc_118 N_VPB_M1004_b N_A_37_107#_M1026_g 0.0426146f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_119 VPB N_A_37_107#_M1026_g 7.4229e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_120 N_VPB_c_117_p N_A_37_107#_M1026_g 0.00416825f $X=16.56 $Y=4.07 $X2=0
+ $Y2=0
cc_121 N_VPB_M1004_b N_A_37_107#_c_290_n 0.016181f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_122 N_VPB_M1004_b N_A_37_107#_c_304_n 0.0271453f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_123 N_VPB_M1004_b N_A_37_107#_c_305_n 0.0316893f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_124 N_VPB_M1004_b N_A_37_107#_c_293_n 0.0204685f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_125 N_VPB_M1004_b N_A_37_107#_c_307_n 0.0423859f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_126 VPB N_A_37_107#_c_307_n 4.92256e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_127 N_VPB_c_117_p N_A_37_107#_c_307_n 0.00490565f $X=16.56 $Y=4.07 $X2=0
+ $Y2=0
cc_128 N_VPB_M1004_b N_A_37_107#_c_310_n 0.0159465f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_129 N_VPB_M1004_b N_A_37_107#_c_294_n 0.0823777f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_130 N_VPB_M1004_b N_A_37_107#_c_312_n 0.00145965f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_131 N_VPB_M1004_b N_A_37_107#_c_313_n 0.0224752f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_132 VPB N_A_37_107#_c_313_n 0.0046234f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_133 N_VPB_c_117_p N_A_37_107#_c_313_n 0.0903565f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_134 N_VPB_M1004_b N_A_37_107#_c_316_n 0.0026545f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_135 VPB N_A_37_107#_c_316_n 5.70856e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_136 N_VPB_c_117_p N_A_37_107#_c_316_n 0.0114989f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_137 N_VPB_M1004_b N_A_37_107#_c_319_n 7.21626e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_138 N_VPB_M1004_b N_A_37_107#_c_320_n 0.00804031f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_139 N_VPB_M1004_b N_A_37_107#_c_321_n 0.0271059f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_140 VPB N_A_37_107#_c_321_n 0.00530737f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_141 N_VPB_c_117_p N_A_37_107#_c_321_n 0.0915483f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_142 N_VPB_M1004_b N_A_37_107#_c_324_n 0.00161351f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_143 VPB N_A_37_107#_c_324_n 5.41341e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_144 N_VPB_c_117_p N_A_37_107#_c_324_n 0.00961156f $X=16.56 $Y=4.07 $X2=0
+ $Y2=0
cc_145 N_VPB_M1004_b N_A_37_107#_c_327_n 0.0557294f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_146 VPB N_A_37_107#_c_327_n 4.55188e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_147 N_VPB_c_117_p N_A_37_107#_c_327_n 0.00306701f $X=16.56 $Y=4.07 $X2=0
+ $Y2=0
cc_148 N_VPB_M1004_b N_A_37_107#_c_330_n 0.00454397f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_149 N_VPB_M1004_b N_A_37_107#_c_331_n 5.15369e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_150 N_VPB_M1004_b N_A_37_107#_c_332_n 0.0127286f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_151 VPB N_A_37_107#_c_332_n 0.00235993f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_152 N_VPB_c_117_p N_A_37_107#_c_332_n 0.0462904f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_153 N_VPB_M1004_b N_A_37_107#_c_335_n 0.00237964f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_154 VPB N_A_37_107#_c_335_n 5.70856e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_155 N_VPB_c_117_p N_A_37_107#_c_335_n 0.0114989f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_156 N_VPB_M1004_b N_A_37_107#_c_338_n 0.0159462f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_157 N_VPB_M1004_b N_A_37_107#_c_339_n 0.00690145f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_158 N_VPB_M1004_b N_A_37_107#_c_340_n 0.00423891f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_159 N_VPB_M1004_b N_A_37_107#_c_296_n 0.0683657f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_160 N_VPB_c_117_p N_A_37_107#_c_296_n 0.0116928f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_161 N_VPB_M1004_b N_A_37_107#_c_343_n 0.00770964f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_162 N_VPB_M1004_b N_RESET_B_M1018_g 0.145066f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=0.745
cc_163 VPB N_RESET_B_M1018_g 5.4063e-19 $X=0 $Y=3.955 $X2=0.72 $Y2=0.745
cc_164 N_VPB_c_117_p N_RESET_B_M1018_g 0.00337783f $X=16.56 $Y=4.07 $X2=0.72
+ $Y2=0.745
cc_165 N_VPB_M1004_b N_RESET_B_c_575_n 0.0387328f $X=-0.33 $Y=1.885 $X2=0.76
+ $Y2=1.28
cc_166 VPB N_RESET_B_c_575_n 7.75595e-19 $X=0 $Y=3.955 $X2=0.76 $Y2=1.28
cc_167 N_VPB_c_117_p N_RESET_B_c_575_n 0.00451113f $X=16.56 $Y=4.07 $X2=0.76
+ $Y2=1.28
cc_168 N_VPB_M1004_b N_RESET_B_M1025_g 0.0675834f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_169 N_VPB_M1004_b N_RESET_B_c_579_n 0.0590788f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_170 N_VPB_M1004_b N_RESET_B_c_554_n 0.00482032f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_171 N_VPB_M1004_b N_RESET_B_c_561_n 0.00660262f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_172 N_VPB_M1004_b N_RESET_B_M1029_g 0.0759662f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_173 N_VPB_M1004_b N_RESET_B_c_570_n 0.00964338f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_174 N_VPB_M1004_b N_D_M1008_g 0.0624639f $X=-0.33 $Y=1.885 $X2=0.72 $Y2=0.745
cc_175 VPB N_D_M1008_g 5.4063e-19 $X=0 $Y=3.955 $X2=0.72 $Y2=0.745
cc_176 N_VPB_c_117_p N_D_M1008_g 0.00344615f $X=16.56 $Y=4.07 $X2=0.72 $Y2=0.745
cc_177 N_VPB_M1004_b N_D_c_751_n 0.0186385f $X=-0.33 $Y=1.885 $X2=0.76 $Y2=1.28
cc_178 N_VPB_M1004_b N_D_c_752_n 0.057111f $X=-0.33 $Y=1.885 $X2=0.76 $Y2=1.28
cc_179 N_VPB_M1004_b N_D_c_746_n 0.0077278f $X=-0.33 $Y=1.885 $X2=0.72 $Y2=3.04
cc_180 N_VPB_M1004_b N_A_350_107#_M1030_g 0.0382772f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=3.04
cc_181 N_VPB_M1004_b N_A_350_107#_c_799_n 0.0302569f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_182 N_VPB_M1004_b N_A_350_107#_c_815_n 0.00388265f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_183 N_VPB_M1004_b N_A_350_107#_c_816_n 0.083605f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_184 N_VPB_M1004_b N_A_350_107#_M1028_g 0.0308576f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_185 N_VPB_M1004_b N_A_350_107#_c_810_n 0.0369048f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_186 N_VPB_M1004_b N_A_350_107#_c_819_n 0.0425252f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_187 N_VPB_M1004_b N_A_1176_466#_c_987_n 0.0778316f $X=-0.33 $Y=1.885 $X2=0.76
+ $Y2=1.28
cc_188 N_VPB_M1004_b N_A_1176_466#_M1022_g 0.0339408f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=3.04
cc_189 N_VPB_c_117_p N_A_1176_466#_M1022_g 0.00212077f $X=16.56 $Y=4.07 $X2=0.72
+ $Y2=3.04
cc_190 N_VPB_M1004_b N_A_1176_466#_c_985_n 0.0399334f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_191 N_VPB_M1004_b N_A_1176_466#_c_991_n 0.0173253f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_192 N_VPB_M1004_b N_A_978_608#_M1009_g 0.0654068f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_193 N_VPB_c_117_p N_A_978_608#_M1009_g 0.0015607f $X=16.56 $Y=4.07 $X2=0
+ $Y2=0
cc_194 N_VPB_M1004_b N_A_978_608#_c_1084_n 0.011425f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_195 N_VPB_M1004_b N_A_978_608#_c_1085_n 0.00201778f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_196 N_VPB_M1004_b N_A_978_608#_c_1077_n 0.00789613f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_197 N_VPB_M1004_b N_A_978_608#_c_1087_n 0.00605308f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_198 N_VPB_M1004_b N_A_978_608#_c_1088_n 0.00167087f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_199 N_VPB_M1004_b N_A_978_608#_c_1089_n 0.00398331f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_200 N_VPB_M1004_b N_A_978_608#_c_1090_n 0.00424815f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_201 N_VPB_M1004_b N_A_978_608#_c_1091_n 7.77693e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_202 N_VPB_M1004_b N_A_978_608#_c_1081_n 0.0128022f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_203 N_VPB_M1004_b N_A_2122_348#_c_1217_n 0.069327f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_204 N_VPB_M1004_b N_A_2122_348#_c_1226_n 0.0024289f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_205 N_VPB_M1004_b N_A_2122_348#_c_1227_n 0.010754f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_206 N_VPB_M1004_b N_A_1900_107#_c_1305_n 0.044955f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_207 N_VPB_M1004_b N_A_1900_107#_c_1295_n 0.0375769f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_208 N_VPB_M1004_b N_A_1900_107#_M1023_g 0.043718f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_209 VPB N_A_1900_107#_M1023_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_210 N_VPB_c_117_p N_A_1900_107#_M1023_g 0.0152133f $X=16.56 $Y=4.07 $X2=0
+ $Y2=0
cc_211 N_VPB_M1004_b N_A_1900_107#_c_1298_n 0.0455069f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_212 N_VPB_M1004_b N_A_1900_107#_M1033_g 0.043238f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_213 N_VPB_M1004_b N_A_1900_107#_c_1300_n 0.0115681f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_214 N_VPB_M1004_b N_A_1900_107#_c_1301_n 0.0162118f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_215 N_VPB_M1004_b N_A_1900_107#_c_1314_n 0.00228659f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_216 N_VPB_M1004_b N_A_1900_107#_c_1315_n 0.0230028f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_217 N_VPB_c_117_p N_A_1900_107#_c_1315_n 0.00319597f $X=16.56 $Y=4.07 $X2=0
+ $Y2=0
cc_218 N_VPB_M1004_b N_A_1900_107#_c_1317_n 4.85926e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_219 N_VPB_M1004_b N_A_1900_107#_c_1302_n 9.99362e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_220 N_VPB_M1004_b N_A_1900_107#_c_1319_n 0.0085255f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_221 N_VPB_M1004_b N_A_1900_107#_c_1320_n 0.0100512f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_222 N_VPB_M1004_b N_A_1900_107#_c_1304_n 0.0282881f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_223 N_VPB_M1004_b N_A_2937_443#_M1010_g 0.0603943f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=3.04
cc_224 VPB N_A_2937_443#_M1010_g 0.00970178f $X=0 $Y=3.955 $X2=0.72 $Y2=3.04
cc_225 N_VPB_c_117_p N_A_2937_443#_M1010_g 0.0162989f $X=16.56 $Y=4.07 $X2=0.72
+ $Y2=3.04
cc_226 N_VPB_M1004_b N_A_2937_443#_c_1453_n 0.0143335f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_227 N_VPB_M1004_b N_A_2937_443#_c_1448_n 0.00537205f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_228 N_VPB_M1004_b N_VPWR_c_1490_n 0.0128551f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1490_n 0.00252021f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_230 N_VPB_c_117_p N_VPWR_c_1490_n 0.0384021f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_231 N_VPB_M1004_b N_VPWR_c_1493_n 0.00646826f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1493_n 4.76526e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_233 N_VPB_c_117_p N_VPWR_c_1493_n 0.00726955f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_234 N_VPB_M1004_b N_VPWR_c_1496_n 0.0062288f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1496_n 0.0026787f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_236 N_VPB_c_117_p N_VPWR_c_1496_n 0.0402679f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_237 N_VPB_M1004_b N_VPWR_c_1499_n 0.0194912f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1499_n 0.00269208f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_239 N_VPB_c_117_p N_VPWR_c_1499_n 0.0409717f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_240 N_VPB_M1004_b N_VPWR_c_1502_n 0.0844032f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1502_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_242 N_VPB_c_117_p N_VPWR_c_1502_n 0.0409968f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_243 N_VPB_M1004_b N_VPWR_c_1505_n 0.0487725f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1505_n 0.00337025f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_245 N_VPB_c_117_p N_VPWR_c_1505_n 0.0454439f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_246 N_VPB_M1004_b N_VPWR_c_1508_n 0.0332888f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1508_n 0.00335473f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_248 N_VPB_c_117_p N_VPWR_c_1508_n 0.0490696f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_249 N_VPB_M1004_b N_VPWR_c_1511_n 0.241938f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1511_n 1.79413f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_251 N_VPB_c_117_p N_VPWR_c_1511_n 0.0842164f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_252 N_VPB_M1004_b N_A_509_608#_c_1619_n 0.0111022f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_253 N_VPB_M1004_b N_A_509_608#_c_1620_n 0.00752592f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_254 N_VPB_M1004_b N_A_509_608#_c_1621_n 0.00831093f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_255 N_VPB_M1004_b N_A_509_608#_c_1617_n 0.0048719f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_256 N_VPB_M1004_b N_A_509_608#_c_1623_n 0.0048816f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_257 N_VPB_M1004_b N_A_509_608#_c_1624_n 0.00290633f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_258 N_VPB_M1004_b N_Q_N_c_1685_n 0.0298952f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=3.04
cc_259 VPB N_Q_N_c_1685_n 7.60114e-19 $X=0 $Y=3.955 $X2=0.72 $Y2=3.04
cc_260 N_VPB_c_117_p N_Q_N_c_1685_n 0.0131049f $X=16.56 $Y=4.07 $X2=0.72
+ $Y2=3.04
cc_261 N_VPB_M1004_b N_Q_c_1709_n 0.0679775f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_262 VPB N_Q_c_1709_n 0.00110823f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_263 N_VPB_c_117_p N_Q_c_1709_n 0.0182942f $X=16.56 $Y=4.07 $X2=0 $Y2=0
cc_264 CLK N_A_37_107#_M1003_g 0.0035357f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_265 N_CLK_M1020_g N_A_37_107#_M1003_g 0.0952851f $X=0.72 $Y=0.745 $X2=0 $Y2=0
cc_266 N_CLK_M1020_g N_A_37_107#_M1026_g 0.0149043f $X=0.72 $Y=0.745 $X2=0 $Y2=0
cc_267 N_CLK_M1020_g N_A_37_107#_c_291_n 0.00602693f $X=0.72 $Y=0.745 $X2=0
+ $Y2=0
cc_268 CLK N_A_37_107#_c_293_n 0.0404148f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_269 N_CLK_M1020_g N_A_37_107#_c_293_n 0.0497587f $X=0.72 $Y=0.745 $X2=0 $Y2=0
cc_270 N_CLK_M1020_g N_A_37_107#_c_307_n 0.0133556f $X=0.72 $Y=0.745 $X2=0 $Y2=0
cc_271 CLK N_A_37_107#_c_310_n 0.00924969f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_272 N_CLK_M1020_g N_A_37_107#_c_310_n 0.0403226f $X=0.72 $Y=0.745 $X2=0 $Y2=0
cc_273 N_CLK_M1020_g N_A_37_107#_c_353_n 0.00165588f $X=0.72 $Y=0.745 $X2=0
+ $Y2=0
cc_274 N_CLK_M1020_g N_A_37_107#_c_312_n 9.82494e-19 $X=0.72 $Y=0.745 $X2=0
+ $Y2=0
cc_275 N_CLK_M1020_g N_A_37_107#_c_298_n 0.00506999f $X=0.72 $Y=0.745 $X2=0
+ $Y2=0
cc_276 N_CLK_M1020_g N_VPWR_c_1490_n 0.0583784f $X=0.72 $Y=0.745 $X2=0 $Y2=0
cc_277 N_CLK_M1020_g N_VPWR_c_1511_n 0.00856946f $X=0.72 $Y=0.745 $X2=0 $Y2=0
cc_278 CLK N_VGND_c_1722_n 0.0189446f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_279 N_CLK_M1020_g N_VGND_c_1722_n 0.0374903f $X=0.72 $Y=0.745 $X2=0 $Y2=0
cc_280 CLK N_VGND_c_1734_n 0.00340663f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_281 N_CLK_M1020_g N_VGND_c_1734_n 0.00922972f $X=0.72 $Y=0.745 $X2=0 $Y2=0
cc_282 N_A_37_107#_c_313_n N_RESET_B_M1018_g 0.00730215f $X=3.035 $Y=3.72 $X2=0
+ $Y2=0
cc_283 N_A_37_107#_c_319_n N_RESET_B_M1018_g 0.0347699f $X=3.12 $Y=3.635 $X2=0
+ $Y2=0
cc_284 N_A_37_107#_c_320_n N_RESET_B_M1018_g 0.0111916f $X=3.735 $Y=2.735 $X2=0
+ $Y2=0
cc_285 N_A_37_107#_c_359_p N_RESET_B_M1018_g 0.00779832f $X=3.205 $Y=2.735 $X2=0
+ $Y2=0
cc_286 N_A_37_107#_c_360_p N_RESET_B_M1018_g 8.83283e-19 $X=3.82 $Y=3.6 $X2=0
+ $Y2=0
cc_287 N_A_37_107#_c_330_n N_RESET_B_c_575_n 0.0100851f $X=6.865 $Y=2.96 $X2=0
+ $Y2=0
cc_288 N_A_37_107#_c_331_n N_RESET_B_c_575_n 0.0237719f $X=6.95 $Y=3.635 $X2=0
+ $Y2=0
cc_289 N_A_37_107#_c_332_n N_RESET_B_c_575_n 0.00465098f $X=7.565 $Y=3.72 $X2=0
+ $Y2=0
cc_290 N_A_37_107#_c_338_n N_RESET_B_c_575_n 0.00251846f $X=7.65 $Y=3.635 $X2=0
+ $Y2=0
cc_291 N_A_37_107#_c_330_n N_RESET_B_c_579_n 0.00858417f $X=6.865 $Y=2.96
+ $X2=8.4 $Y2=0
cc_292 N_A_37_107#_c_338_n N_RESET_B_c_579_n 9.45457e-19 $X=7.65 $Y=3.635
+ $X2=8.4 $Y2=0
cc_293 N_A_37_107#_c_340_n N_RESET_B_c_579_n 0.00288729f $X=7.735 $Y=2.785
+ $X2=8.4 $Y2=0
cc_294 N_A_37_107#_M1006_g N_RESET_B_c_555_n 0.0218926f $X=4.88 $Y=1.075 $X2=0
+ $Y2=0
cc_295 N_A_37_107#_M1005_g N_RESET_B_c_562_n 0.01476f $X=10.32 $Y=0.745 $X2=0
+ $Y2=0
cc_296 N_A_37_107#_M1005_g N_RESET_B_c_598_n 0.00175194f $X=10.32 $Y=0.745 $X2=0
+ $Y2=0
cc_297 N_A_37_107#_c_319_n N_D_M1008_g 8.83283e-19 $X=3.12 $Y=3.635 $X2=0 $Y2=0
cc_298 N_A_37_107#_c_320_n N_D_M1008_g 0.0190932f $X=3.735 $Y=2.735 $X2=0 $Y2=0
cc_299 N_A_37_107#_c_360_p N_D_M1008_g 0.0340448f $X=3.82 $Y=3.6 $X2=0 $Y2=0
cc_300 N_A_37_107#_c_321_n N_D_M1008_g 0.00774274f $X=5.395 $Y=3.685 $X2=0 $Y2=0
cc_301 N_A_37_107#_c_290_n N_D_c_746_n 0.0187614f $X=4.997 $Y=1.915 $X2=0.24
+ $Y2=0
cc_302 N_A_37_107#_M1006_g D 2.44045e-19 $X=4.88 $Y=1.075 $X2=0.24 $Y2=0
cc_303 N_A_37_107#_M1006_g N_D_M1014_g 0.0187614f $X=4.88 $Y=1.075 $X2=16.56
+ $Y2=0
cc_304 N_A_37_107#_c_360_p N_A_350_107#_M1030_g 0.00112553f $X=3.82 $Y=3.6 $X2=0
+ $Y2=0
cc_305 N_A_37_107#_c_321_n N_A_350_107#_M1030_g 0.0175848f $X=5.395 $Y=3.685
+ $X2=0 $Y2=0
cc_306 N_A_37_107#_c_327_n N_A_350_107#_M1030_g 0.0140517f $X=5.485 $Y=2.715
+ $X2=0 $Y2=0
cc_307 N_A_37_107#_c_381_p N_A_350_107#_M1030_g 0.00105516f $X=5.48 $Y=3.6 $X2=0
+ $Y2=0
cc_308 N_A_37_107#_c_297_n N_A_350_107#_c_796_n 0.00804347f $X=10.09 $Y=1.315
+ $X2=0.24 $Y2=0
cc_309 N_A_37_107#_c_383_p N_A_350_107#_c_796_n 0.00978694f $X=9.375 $Y=1.315
+ $X2=0.24 $Y2=0
cc_310 N_A_37_107#_c_384_p N_A_350_107#_c_796_n 0.00103296f $X=10.255 $Y=1.235
+ $X2=0.24 $Y2=0
cc_311 N_A_37_107#_M1005_g N_A_350_107#_c_796_n 0.0188856f $X=10.32 $Y=0.745
+ $X2=0.24 $Y2=0
cc_312 N_A_37_107#_c_297_n N_A_350_107#_c_797_n 0.0114225f $X=10.09 $Y=1.315
+ $X2=0 $Y2=0
cc_313 N_A_37_107#_M1005_g N_A_350_107#_c_797_n 0.0103535f $X=10.32 $Y=0.745
+ $X2=0 $Y2=0
cc_314 N_A_37_107#_c_295_n N_A_350_107#_c_798_n 0.011277f $X=9.29 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_A_37_107#_c_296_n N_A_350_107#_c_798_n 0.0367675f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_316 N_A_37_107#_c_297_n N_A_350_107#_c_798_n 7.2577e-19 $X=10.09 $Y=1.315
+ $X2=0 $Y2=0
cc_317 N_A_37_107#_c_353_n N_A_350_107#_c_799_n 0.0278582f $X=1.67 $Y=2 $X2=0
+ $Y2=0
cc_318 N_A_37_107#_c_294_n N_A_350_107#_c_799_n 0.0310609f $X=1.67 $Y=2 $X2=0
+ $Y2=0
cc_319 N_A_37_107#_c_312_n N_A_350_107#_c_799_n 0.0425078f $X=1.75 $Y=3.635
+ $X2=0 $Y2=0
cc_320 N_A_37_107#_c_313_n N_A_350_107#_c_799_n 0.0176725f $X=3.035 $Y=3.72
+ $X2=0 $Y2=0
cc_321 N_A_37_107#_c_395_p N_A_350_107#_c_799_n 0.0134164f $X=1.67 $Y=2.36 $X2=0
+ $Y2=0
cc_322 N_A_37_107#_c_290_n N_A_350_107#_c_815_n 0.0101713f $X=4.997 $Y=1.915
+ $X2=0 $Y2=0
cc_323 N_A_37_107#_c_305_n N_A_350_107#_c_815_n 0.00747067f $X=5.42 $Y=2.41
+ $X2=0 $Y2=0
cc_324 N_A_37_107#_c_290_n N_A_350_107#_c_816_n 0.0232749f $X=4.997 $Y=1.915
+ $X2=0 $Y2=0
cc_325 N_A_37_107#_c_305_n N_A_350_107#_c_816_n 0.050556f $X=5.42 $Y=2.41 $X2=0
+ $Y2=0
cc_326 N_A_37_107#_M1003_g N_A_350_107#_c_800_n 0.00275918f $X=1.5 $Y=0.745
+ $X2=0 $Y2=0
cc_327 N_A_37_107#_c_290_n N_A_350_107#_c_843_n 0.0144976f $X=4.997 $Y=1.915
+ $X2=0 $Y2=0
cc_328 N_A_37_107#_c_290_n N_A_350_107#_c_844_n 0.00183185f $X=4.997 $Y=1.915
+ $X2=0 $Y2=0
cc_329 N_A_37_107#_c_290_n N_A_350_107#_c_802_n 0.0429192f $X=4.997 $Y=1.915
+ $X2=0 $Y2=0
cc_330 N_A_37_107#_c_290_n N_A_350_107#_c_803_n 0.00390195f $X=4.997 $Y=1.915
+ $X2=0 $Y2=0
cc_331 N_A_37_107#_M1003_g N_A_350_107#_c_804_n 0.00679362f $X=1.5 $Y=0.745
+ $X2=0 $Y2=0
cc_332 N_A_37_107#_c_295_n N_A_350_107#_c_805_n 0.0147789f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_333 N_A_37_107#_c_296_n N_A_350_107#_c_805_n 0.00439311f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_334 N_A_37_107#_c_297_n N_A_350_107#_c_805_n 0.0129217f $X=10.09 $Y=1.315
+ $X2=0 $Y2=0
cc_335 N_A_37_107#_c_290_n N_A_350_107#_c_851_n 0.00582843f $X=4.997 $Y=1.915
+ $X2=0 $Y2=0
cc_336 N_A_37_107#_c_295_n N_A_350_107#_c_807_n 0.002581f $X=9.29 $Y=1.985 $X2=0
+ $Y2=0
cc_337 N_A_37_107#_c_297_n N_A_350_107#_c_807_n 0.00796764f $X=10.09 $Y=1.315
+ $X2=0 $Y2=0
cc_338 N_A_37_107#_c_295_n N_A_350_107#_c_808_n 0.0185074f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_339 N_A_37_107#_c_296_n N_A_350_107#_c_808_n 0.00115691f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_340 N_A_37_107#_c_297_n N_A_350_107#_c_808_n 0.0213394f $X=10.09 $Y=1.315
+ $X2=0 $Y2=0
cc_341 N_A_37_107#_M1006_g N_A_350_107#_M1028_g 0.013837f $X=4.88 $Y=1.075 $X2=0
+ $Y2=0
cc_342 N_A_37_107#_c_290_n N_A_350_107#_M1028_g 0.0497914f $X=4.997 $Y=1.915
+ $X2=0 $Y2=0
cc_343 N_A_37_107#_c_304_n N_A_350_107#_M1028_g 0.00400771f $X=5.42 $Y=2.66
+ $X2=0 $Y2=0
cc_344 N_A_37_107#_c_295_n N_A_350_107#_c_810_n 0.00160991f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_345 N_A_37_107#_c_296_n N_A_350_107#_c_810_n 0.0280569f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_346 N_A_37_107#_c_297_n N_A_350_107#_c_810_n 0.00143484f $X=10.09 $Y=1.315
+ $X2=0 $Y2=0
cc_347 N_A_37_107#_c_384_p N_A_350_107#_c_810_n 0.001357f $X=10.255 $Y=1.235
+ $X2=0 $Y2=0
cc_348 N_A_37_107#_M1005_g N_A_350_107#_c_810_n 0.0247338f $X=10.32 $Y=0.745
+ $X2=0 $Y2=0
cc_349 N_A_37_107#_c_295_n N_A_350_107#_c_811_n 0.00289391f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_350 N_A_37_107#_c_295_n N_A_350_107#_c_819_n 5.55519e-19 $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_351 N_A_37_107#_c_296_n N_A_350_107#_c_819_n 0.0109215f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_352 N_A_37_107#_M1003_g N_A_350_107#_c_812_n 0.0285165f $X=1.5 $Y=0.745 $X2=0
+ $Y2=0
cc_353 N_A_37_107#_c_339_n N_A_1176_466#_M1009_d 0.00430106f $X=9.205 $Y=2.785
+ $X2=0 $Y2=0
cc_354 N_A_37_107#_c_304_n N_A_1176_466#_c_987_n 0.0407688f $X=5.42 $Y=2.66
+ $X2=0 $Y2=0
cc_355 N_A_37_107#_c_305_n N_A_1176_466#_c_987_n 0.00184888f $X=5.42 $Y=2.41
+ $X2=0 $Y2=0
cc_356 N_A_37_107#_c_430_p N_A_1176_466#_c_987_n 0.00190692f $X=5.485 $Y=2.715
+ $X2=0 $Y2=0
cc_357 N_A_37_107#_c_330_n N_A_1176_466#_c_987_n 0.0140965f $X=6.865 $Y=2.96
+ $X2=0 $Y2=0
cc_358 N_A_37_107#_c_327_n N_A_1176_466#_M1022_g 0.0407688f $X=5.485 $Y=2.715
+ $X2=0 $Y2=0
cc_359 N_A_37_107#_c_381_p N_A_1176_466#_M1022_g 0.00142735f $X=5.48 $Y=3.6
+ $X2=0 $Y2=0
cc_360 N_A_37_107#_c_330_n N_A_1176_466#_M1022_g 0.0160235f $X=6.865 $Y=2.96
+ $X2=0 $Y2=0
cc_361 N_A_37_107#_c_331_n N_A_1176_466#_M1022_g 8.03185e-19 $X=6.95 $Y=3.635
+ $X2=0 $Y2=0
cc_362 N_A_37_107#_c_339_n N_A_1176_466#_c_991_n 0.0365002f $X=9.205 $Y=2.785
+ $X2=0 $Y2=0
cc_363 N_A_37_107#_c_340_n N_A_1176_466#_c_991_n 0.00861088f $X=7.735 $Y=2.785
+ $X2=0 $Y2=0
cc_364 N_A_37_107#_c_295_n N_A_1176_466#_c_986_n 0.0767638f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_365 N_A_37_107#_c_296_n N_A_1176_466#_c_986_n 0.0108082f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_366 N_A_37_107#_c_383_p N_A_1176_466#_c_986_n 0.0128825f $X=9.375 $Y=1.315
+ $X2=0 $Y2=0
cc_367 N_A_37_107#_c_339_n N_A_1176_466#_c_1006_n 0.0163515f $X=9.205 $Y=2.785
+ $X2=0 $Y2=0
cc_368 N_A_37_107#_c_296_n N_A_1176_466#_c_1006_n 0.00768216f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_369 N_A_37_107#_c_338_n N_A_978_608#_M1009_g 0.00392464f $X=7.65 $Y=3.635
+ $X2=0 $Y2=0
cc_370 N_A_37_107#_c_339_n N_A_978_608#_M1009_g 0.0304058f $X=9.205 $Y=2.785
+ $X2=0 $Y2=0
cc_371 N_A_37_107#_c_295_n N_A_978_608#_M1009_g 5.99284e-19 $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_372 N_A_37_107#_c_304_n N_A_978_608#_c_1084_n 0.00800423f $X=5.42 $Y=2.66
+ $X2=0 $Y2=0
cc_373 N_A_37_107#_c_305_n N_A_978_608#_c_1084_n 0.0160578f $X=5.42 $Y=2.41
+ $X2=0 $Y2=0
cc_374 N_A_37_107#_c_430_p N_A_978_608#_c_1084_n 0.0191957f $X=5.485 $Y=2.715
+ $X2=0 $Y2=0
cc_375 N_A_37_107#_c_330_n N_A_978_608#_c_1084_n 0.0143192f $X=6.865 $Y=2.96
+ $X2=0 $Y2=0
cc_376 N_A_37_107#_c_290_n N_A_978_608#_c_1085_n 0.00329456f $X=4.997 $Y=1.915
+ $X2=0 $Y2=0
cc_377 N_A_37_107#_c_305_n N_A_978_608#_c_1085_n 0.00262624f $X=5.42 $Y=2.41
+ $X2=0 $Y2=0
cc_378 N_A_37_107#_c_304_n N_A_978_608#_c_1102_n 5.34958e-19 $X=5.42 $Y=2.66
+ $X2=0 $Y2=0
cc_379 N_A_37_107#_c_330_n N_A_978_608#_c_1087_n 0.0520926f $X=6.865 $Y=2.96
+ $X2=0 $Y2=0
cc_380 N_A_37_107#_c_304_n N_A_978_608#_c_1104_n 5.03523e-19 $X=5.42 $Y=2.66
+ $X2=0 $Y2=0
cc_381 N_A_37_107#_c_430_p N_A_978_608#_c_1104_n 0.00508234f $X=5.485 $Y=2.715
+ $X2=0 $Y2=0
cc_382 N_A_37_107#_c_330_n N_A_978_608#_c_1104_n 0.0123662f $X=6.865 $Y=2.96
+ $X2=0 $Y2=0
cc_383 N_A_37_107#_c_330_n N_A_978_608#_c_1088_n 0.0125408f $X=6.865 $Y=2.96
+ $X2=0 $Y2=0
cc_384 N_A_37_107#_c_331_n N_A_978_608#_c_1088_n 0.0133874f $X=6.95 $Y=3.635
+ $X2=0 $Y2=0
cc_385 N_A_37_107#_c_332_n N_A_978_608#_c_1088_n 0.0112524f $X=7.565 $Y=3.72
+ $X2=0 $Y2=0
cc_386 N_A_37_107#_c_338_n N_A_978_608#_c_1088_n 0.0414296f $X=7.65 $Y=3.635
+ $X2=0 $Y2=0
cc_387 N_A_37_107#_c_340_n N_A_978_608#_c_1088_n 0.0131377f $X=7.735 $Y=2.785
+ $X2=0 $Y2=0
cc_388 N_A_37_107#_c_321_n N_A_978_608#_c_1089_n 0.0188079f $X=5.395 $Y=3.685
+ $X2=0 $Y2=0
cc_389 N_A_37_107#_c_327_n N_A_978_608#_c_1089_n 0.0086799f $X=5.485 $Y=2.715
+ $X2=0 $Y2=0
cc_390 N_A_37_107#_c_381_p N_A_978_608#_c_1089_n 0.0256692f $X=5.48 $Y=3.6 $X2=0
+ $Y2=0
cc_391 N_A_37_107#_c_304_n N_A_978_608#_c_1090_n 0.00661301f $X=5.42 $Y=2.66
+ $X2=0 $Y2=0
cc_392 N_A_37_107#_c_305_n N_A_978_608#_c_1090_n 0.00105638f $X=5.42 $Y=2.41
+ $X2=0 $Y2=0
cc_393 N_A_37_107#_c_430_p N_A_978_608#_c_1090_n 0.0216168f $X=5.485 $Y=2.715
+ $X2=0 $Y2=0
cc_394 N_A_37_107#_c_327_n N_A_978_608#_c_1090_n 0.00786869f $X=5.485 $Y=2.715
+ $X2=0 $Y2=0
cc_395 N_A_37_107#_c_469_p N_A_978_608#_c_1090_n 0.0125052f $X=5.522 $Y=2.96
+ $X2=0 $Y2=0
cc_396 N_A_37_107#_M1006_g N_A_978_608#_c_1079_n 0.00758143f $X=4.88 $Y=1.075
+ $X2=0 $Y2=0
cc_397 N_A_37_107#_c_290_n N_A_978_608#_c_1079_n 0.00280787f $X=4.997 $Y=1.915
+ $X2=0 $Y2=0
cc_398 N_A_37_107#_c_295_n N_A_978_608#_c_1081_n 0.00116227f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_399 N_A_37_107#_c_296_n N_A_978_608#_c_1081_n 0.0631167f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_400 N_A_37_107#_M1005_g N_A_2122_348#_M1007_g 0.0732905f $X=10.32 $Y=0.745
+ $X2=0 $Y2=0
cc_401 N_A_37_107#_c_297_n N_A_1900_107#_M1016_d 0.0025225f $X=10.09 $Y=1.315
+ $X2=0 $Y2=0
cc_402 N_A_37_107#_c_295_n N_A_1900_107#_c_1314_n 0.00727363f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_403 N_A_37_107#_c_296_n N_A_1900_107#_c_1314_n 4.57034e-19 $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_404 N_A_37_107#_c_296_n N_A_1900_107#_c_1315_n 0.00184621f $X=9.29 $Y=1.985
+ $X2=0 $Y2=0
cc_405 N_A_37_107#_c_297_n N_A_1900_107#_c_1326_n 0.00448304f $X=10.09 $Y=1.315
+ $X2=0 $Y2=0
cc_406 N_A_37_107#_c_384_p N_A_1900_107#_c_1326_n 0.0118001f $X=10.255 $Y=1.235
+ $X2=0 $Y2=0
cc_407 N_A_37_107#_M1005_g N_A_1900_107#_c_1326_n 0.0294086f $X=10.32 $Y=0.745
+ $X2=0 $Y2=0
cc_408 N_A_37_107#_c_384_p N_A_1900_107#_c_1302_n 0.0222477f $X=10.255 $Y=1.235
+ $X2=0 $Y2=0
cc_409 N_A_37_107#_M1005_g N_A_1900_107#_c_1302_n 0.0213242f $X=10.32 $Y=0.745
+ $X2=0 $Y2=0
cc_410 N_A_37_107#_c_384_p N_A_1900_107#_c_1320_n 0.00363417f $X=10.255 $Y=1.235
+ $X2=0 $Y2=0
cc_411 N_A_37_107#_M1005_g N_A_1900_107#_c_1320_n 0.0053771f $X=10.32 $Y=0.745
+ $X2=0 $Y2=0
cc_412 N_A_37_107#_c_297_n N_A_1900_107#_c_1303_n 0.0181887f $X=10.09 $Y=1.315
+ $X2=0 $Y2=0
cc_413 N_A_37_107#_M1005_g N_A_1900_107#_c_1303_n 0.00343208f $X=10.32 $Y=0.745
+ $X2=0 $Y2=0
cc_414 N_A_37_107#_c_330_n N_VPWR_M1022_d 0.00174261f $X=6.865 $Y=2.96 $X2=0
+ $Y2=0
cc_415 N_A_37_107#_c_339_n N_VPWR_M1009_s 0.00685713f $X=9.205 $Y=2.785 $X2=0
+ $Y2=0
cc_416 N_A_37_107#_M1026_g N_VPWR_c_1490_n 0.0322309f $X=1.71 $Y=3.04 $X2=0
+ $Y2=0
cc_417 N_A_37_107#_c_307_n N_VPWR_c_1490_n 0.036089f $X=0.33 $Y=2.79 $X2=0 $Y2=0
cc_418 N_A_37_107#_c_310_n N_VPWR_c_1490_n 0.0678906f $X=1.505 $Y=2.36 $X2=0
+ $Y2=0
cc_419 N_A_37_107#_c_294_n N_VPWR_c_1490_n 0.00633626f $X=1.67 $Y=2 $X2=0 $Y2=0
cc_420 N_A_37_107#_c_312_n N_VPWR_c_1490_n 0.0716056f $X=1.75 $Y=3.635 $X2=0
+ $Y2=0
cc_421 N_A_37_107#_c_316_n N_VPWR_c_1490_n 0.00489946f $X=1.835 $Y=3.72 $X2=0
+ $Y2=0
cc_422 N_A_37_107#_c_313_n N_VPWR_c_1493_n 0.00479486f $X=3.035 $Y=3.72 $X2=0
+ $Y2=0
cc_423 N_A_37_107#_c_319_n N_VPWR_c_1493_n 0.0277594f $X=3.12 $Y=3.635 $X2=0
+ $Y2=0
cc_424 N_A_37_107#_c_320_n N_VPWR_c_1493_n 0.0136666f $X=3.735 $Y=2.735 $X2=0
+ $Y2=0
cc_425 N_A_37_107#_c_360_p N_VPWR_c_1493_n 0.0254272f $X=3.82 $Y=3.6 $X2=0 $Y2=0
cc_426 N_A_37_107#_c_324_n N_VPWR_c_1493_n 0.00719229f $X=3.905 $Y=3.685 $X2=0
+ $Y2=0
cc_427 N_A_37_107#_c_321_n N_VPWR_c_1496_n 0.0073198f $X=5.395 $Y=3.685 $X2=0
+ $Y2=0
cc_428 N_A_37_107#_c_327_n N_VPWR_c_1496_n 0.00260875f $X=5.485 $Y=2.715 $X2=0
+ $Y2=0
cc_429 N_A_37_107#_c_381_p N_VPWR_c_1496_n 0.0266834f $X=5.48 $Y=3.6 $X2=0 $Y2=0
cc_430 N_A_37_107#_c_330_n N_VPWR_c_1496_n 0.0523546f $X=6.865 $Y=2.96 $X2=0
+ $Y2=0
cc_431 N_A_37_107#_c_331_n N_VPWR_c_1496_n 0.0279156f $X=6.95 $Y=3.635 $X2=0
+ $Y2=0
cc_432 N_A_37_107#_c_335_n N_VPWR_c_1496_n 0.00485641f $X=7.035 $Y=3.72 $X2=0
+ $Y2=0
cc_433 N_A_37_107#_c_332_n N_VPWR_c_1499_n 0.00489946f $X=7.565 $Y=3.72 $X2=0
+ $Y2=0
cc_434 N_A_37_107#_c_338_n N_VPWR_c_1499_n 0.0448205f $X=7.65 $Y=3.635 $X2=0
+ $Y2=0
cc_435 N_A_37_107#_c_339_n N_VPWR_c_1499_n 0.060499f $X=9.205 $Y=2.785 $X2=0
+ $Y2=0
cc_436 N_A_37_107#_c_296_n N_VPWR_c_1499_n 0.0116259f $X=9.29 $Y=1.985 $X2=0
+ $Y2=0
cc_437 N_A_37_107#_M1026_g N_VPWR_c_1511_n 0.0192291f $X=1.71 $Y=3.04 $X2=0
+ $Y2=0
cc_438 N_A_37_107#_c_307_n N_VPWR_c_1511_n 0.0199094f $X=0.33 $Y=2.79 $X2=0
+ $Y2=0
cc_439 N_A_37_107#_c_312_n N_VPWR_c_1511_n 0.0206969f $X=1.75 $Y=3.635 $X2=0
+ $Y2=0
cc_440 N_A_37_107#_c_313_n N_VPWR_c_1511_n 0.054585f $X=3.035 $Y=3.72 $X2=0
+ $Y2=0
cc_441 N_A_37_107#_c_316_n N_VPWR_c_1511_n 0.00776931f $X=1.835 $Y=3.72 $X2=0
+ $Y2=0
cc_442 N_A_37_107#_c_319_n N_VPWR_c_1511_n 0.0204951f $X=3.12 $Y=3.635 $X2=0
+ $Y2=0
cc_443 N_A_37_107#_c_360_p N_VPWR_c_1511_n 0.0182728f $X=3.82 $Y=3.6 $X2=0 $Y2=0
cc_444 N_A_37_107#_c_321_n N_VPWR_c_1511_n 0.0663306f $X=5.395 $Y=3.685 $X2=0
+ $Y2=0
cc_445 N_A_37_107#_c_324_n N_VPWR_c_1511_n 0.00655263f $X=3.905 $Y=3.685 $X2=0
+ $Y2=0
cc_446 N_A_37_107#_c_327_n N_VPWR_c_1511_n 0.0157316f $X=5.485 $Y=2.715 $X2=0
+ $Y2=0
cc_447 N_A_37_107#_c_381_p N_VPWR_c_1511_n 0.018265f $X=5.48 $Y=3.6 $X2=0 $Y2=0
cc_448 N_A_37_107#_c_330_n N_VPWR_c_1511_n 0.0135811f $X=6.865 $Y=2.96 $X2=0
+ $Y2=0
cc_449 N_A_37_107#_c_331_n N_VPWR_c_1511_n 0.0191126f $X=6.95 $Y=3.635 $X2=0
+ $Y2=0
cc_450 N_A_37_107#_c_332_n N_VPWR_c_1511_n 0.0304574f $X=7.565 $Y=3.72 $X2=0
+ $Y2=0
cc_451 N_A_37_107#_c_335_n N_VPWR_c_1511_n 0.00779018f $X=7.035 $Y=3.72 $X2=0
+ $Y2=0
cc_452 N_A_37_107#_c_338_n N_VPWR_c_1511_n 0.0194693f $X=7.65 $Y=3.635 $X2=0
+ $Y2=0
cc_453 N_A_37_107#_c_339_n N_VPWR_c_1511_n 0.0261168f $X=9.205 $Y=2.785 $X2=0
+ $Y2=0
cc_454 N_A_37_107#_c_296_n N_VPWR_c_1511_n 0.0173821f $X=9.29 $Y=1.985 $X2=0
+ $Y2=0
cc_455 N_A_37_107#_c_469_p N_VPWR_c_1511_n 0.00309396f $X=5.522 $Y=2.96 $X2=0
+ $Y2=0
cc_456 N_A_37_107#_c_313_n N_A_509_608#_c_1619_n 0.016277f $X=3.035 $Y=3.72
+ $X2=0 $Y2=0
cc_457 N_A_37_107#_c_319_n N_A_509_608#_c_1619_n 0.0408955f $X=3.12 $Y=3.635
+ $X2=0 $Y2=0
cc_458 N_A_37_107#_c_359_p N_A_509_608#_c_1619_n 0.0129587f $X=3.205 $Y=2.735
+ $X2=0 $Y2=0
cc_459 N_A_37_107#_c_320_n N_A_509_608#_c_1620_n 0.0487392f $X=3.735 $Y=2.735
+ $X2=0 $Y2=0
cc_460 N_A_37_107#_c_359_p N_A_509_608#_c_1620_n 0.0123662f $X=3.205 $Y=2.735
+ $X2=0 $Y2=0
cc_461 N_A_37_107#_M1006_g N_A_509_608#_c_1616_n 0.0100797f $X=4.88 $Y=1.075
+ $X2=0 $Y2=0
cc_462 N_A_37_107#_M1006_g N_A_509_608#_c_1617_n 0.0071608f $X=4.88 $Y=1.075
+ $X2=8.4 $Y2=0
cc_463 N_A_37_107#_c_320_n N_A_509_608#_c_1623_n 0.0066181f $X=3.735 $Y=2.735
+ $X2=8.4 $Y2=0.057
cc_464 N_A_37_107#_c_360_p N_A_509_608#_c_1623_n 0.00630942f $X=3.82 $Y=3.6
+ $X2=8.4 $Y2=0.057
cc_465 N_A_37_107#_c_360_p N_A_509_608#_c_1624_n 0.0292737f $X=3.82 $Y=3.6 $X2=0
+ $Y2=0
cc_466 N_A_37_107#_c_321_n N_A_509_608#_c_1624_n 0.0234562f $X=5.395 $Y=3.685
+ $X2=0 $Y2=0
cc_467 N_A_37_107#_M1006_g N_A_509_608#_c_1618_n 0.00526825f $X=4.88 $Y=1.075
+ $X2=0 $Y2=0
cc_468 N_A_37_107#_c_330_n A_1134_608# 0.00111857f $X=6.865 $Y=2.96 $X2=0 $Y2=0
cc_469 N_A_37_107#_M1003_g N_VGND_c_1722_n 0.0534923f $X=1.5 $Y=0.745 $X2=0
+ $Y2=0
cc_470 N_A_37_107#_c_291_n N_VGND_c_1722_n 0.0360269f $X=0.33 $Y=0.745 $X2=0
+ $Y2=0
cc_471 N_A_37_107#_M1003_g N_VGND_c_1724_n 0.00245457f $X=1.5 $Y=0.745 $X2=0
+ $Y2=0
cc_472 N_A_37_107#_M1003_g N_VGND_c_1734_n 0.00935388f $X=1.5 $Y=0.745 $X2=0
+ $Y2=0
cc_473 N_A_37_107#_c_291_n N_VGND_c_1734_n 0.0329542f $X=0.33 $Y=0.745 $X2=0
+ $Y2=0
cc_474 N_A_37_107#_c_297_n N_VGND_c_1734_n 0.00805752f $X=10.09 $Y=1.315 $X2=0
+ $Y2=0
cc_475 N_A_37_107#_c_383_p N_VGND_c_1734_n 0.00518526f $X=9.375 $Y=1.315 $X2=0
+ $Y2=0
cc_476 N_A_37_107#_c_384_p N_VGND_c_1734_n 0.00141706f $X=10.255 $Y=1.235 $X2=0
+ $Y2=0
cc_477 N_A_37_107#_M1005_g N_VGND_c_1734_n 0.00281472f $X=10.32 $Y=0.745 $X2=0
+ $Y2=0
cc_478 N_RESET_B_M1018_g N_D_c_752_n 0.05537f $X=3.08 $Y=3.25 $X2=0 $Y2=0
cc_479 N_RESET_B_c_554_n N_D_c_752_n 0.00112279f $X=3.58 $Y=1.505 $X2=0 $Y2=0
cc_480 N_RESET_B_c_570_n N_D_c_752_n 0.00165401f $X=3.39 $Y=1.645 $X2=0 $Y2=0
cc_481 N_RESET_B_M1018_g N_D_c_746_n 0.00433691f $X=3.08 $Y=3.25 $X2=0.24 $Y2=0
cc_482 N_RESET_B_c_570_n N_D_c_746_n 0.0378236f $X=3.39 $Y=1.645 $X2=0.24 $Y2=0
cc_483 N_RESET_B_c_552_n D 8.25959e-19 $X=3.39 $Y=1.395 $X2=0.24 $Y2=0
cc_484 N_RESET_B_c_554_n D 0.0790254f $X=3.58 $Y=1.505 $X2=0.24 $Y2=0
cc_485 N_RESET_B_c_555_n D 0.0214269f $X=6.455 $Y=0.545 $X2=0.24 $Y2=0
cc_486 N_RESET_B_c_570_n D 5.47031e-19 $X=3.39 $Y=1.645 $X2=0.24 $Y2=0
cc_487 N_RESET_B_c_552_n N_D_M1014_g 0.0378236f $X=3.39 $Y=1.395 $X2=16.56 $Y2=0
cc_488 N_RESET_B_c_554_n N_D_M1014_g 0.00914406f $X=3.58 $Y=1.505 $X2=16.56
+ $Y2=0
cc_489 N_RESET_B_c_555_n N_D_M1014_g 0.0172053f $X=6.455 $Y=0.545 $X2=16.56
+ $Y2=0
cc_490 N_RESET_B_c_611_p N_A_350_107#_c_796_n 0.00120637f $X=8.43 $Y=1.125
+ $X2=0.24 $Y2=0
cc_491 N_RESET_B_c_562_n N_A_350_107#_c_796_n 0.0224685f $X=10.905 $Y=0.35
+ $X2=0.24 $Y2=0
cc_492 N_RESET_B_M1018_g N_A_350_107#_c_799_n 0.0133646f $X=3.08 $Y=3.25 $X2=0
+ $Y2=0
cc_493 N_RESET_B_c_554_n N_A_350_107#_c_803_n 0.0440611f $X=3.58 $Y=1.505 $X2=0
+ $Y2=0
cc_494 N_RESET_B_c_570_n N_A_350_107#_c_803_n 0.00610993f $X=3.39 $Y=1.645 $X2=0
+ $Y2=0
cc_495 N_RESET_B_c_570_n N_A_350_107#_c_804_n 0.00222945f $X=3.39 $Y=1.645 $X2=0
+ $Y2=0
cc_496 N_RESET_B_c_560_n N_A_350_107#_c_805_n 0.0124639f $X=8.345 $Y=1.21 $X2=0
+ $Y2=0
cc_497 N_RESET_B_c_618_p N_A_350_107#_c_805_n 0.00102093f $X=6.625 $Y=1.21 $X2=0
+ $Y2=0
cc_498 N_RESET_B_c_561_n N_A_350_107#_c_805_n 0.0298798f $X=8.345 $Y=1.91 $X2=0
+ $Y2=0
cc_499 N_RESET_B_c_620_p N_A_350_107#_c_805_n 0.0185494f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_500 N_RESET_B_M1029_g N_A_350_107#_c_805_n 0.00584887f $X=7.265 $Y=1.075
+ $X2=0 $Y2=0
cc_501 N_RESET_B_c_570_n N_A_350_107#_c_806_n 0.0094077f $X=3.39 $Y=1.645 $X2=0
+ $Y2=0
cc_502 N_RESET_B_c_555_n N_A_350_107#_M1028_g 0.0162148f $X=6.455 $Y=0.545 $X2=0
+ $Y2=0
cc_503 N_RESET_B_c_559_n N_A_350_107#_M1028_g 0.00201786f $X=6.54 $Y=1.125 $X2=0
+ $Y2=0
cc_504 N_RESET_B_c_618_p N_A_350_107#_M1028_g 2.48855e-19 $X=6.625 $Y=1.21 $X2=0
+ $Y2=0
cc_505 N_RESET_B_c_570_n N_A_350_107#_c_812_n 0.0039277f $X=3.39 $Y=1.645 $X2=0
+ $Y2=0
cc_506 N_RESET_B_c_579_n N_A_1176_466#_c_987_n 0.0299234f $X=7.265 $Y=2.645
+ $X2=0 $Y2=0
cc_507 N_RESET_B_M1029_g N_A_1176_466#_c_987_n 0.00478065f $X=7.265 $Y=1.075
+ $X2=0 $Y2=0
cc_508 N_RESET_B_c_579_n N_A_1176_466#_M1022_g 0.0164991f $X=7.265 $Y=2.645
+ $X2=0 $Y2=0
cc_509 N_RESET_B_c_555_n N_A_1176_466#_M1031_g 0.00755369f $X=6.455 $Y=0.545
+ $X2=0 $Y2=0
cc_510 N_RESET_B_c_559_n N_A_1176_466#_M1031_g 0.0214101f $X=6.54 $Y=1.125 $X2=0
+ $Y2=0
cc_511 N_RESET_B_c_560_n N_A_1176_466#_M1031_g 0.00961899f $X=8.345 $Y=1.21
+ $X2=0 $Y2=0
cc_512 N_RESET_B_c_618_p N_A_1176_466#_M1031_g 0.00695687f $X=6.625 $Y=1.21
+ $X2=0 $Y2=0
cc_513 N_RESET_B_M1029_g N_A_1176_466#_M1031_g 0.0438714f $X=7.265 $Y=1.075
+ $X2=0 $Y2=0
cc_514 N_RESET_B_c_560_n N_A_1176_466#_c_984_n 5.6143e-19 $X=8.345 $Y=1.21 $X2=0
+ $Y2=0
cc_515 N_RESET_B_M1029_g N_A_1176_466#_c_984_n 0.0723084f $X=7.265 $Y=1.075
+ $X2=0 $Y2=0
cc_516 N_RESET_B_c_561_n N_A_1176_466#_c_1018_n 0.00700402f $X=8.345 $Y=1.91
+ $X2=0 $Y2=0
cc_517 N_RESET_B_M1029_g N_A_1176_466#_c_1018_n 0.00195494f $X=7.265 $Y=1.075
+ $X2=0 $Y2=0
cc_518 N_RESET_B_c_561_n N_A_1176_466#_c_985_n 5.10968e-19 $X=8.345 $Y=1.91
+ $X2=8.4 $Y2=0.057
cc_519 N_RESET_B_c_579_n N_A_1176_466#_c_991_n 0.00109361f $X=7.265 $Y=2.645
+ $X2=0 $Y2=0
cc_520 N_RESET_B_c_561_n N_A_1176_466#_c_991_n 0.0894381f $X=8.345 $Y=1.91 $X2=0
+ $Y2=0
cc_521 N_RESET_B_M1029_g N_A_1176_466#_c_991_n 0.032279f $X=7.265 $Y=1.075 $X2=0
+ $Y2=0
cc_522 N_RESET_B_c_561_n N_A_1176_466#_c_986_n 0.0128825f $X=8.345 $Y=1.91 $X2=0
+ $Y2=0
cc_523 N_RESET_B_c_611_p N_A_1176_466#_c_986_n 0.0346849f $X=8.43 $Y=1.125 $X2=0
+ $Y2=0
cc_524 N_RESET_B_c_620_p N_A_1176_466#_c_986_n 0.0350191f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_525 N_RESET_B_c_562_n N_A_1176_466#_c_986_n 0.0199321f $X=10.905 $Y=0.35
+ $X2=0 $Y2=0
cc_526 N_RESET_B_c_647_p N_A_1176_466#_c_986_n 0.0129587f $X=8.43 $Y=1.21 $X2=0
+ $Y2=0
cc_527 N_RESET_B_c_560_n N_A_978_608#_c_1073_n 0.0111401f $X=8.345 $Y=1.21
+ $X2=0.24 $Y2=0
cc_528 N_RESET_B_c_611_p N_A_978_608#_c_1073_n 0.0318677f $X=8.43 $Y=1.125
+ $X2=0.24 $Y2=0
cc_529 N_RESET_B_c_620_p N_A_978_608#_c_1073_n 0.00659601f $X=8.43 $Y=1.825
+ $X2=0.24 $Y2=0
cc_530 N_RESET_B_c_562_n N_A_978_608#_c_1073_n 0.00891555f $X=10.905 $Y=0.35
+ $X2=0.24 $Y2=0
cc_531 N_RESET_B_c_564_n N_A_978_608#_c_1073_n 0.00353941f $X=8.515 $Y=0.35
+ $X2=0.24 $Y2=0
cc_532 N_RESET_B_c_647_p N_A_978_608#_c_1073_n 0.00513124f $X=8.43 $Y=1.21
+ $X2=0.24 $Y2=0
cc_533 N_RESET_B_M1029_g N_A_978_608#_c_1073_n 0.0109138f $X=7.265 $Y=1.075
+ $X2=0.24 $Y2=0
cc_534 N_RESET_B_c_561_n N_A_978_608#_M1009_g 0.0104906f $X=8.345 $Y=1.91 $X2=0
+ $Y2=0
cc_535 N_RESET_B_M1029_g N_A_978_608#_M1009_g 0.0188667f $X=7.265 $Y=1.075 $X2=0
+ $Y2=0
cc_536 N_RESET_B_c_555_n N_A_978_608#_c_1075_n 0.0164585f $X=6.455 $Y=0.545
+ $X2=8.4 $Y2=0
cc_537 N_RESET_B_c_618_p N_A_978_608#_c_1075_n 0.00606097f $X=6.625 $Y=1.21
+ $X2=8.4 $Y2=0
cc_538 N_RESET_B_c_560_n N_A_978_608#_c_1078_n 0.0967999f $X=8.345 $Y=1.21 $X2=0
+ $Y2=0
cc_539 N_RESET_B_c_618_p N_A_978_608#_c_1078_n 0.0112593f $X=6.625 $Y=1.21 $X2=0
+ $Y2=0
cc_540 N_RESET_B_c_561_n N_A_978_608#_c_1078_n 0.0569956f $X=8.345 $Y=1.91 $X2=0
+ $Y2=0
cc_541 N_RESET_B_c_620_p N_A_978_608#_c_1078_n 0.0116761f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_542 N_RESET_B_M1029_g N_A_978_608#_c_1078_n 0.024145f $X=7.265 $Y=1.075 $X2=0
+ $Y2=0
cc_543 N_RESET_B_c_579_n N_A_978_608#_c_1087_n 0.0231935f $X=7.265 $Y=2.645
+ $X2=0 $Y2=0
cc_544 N_RESET_B_M1029_g N_A_978_608#_c_1087_n 0.0170584f $X=7.265 $Y=1.075
+ $X2=0 $Y2=0
cc_545 N_RESET_B_c_575_n N_A_978_608#_c_1088_n 0.00389904f $X=6.91 $Y=2.93 $X2=0
+ $Y2=0
cc_546 N_RESET_B_c_579_n N_A_978_608#_c_1088_n 0.0178638f $X=7.265 $Y=2.645
+ $X2=0 $Y2=0
cc_547 N_RESET_B_c_555_n N_A_978_608#_c_1079_n 0.0215139f $X=6.455 $Y=0.545
+ $X2=0 $Y2=0
cc_548 N_RESET_B_c_560_n N_A_978_608#_c_1081_n 0.0110232f $X=8.345 $Y=1.21 $X2=0
+ $Y2=0
cc_549 N_RESET_B_c_561_n N_A_978_608#_c_1081_n 0.0214908f $X=8.345 $Y=1.91 $X2=0
+ $Y2=0
cc_550 N_RESET_B_c_620_p N_A_978_608#_c_1081_n 0.0231276f $X=8.43 $Y=1.825 $X2=0
+ $Y2=0
cc_551 N_RESET_B_M1029_g N_A_978_608#_c_1081_n 0.0244647f $X=7.265 $Y=1.075
+ $X2=0 $Y2=0
cc_552 N_RESET_B_M1025_g N_A_2122_348#_c_1217_n 0.0567774f $X=11.74 $Y=2.52
+ $X2=0 $Y2=0
cc_553 N_RESET_B_M1025_g N_A_2122_348#_c_1218_n 0.0324759f $X=11.74 $Y=2.52
+ $X2=0 $Y2=0
cc_554 N_RESET_B_c_566_n N_A_2122_348#_c_1218_n 0.0101169f $X=11.51 $Y=1.045
+ $X2=0 $Y2=0
cc_555 N_RESET_B_c_567_n N_A_2122_348#_c_1218_n 0.0227892f $X=11.675 $Y=1.045
+ $X2=0 $Y2=0
cc_556 N_RESET_B_c_568_n N_A_2122_348#_c_1218_n 0.00348073f $X=11.675 $Y=1.25
+ $X2=0 $Y2=0
cc_557 N_RESET_B_c_568_n N_A_2122_348#_c_1219_n 0.00121827f $X=11.675 $Y=1.25
+ $X2=0 $Y2=0
cc_558 N_RESET_B_M1025_g N_A_2122_348#_c_1235_n 9.48226e-19 $X=11.74 $Y=2.52
+ $X2=0 $Y2=0
cc_559 N_RESET_B_c_566_n N_A_2122_348#_c_1235_n 0.0130351f $X=11.51 $Y=1.045
+ $X2=0 $Y2=0
cc_560 N_RESET_B_c_681_p N_A_2122_348#_c_1235_n 0.011388f $X=11.075 $Y=1.045
+ $X2=0 $Y2=0
cc_561 N_RESET_B_c_567_n N_A_2122_348#_c_1235_n 0.00220576f $X=11.675 $Y=1.045
+ $X2=0 $Y2=0
cc_562 N_RESET_B_c_568_n N_A_2122_348#_c_1235_n 0.00144299f $X=11.675 $Y=1.25
+ $X2=0 $Y2=0
cc_563 N_RESET_B_M1025_g N_A_2122_348#_c_1227_n 0.0127095f $X=11.74 $Y=2.52
+ $X2=0 $Y2=0
cc_564 N_RESET_B_c_571_n N_A_2122_348#_c_1220_n 0.00143997f $X=11.775 $Y=1.065
+ $X2=0 $Y2=0
cc_565 N_RESET_B_c_562_n N_A_2122_348#_M1007_g 0.00934051f $X=10.905 $Y=0.35
+ $X2=0 $Y2=0
cc_566 N_RESET_B_c_598_n N_A_2122_348#_M1007_g 0.0209646f $X=10.99 $Y=0.96 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_566_n N_A_2122_348#_M1007_g 0.0112453f $X=11.51 $Y=1.045
+ $X2=0 $Y2=0
cc_568 N_RESET_B_c_681_p N_A_2122_348#_M1007_g 0.0075568f $X=11.075 $Y=1.045
+ $X2=0 $Y2=0
cc_569 N_RESET_B_c_567_n N_A_2122_348#_M1007_g 0.00154335f $X=11.675 $Y=1.045
+ $X2=0 $Y2=0
cc_570 N_RESET_B_c_568_n N_A_2122_348#_M1007_g 0.0405493f $X=11.675 $Y=1.25
+ $X2=0 $Y2=0
cc_571 N_RESET_B_c_571_n N_A_2122_348#_M1007_g 0.0157013f $X=11.775 $Y=1.065
+ $X2=0 $Y2=0
cc_572 N_RESET_B_M1025_g N_A_1900_107#_M1001_g 0.0102357f $X=11.74 $Y=2.52 $X2=0
+ $Y2=0
cc_573 N_RESET_B_c_567_n N_A_1900_107#_M1001_g 0.00182015f $X=11.675 $Y=1.045
+ $X2=0 $Y2=0
cc_574 N_RESET_B_c_571_n N_A_1900_107#_M1001_g 0.0806803f $X=11.775 $Y=1.065
+ $X2=0 $Y2=0
cc_575 N_RESET_B_M1025_g N_A_1900_107#_c_1305_n 0.0155799f $X=11.74 $Y=2.52
+ $X2=0.24 $Y2=0
cc_576 N_RESET_B_c_562_n N_A_1900_107#_c_1326_n 0.0103975f $X=10.905 $Y=0.35
+ $X2=0 $Y2=0
cc_577 N_RESET_B_c_598_n N_A_1900_107#_c_1326_n 0.00568401f $X=10.99 $Y=0.96
+ $X2=0 $Y2=0
cc_578 N_RESET_B_c_598_n N_A_1900_107#_c_1302_n 0.00577724f $X=10.99 $Y=0.96
+ $X2=0 $Y2=0
cc_579 N_RESET_B_c_681_p N_A_1900_107#_c_1302_n 0.0128864f $X=11.075 $Y=1.045
+ $X2=0 $Y2=0
cc_580 N_RESET_B_M1025_g N_A_1900_107#_c_1319_n 0.0401969f $X=11.74 $Y=2.52
+ $X2=0 $Y2=0
cc_581 N_RESET_B_c_562_n N_A_1900_107#_c_1303_n 0.0609551f $X=10.905 $Y=0.35
+ $X2=0 $Y2=0
cc_582 N_RESET_B_M1025_g N_A_1900_107#_c_1345_n 0.00100296f $X=11.74 $Y=2.52
+ $X2=0 $Y2=0
cc_583 N_RESET_B_M1025_g N_A_1900_107#_c_1304_n 0.0342216f $X=11.74 $Y=2.52
+ $X2=0 $Y2=0
cc_584 N_RESET_B_M1018_g N_VPWR_c_1493_n 0.00136844f $X=3.08 $Y=3.25 $X2=0 $Y2=0
cc_585 N_RESET_B_c_575_n N_VPWR_c_1496_n 0.00755674f $X=6.91 $Y=2.93 $X2=0 $Y2=0
cc_586 N_RESET_B_M1025_g N_VPWR_c_1502_n 0.0264777f $X=11.74 $Y=2.52 $X2=0 $Y2=0
cc_587 N_RESET_B_M1018_g N_VPWR_c_1511_n 0.0216125f $X=3.08 $Y=3.25 $X2=0 $Y2=0
cc_588 N_RESET_B_c_575_n N_VPWR_c_1511_n 0.013947f $X=6.91 $Y=2.93 $X2=0 $Y2=0
cc_589 N_RESET_B_M1025_g N_VPWR_c_1511_n 0.0111527f $X=11.74 $Y=2.52 $X2=0 $Y2=0
cc_590 N_RESET_B_c_579_n N_VPWR_c_1511_n 0.00479281f $X=7.265 $Y=2.645 $X2=0
+ $Y2=0
cc_591 N_RESET_B_M1018_g N_A_509_608#_c_1619_n 0.0332857f $X=3.08 $Y=3.25 $X2=0
+ $Y2=0
cc_592 N_RESET_B_M1018_g N_A_509_608#_c_1620_n 0.0293885f $X=3.08 $Y=3.25 $X2=0
+ $Y2=0
cc_593 N_RESET_B_c_554_n N_A_509_608#_c_1620_n 0.0502318f $X=3.58 $Y=1.505 $X2=0
+ $Y2=0
cc_594 N_RESET_B_c_570_n N_A_509_608#_c_1620_n 0.00118209f $X=3.39 $Y=1.645
+ $X2=0 $Y2=0
cc_595 N_RESET_B_M1018_g N_A_509_608#_c_1621_n 0.0045224f $X=3.08 $Y=3.25 $X2=0
+ $Y2=0
cc_596 N_RESET_B_c_555_n N_A_509_608#_c_1616_n 0.0204346f $X=6.455 $Y=0.545
+ $X2=0 $Y2=0
cc_597 N_RESET_B_c_560_n N_VGND_M1029_d 0.00933647f $X=8.345 $Y=1.21 $X2=0 $Y2=0
cc_598 N_RESET_B_c_552_n N_VGND_c_1724_n 0.0292763f $X=3.39 $Y=1.395 $X2=0 $Y2=0
cc_599 N_RESET_B_c_554_n N_VGND_c_1724_n 0.07623f $X=3.58 $Y=1.505 $X2=0 $Y2=0
cc_600 N_RESET_B_c_557_n N_VGND_c_1724_n 0.0119967f $X=3.665 $Y=0.545 $X2=0
+ $Y2=0
cc_601 N_RESET_B_c_570_n N_VGND_c_1724_n 0.0130403f $X=3.39 $Y=1.645 $X2=0 $Y2=0
cc_602 N_RESET_B_c_555_n N_VGND_c_1726_n 0.00325109f $X=6.455 $Y=0.545 $X2=0
+ $Y2=0
cc_603 N_RESET_B_c_559_n N_VGND_c_1726_n 0.00938421f $X=6.54 $Y=1.125 $X2=0
+ $Y2=0
cc_604 N_RESET_B_c_560_n N_VGND_c_1726_n 0.0642307f $X=8.345 $Y=1.21 $X2=0 $Y2=0
cc_605 N_RESET_B_c_611_p N_VGND_c_1726_n 0.0212201f $X=8.43 $Y=1.125 $X2=0 $Y2=0
cc_606 N_RESET_B_c_564_n N_VGND_c_1726_n 0.00473621f $X=8.515 $Y=0.35 $X2=0
+ $Y2=0
cc_607 N_RESET_B_M1029_g N_VGND_c_1726_n 0.02468f $X=7.265 $Y=1.075 $X2=0 $Y2=0
cc_608 N_RESET_B_c_562_n N_VGND_c_1728_n 0.00461601f $X=10.905 $Y=0.35 $X2=0
+ $Y2=0
cc_609 N_RESET_B_c_598_n N_VGND_c_1728_n 0.022881f $X=10.99 $Y=0.96 $X2=0 $Y2=0
cc_610 N_RESET_B_c_566_n N_VGND_c_1728_n 0.0153548f $X=11.51 $Y=1.045 $X2=0
+ $Y2=0
cc_611 N_RESET_B_c_567_n N_VGND_c_1728_n 0.0210012f $X=11.675 $Y=1.045 $X2=0
+ $Y2=0
cc_612 N_RESET_B_c_571_n N_VGND_c_1728_n 0.0434618f $X=11.775 $Y=1.065 $X2=0
+ $Y2=0
cc_613 N_RESET_B_c_552_n N_VGND_c_1734_n 0.00593019f $X=3.39 $Y=1.395 $X2=0
+ $Y2=0
cc_614 N_RESET_B_c_555_n N_VGND_c_1734_n 0.159696f $X=6.455 $Y=0.545 $X2=0 $Y2=0
cc_615 N_RESET_B_c_557_n N_VGND_c_1734_n 0.0127114f $X=3.665 $Y=0.545 $X2=0
+ $Y2=0
cc_616 N_RESET_B_c_560_n N_VGND_c_1734_n 0.0294584f $X=8.345 $Y=1.21 $X2=0 $Y2=0
cc_617 N_RESET_B_c_611_p N_VGND_c_1734_n 0.0199533f $X=8.43 $Y=1.125 $X2=0 $Y2=0
cc_618 N_RESET_B_c_562_n N_VGND_c_1734_n 0.089453f $X=10.905 $Y=0.35 $X2=0 $Y2=0
cc_619 N_RESET_B_c_564_n N_VGND_c_1734_n 0.00776561f $X=8.515 $Y=0.35 $X2=0
+ $Y2=0
cc_620 N_RESET_B_c_598_n N_VGND_c_1734_n 0.019173f $X=10.99 $Y=0.96 $X2=0 $Y2=0
cc_621 N_RESET_B_c_566_n N_VGND_c_1734_n 0.0076026f $X=11.51 $Y=1.045 $X2=0
+ $Y2=0
cc_622 N_RESET_B_c_567_n N_VGND_c_1734_n 0.00169922f $X=11.675 $Y=1.045 $X2=0
+ $Y2=0
cc_623 N_RESET_B_M1029_g N_VGND_c_1734_n 0.0065328f $X=7.265 $Y=1.075 $X2=0
+ $Y2=0
cc_624 N_RESET_B_c_560_n A_1357_173# 0.00213952f $X=8.345 $Y=1.21 $X2=0 $Y2=0
cc_625 N_D_M1008_g N_A_350_107#_c_816_n 0.0265195f $X=3.86 $Y=3.25 $X2=0 $Y2=0
cc_626 N_D_c_751_n N_A_350_107#_c_816_n 0.0329278f $X=3.895 $Y=2.135 $X2=0 $Y2=0
cc_627 N_D_M1014_g N_A_350_107#_c_843_n 3.1021e-19 $X=4.1 $Y=1.075 $X2=0 $Y2=0
cc_628 N_D_c_752_n N_A_350_107#_c_803_n 0.00450193f $X=3.895 $Y=2.635 $X2=0
+ $Y2=0
cc_629 N_D_c_746_n N_A_350_107#_c_803_n 0.00263833f $X=4.1 $Y=1.915 $X2=0 $Y2=0
cc_630 D N_A_350_107#_c_803_n 0.0302969f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_631 N_D_M1014_g N_A_350_107#_c_803_n 0.00782181f $X=4.1 $Y=1.075 $X2=0 $Y2=0
cc_632 N_D_M1008_g N_VPWR_c_1493_n 0.00136844f $X=3.86 $Y=3.25 $X2=0 $Y2=0
cc_633 N_D_M1008_g N_VPWR_c_1511_n 0.0199373f $X=3.86 $Y=3.25 $X2=0 $Y2=0
cc_634 N_D_c_752_n N_A_509_608#_c_1620_n 0.0358096f $X=3.895 $Y=2.635 $X2=0
+ $Y2=0
cc_635 N_D_c_746_n N_A_509_608#_c_1620_n 0.00543882f $X=4.1 $Y=1.915 $X2=0 $Y2=0
cc_636 D N_A_509_608#_c_1620_n 0.0205917f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_637 D N_A_509_608#_c_1616_n 0.088204f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_638 N_D_M1014_g N_A_509_608#_c_1616_n 0.00573446f $X=4.1 $Y=1.075 $X2=0 $Y2=0
cc_639 N_D_c_751_n N_A_509_608#_c_1617_n 0.00877159f $X=3.895 $Y=2.135 $X2=8.4
+ $Y2=0
cc_640 N_D_c_746_n N_A_509_608#_c_1617_n 0.00513274f $X=4.1 $Y=1.915 $X2=8.4
+ $Y2=0
cc_641 N_D_M1014_g N_A_509_608#_c_1617_n 0.00709523f $X=4.1 $Y=1.075 $X2=8.4
+ $Y2=0
cc_642 N_D_M1008_g N_A_509_608#_c_1623_n 0.00323081f $X=3.86 $Y=3.25 $X2=8.4
+ $Y2=0.057
cc_643 N_D_c_752_n N_A_509_608#_c_1623_n 0.0034404f $X=3.895 $Y=2.635 $X2=8.4
+ $Y2=0.057
cc_644 N_D_M1008_g N_A_509_608#_c_1624_n 0.00855431f $X=3.86 $Y=3.25 $X2=0 $Y2=0
cc_645 N_D_c_752_n N_A_509_608#_c_1624_n 0.00173516f $X=3.895 $Y=2.635 $X2=0
+ $Y2=0
cc_646 N_D_M1014_g N_A_509_608#_c_1618_n 0.00294597f $X=4.1 $Y=1.075 $X2=0 $Y2=0
cc_647 D N_VGND_c_1734_n 0.00242412f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_648 N_A_350_107#_c_805_n N_A_1176_466#_c_987_n 2.4715e-19 $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_649 N_A_350_107#_M1028_g N_A_1176_466#_c_987_n 0.0128285f $X=5.825 $Y=1.075
+ $X2=0 $Y2=0
cc_650 N_A_350_107#_M1028_g N_A_1176_466#_M1031_g 0.0920651f $X=5.825 $Y=1.075
+ $X2=0 $Y2=0
cc_651 N_A_350_107#_c_844_n N_A_1176_466#_c_984_n 2.89102e-19 $X=5.76 $Y=1.595
+ $X2=0 $Y2=0
cc_652 N_A_350_107#_c_805_n N_A_1176_466#_c_984_n 3.0408e-19 $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_653 N_A_350_107#_c_805_n N_A_1176_466#_c_1018_n 0.00799912f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_654 N_A_350_107#_c_805_n N_A_1176_466#_c_985_n 0.0105968f $X=9.695 $Y=1.665
+ $X2=8.4 $Y2=0.057
cc_655 N_A_350_107#_c_805_n N_A_1176_466#_c_991_n 0.0154939f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_656 N_A_350_107#_c_796_n N_A_1176_466#_c_986_n 0.0257611f $X=9.25 $Y=1.395
+ $X2=0 $Y2=0
cc_657 N_A_350_107#_c_798_n N_A_1176_466#_c_986_n 0.00582222f $X=9.5 $Y=1.492
+ $X2=0 $Y2=0
cc_658 N_A_350_107#_c_805_n N_A_1176_466#_c_986_n 0.041779f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_659 N_A_350_107#_c_796_n N_A_978_608#_c_1073_n 0.0118378f $X=9.25 $Y=1.395
+ $X2=0.24 $Y2=0
cc_660 N_A_350_107#_c_844_n N_A_978_608#_c_1084_n 0.0234651f $X=5.76 $Y=1.595
+ $X2=0 $Y2=0
cc_661 N_A_350_107#_c_802_n N_A_978_608#_c_1084_n 0.0120811f $X=5.595 $Y=1.642
+ $X2=0 $Y2=0
cc_662 N_A_350_107#_c_805_n N_A_978_608#_c_1084_n 0.00933264f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_663 N_A_350_107#_M1028_g N_A_978_608#_c_1084_n 0.0109485f $X=5.825 $Y=1.075
+ $X2=0 $Y2=0
cc_664 N_A_350_107#_c_815_n N_A_978_608#_c_1085_n 0.0131382f $X=4.78 $Y=2.315
+ $X2=0 $Y2=0
cc_665 N_A_350_107#_c_816_n N_A_978_608#_c_1085_n 0.00135507f $X=4.78 $Y=2.315
+ $X2=0 $Y2=0
cc_666 N_A_350_107#_c_802_n N_A_978_608#_c_1085_n 0.00450453f $X=5.595 $Y=1.642
+ $X2=0 $Y2=0
cc_667 N_A_350_107#_c_851_n N_A_978_608#_c_1085_n 0.00295568f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_668 N_A_350_107#_c_844_n N_A_978_608#_c_1075_n 0.0212997f $X=5.76 $Y=1.595
+ $X2=8.4 $Y2=0
cc_669 N_A_350_107#_c_805_n N_A_978_608#_c_1075_n 0.00816987f $X=9.695 $Y=1.665
+ $X2=8.4 $Y2=0
cc_670 N_A_350_107#_M1028_g N_A_978_608#_c_1075_n 0.0266026f $X=5.825 $Y=1.075
+ $X2=8.4 $Y2=0
cc_671 N_A_350_107#_M1028_g N_A_978_608#_c_1076_n 0.00366742f $X=5.825 $Y=1.075
+ $X2=0 $Y2=0
cc_672 N_A_350_107#_c_844_n N_A_978_608#_c_1077_n 0.0262336f $X=5.76 $Y=1.595
+ $X2=0 $Y2=0
cc_673 N_A_350_107#_c_805_n N_A_978_608#_c_1077_n 0.0105865f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_674 N_A_350_107#_M1028_g N_A_978_608#_c_1077_n 0.00518844f $X=5.825 $Y=1.075
+ $X2=0 $Y2=0
cc_675 N_A_350_107#_c_805_n N_A_978_608#_c_1078_n 0.0547824f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_676 N_A_350_107#_M1030_g N_A_978_608#_c_1089_n 0.0117121f $X=4.64 $Y=3.25
+ $X2=0 $Y2=0
cc_677 N_A_350_107#_c_816_n N_A_978_608#_c_1089_n 0.00348119f $X=4.78 $Y=2.315
+ $X2=0 $Y2=0
cc_678 N_A_350_107#_M1030_g N_A_978_608#_c_1090_n 9.45538e-19 $X=4.64 $Y=3.25
+ $X2=0 $Y2=0
cc_679 N_A_350_107#_c_815_n N_A_978_608#_c_1090_n 0.030793f $X=4.78 $Y=2.315
+ $X2=0 $Y2=0
cc_680 N_A_350_107#_c_816_n N_A_978_608#_c_1090_n 0.00409847f $X=4.78 $Y=2.315
+ $X2=0 $Y2=0
cc_681 N_A_350_107#_c_802_n N_A_978_608#_c_1079_n 0.0236956f $X=5.595 $Y=1.642
+ $X2=0 $Y2=0
cc_682 N_A_350_107#_c_805_n N_A_978_608#_c_1079_n 0.00218096f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_683 N_A_350_107#_M1028_g N_A_978_608#_c_1079_n 0.0109118f $X=5.825 $Y=1.075
+ $X2=0 $Y2=0
cc_684 N_A_350_107#_c_844_n N_A_978_608#_c_1080_n 0.0105589f $X=5.76 $Y=1.595
+ $X2=0 $Y2=0
cc_685 N_A_350_107#_c_805_n N_A_978_608#_c_1080_n 0.00973981f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_686 N_A_350_107#_M1028_g N_A_978_608#_c_1080_n 0.00210817f $X=5.825 $Y=1.075
+ $X2=0 $Y2=0
cc_687 N_A_350_107#_c_798_n N_A_978_608#_c_1081_n 0.0118378f $X=9.5 $Y=1.492
+ $X2=0 $Y2=0
cc_688 N_A_350_107#_c_805_n N_A_978_608#_c_1081_n 0.0161474f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_689 N_A_350_107#_c_808_n N_A_2122_348#_c_1217_n 2.38523e-19 $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_690 N_A_350_107#_c_810_n N_A_2122_348#_c_1217_n 0.0354737f $X=9.895 $Y=1.925
+ $X2=0 $Y2=0
cc_691 N_A_350_107#_c_819_n N_A_2122_348#_c_1217_n 0.0354737f $X=10.052 $Y=2.2
+ $X2=0 $Y2=0
cc_692 N_A_350_107#_c_797_n N_A_1900_107#_c_1314_n 0.00378462f $X=9.71 $Y=1.492
+ $X2=0 $Y2=0
cc_693 N_A_350_107#_c_805_n N_A_1900_107#_c_1314_n 0.005196f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_694 N_A_350_107#_c_807_n N_A_1900_107#_c_1314_n 0.00155292f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_695 N_A_350_107#_c_808_n N_A_1900_107#_c_1314_n 0.00631227f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_696 N_A_350_107#_c_810_n N_A_1900_107#_c_1314_n 0.00330429f $X=9.895 $Y=1.925
+ $X2=0 $Y2=0
cc_697 N_A_350_107#_c_819_n N_A_1900_107#_c_1315_n 0.0115771f $X=10.052 $Y=2.2
+ $X2=0 $Y2=0
cc_698 N_A_350_107#_c_807_n N_A_1900_107#_c_1317_n 6.82026e-19 $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_699 N_A_350_107#_c_808_n N_A_1900_107#_c_1317_n 0.0178269f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_700 N_A_350_107#_c_810_n N_A_1900_107#_c_1317_n 0.00258485f $X=9.895 $Y=1.925
+ $X2=0 $Y2=0
cc_701 N_A_350_107#_c_819_n N_A_1900_107#_c_1317_n 0.0317034f $X=10.052 $Y=2.2
+ $X2=0 $Y2=0
cc_702 N_A_350_107#_c_797_n N_A_1900_107#_c_1302_n 0.00202798f $X=9.71 $Y=1.492
+ $X2=0 $Y2=0
cc_703 N_A_350_107#_c_807_n N_A_1900_107#_c_1302_n 0.00215053f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_704 N_A_350_107#_c_808_n N_A_1900_107#_c_1302_n 0.0134639f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_705 N_A_350_107#_c_810_n N_A_1900_107#_c_1302_n 0.00246641f $X=9.895 $Y=1.925
+ $X2=0 $Y2=0
cc_706 N_A_350_107#_c_808_n N_A_1900_107#_c_1320_n 0.00686795f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_707 N_A_350_107#_c_810_n N_A_1900_107#_c_1320_n 0.0140448f $X=9.895 $Y=1.925
+ $X2=0 $Y2=0
cc_708 N_A_350_107#_c_819_n N_A_1900_107#_c_1320_n 0.0138037f $X=10.052 $Y=2.2
+ $X2=0 $Y2=0
cc_709 N_A_350_107#_c_796_n N_A_1900_107#_c_1303_n 0.00705752f $X=9.25 $Y=1.395
+ $X2=0 $Y2=0
cc_710 N_A_350_107#_c_797_n N_A_1900_107#_c_1303_n 0.00140822f $X=9.71 $Y=1.492
+ $X2=0 $Y2=0
cc_711 N_A_350_107#_c_819_n N_VPWR_c_1502_n 0.00441791f $X=10.052 $Y=2.2 $X2=0
+ $Y2=0
cc_712 N_A_350_107#_M1030_g N_VPWR_c_1511_n 0.0259948f $X=4.64 $Y=3.25 $X2=0
+ $Y2=0
cc_713 N_A_350_107#_c_799_n N_VPWR_c_1511_n 0.0183374f $X=2.1 $Y=2.79 $X2=0
+ $Y2=0
cc_714 N_A_350_107#_c_819_n N_VPWR_c_1511_n 0.0123644f $X=10.052 $Y=2.2 $X2=0
+ $Y2=0
cc_715 N_A_350_107#_c_799_n N_A_509_608#_c_1619_n 0.0593634f $X=2.1 $Y=2.79
+ $X2=0 $Y2=0
cc_716 N_A_350_107#_c_803_n N_A_509_608#_c_1620_n 0.0165907f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_717 N_A_350_107#_c_799_n N_A_509_608#_c_1621_n 0.0112865f $X=2.1 $Y=2.79
+ $X2=0 $Y2=0
cc_718 N_A_350_107#_c_803_n N_A_509_608#_c_1621_n 0.0117795f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_719 N_A_350_107#_c_815_n N_A_509_608#_c_1617_n 0.0357411f $X=4.78 $Y=2.315
+ $X2=8.4 $Y2=0
cc_720 N_A_350_107#_c_816_n N_A_509_608#_c_1617_n 0.00785165f $X=4.78 $Y=2.315
+ $X2=8.4 $Y2=0
cc_721 N_A_350_107#_c_843_n N_A_509_608#_c_1617_n 0.018971f $X=4.865 $Y=1.642
+ $X2=8.4 $Y2=0
cc_722 N_A_350_107#_c_803_n N_A_509_608#_c_1617_n 0.0202049f $X=4.895 $Y=1.665
+ $X2=8.4 $Y2=0
cc_723 N_A_350_107#_c_851_n N_A_509_608#_c_1617_n 4.2434e-19 $X=5.185 $Y=1.665
+ $X2=8.4 $Y2=0
cc_724 N_A_350_107#_M1030_g N_A_509_608#_c_1623_n 0.00402436f $X=4.64 $Y=3.25
+ $X2=8.4 $Y2=0.057
cc_725 N_A_350_107#_c_815_n N_A_509_608#_c_1623_n 0.0226279f $X=4.78 $Y=2.315
+ $X2=8.4 $Y2=0.057
cc_726 N_A_350_107#_c_816_n N_A_509_608#_c_1623_n 0.013469f $X=4.78 $Y=2.315
+ $X2=8.4 $Y2=0.057
cc_727 N_A_350_107#_M1030_g N_A_509_608#_c_1624_n 0.0155308f $X=4.64 $Y=3.25
+ $X2=0 $Y2=0
cc_728 N_A_350_107#_c_803_n N_A_509_608#_c_1618_n 0.00622714f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_729 N_A_350_107#_c_815_n N_A_509_608#_c_1670_n 0.0123662f $X=4.78 $Y=2.315
+ $X2=0 $Y2=0
cc_730 N_A_350_107#_c_816_n N_A_509_608#_c_1670_n 0.00602522f $X=4.78 $Y=2.315
+ $X2=0 $Y2=0
cc_731 N_A_350_107#_c_800_n N_VGND_c_1722_n 0.0232694f $X=2.1 $Y=0.745 $X2=0
+ $Y2=0
cc_732 N_A_350_107#_c_800_n N_VGND_c_1724_n 0.0406247f $X=2.1 $Y=0.745 $X2=0
+ $Y2=0
cc_733 N_A_350_107#_c_803_n N_VGND_c_1724_n 0.0309883f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_734 N_A_350_107#_c_812_n N_VGND_c_1724_n 0.02666f $X=2.145 $Y=1.55 $X2=0
+ $Y2=0
cc_735 N_A_350_107#_M1003_d N_VGND_c_1734_n 0.00221032f $X=1.75 $Y=0.535 $X2=0
+ $Y2=0
cc_736 N_A_350_107#_c_796_n N_VGND_c_1734_n 0.0170573f $X=9.25 $Y=1.395 $X2=0
+ $Y2=0
cc_737 N_A_350_107#_c_800_n N_VGND_c_1734_n 0.0276225f $X=2.1 $Y=0.745 $X2=0
+ $Y2=0
cc_738 N_A_350_107#_c_812_n N_VGND_c_1734_n 4.53502e-19 $X=2.145 $Y=1.55 $X2=0
+ $Y2=0
cc_739 N_A_1176_466#_c_986_n N_A_978_608#_c_1073_n 0.0152055f $X=8.86 $Y=0.7
+ $X2=0.24 $Y2=0
cc_740 N_A_1176_466#_c_991_n N_A_978_608#_M1009_g 0.0291241f $X=8.695 $Y=2.26
+ $X2=0 $Y2=0
cc_741 N_A_1176_466#_c_986_n N_A_978_608#_M1009_g 0.013369f $X=8.86 $Y=0.7 $X2=0
+ $Y2=0
cc_742 N_A_1176_466#_c_1006_n N_A_978_608#_M1009_g 0.0111093f $X=8.86 $Y=2.26
+ $X2=0 $Y2=0
cc_743 N_A_1176_466#_c_987_n N_A_978_608#_c_1084_n 0.00860495f $X=6.13 $Y=2.91
+ $X2=0 $Y2=0
cc_744 N_A_1176_466#_M1031_g N_A_978_608#_c_1075_n 0.00169455f $X=6.535 $Y=1.075
+ $X2=8.4 $Y2=0
cc_745 N_A_1176_466#_M1031_g N_A_978_608#_c_1076_n 0.00376182f $X=6.535 $Y=1.075
+ $X2=0 $Y2=0
cc_746 N_A_1176_466#_c_984_n N_A_978_608#_c_1077_n 0.00897168f $X=6.545 $Y=1.675
+ $X2=0 $Y2=0
cc_747 N_A_1176_466#_c_1018_n N_A_978_608#_c_1077_n 0.0251553f $X=6.62 $Y=1.91
+ $X2=0 $Y2=0
cc_748 N_A_1176_466#_c_1049_p N_A_978_608#_c_1077_n 0.00187626f $X=6.785 $Y=2.26
+ $X2=0 $Y2=0
cc_749 N_A_1176_466#_c_987_n N_A_978_608#_c_1102_n 0.0118821f $X=6.13 $Y=2.91
+ $X2=0 $Y2=0
cc_750 N_A_1176_466#_c_984_n N_A_978_608#_c_1078_n 0.0302172f $X=6.545 $Y=1.675
+ $X2=0 $Y2=0
cc_751 N_A_1176_466#_c_1018_n N_A_978_608#_c_1078_n 0.0197788f $X=6.62 $Y=1.91
+ $X2=0 $Y2=0
cc_752 N_A_1176_466#_c_991_n N_A_978_608#_c_1078_n 0.00653266f $X=8.695 $Y=2.26
+ $X2=0 $Y2=0
cc_753 N_A_1176_466#_c_987_n N_A_978_608#_c_1087_n 0.0227888f $X=6.13 $Y=2.91
+ $X2=0 $Y2=0
cc_754 N_A_1176_466#_c_991_n N_A_978_608#_c_1087_n 0.0418079f $X=8.695 $Y=2.26
+ $X2=0 $Y2=0
cc_755 N_A_1176_466#_c_1049_p N_A_978_608#_c_1087_n 0.0247192f $X=6.785 $Y=2.26
+ $X2=0 $Y2=0
cc_756 N_A_1176_466#_c_987_n N_A_978_608#_c_1104_n 0.00804903f $X=6.13 $Y=2.91
+ $X2=0 $Y2=0
cc_757 N_A_1176_466#_c_987_n N_A_978_608#_c_1090_n 7.41631e-19 $X=6.13 $Y=2.91
+ $X2=0 $Y2=0
cc_758 N_A_1176_466#_M1031_g N_A_978_608#_c_1079_n 0.00101042f $X=6.535 $Y=1.075
+ $X2=0 $Y2=0
cc_759 N_A_1176_466#_c_987_n N_A_978_608#_c_1091_n 0.00634819f $X=6.13 $Y=2.91
+ $X2=0 $Y2=0
cc_760 N_A_1176_466#_c_985_n N_A_978_608#_c_1091_n 0.00403169f $X=6.62 $Y=1.91
+ $X2=0 $Y2=0
cc_761 N_A_1176_466#_c_1049_p N_A_978_608#_c_1091_n 0.0122668f $X=6.785 $Y=2.26
+ $X2=0 $Y2=0
cc_762 N_A_1176_466#_c_991_n N_A_978_608#_c_1081_n 0.00218303f $X=8.695 $Y=2.26
+ $X2=0 $Y2=0
cc_763 N_A_1176_466#_c_986_n N_A_978_608#_c_1081_n 0.0151782f $X=8.86 $Y=0.7
+ $X2=0 $Y2=0
cc_764 N_A_1176_466#_c_986_n N_A_1900_107#_c_1303_n 0.0117897f $X=8.86 $Y=0.7
+ $X2=0 $Y2=0
cc_765 N_A_1176_466#_c_991_n N_VPWR_M1009_s 0.00363461f $X=8.695 $Y=2.26 $X2=0
+ $Y2=0
cc_766 N_A_1176_466#_c_987_n N_VPWR_c_1496_n 2.53921e-19 $X=6.13 $Y=2.91 $X2=0
+ $Y2=0
cc_767 N_A_1176_466#_M1022_g N_VPWR_c_1496_n 0.036216f $X=6.13 $Y=3.25 $X2=0
+ $Y2=0
cc_768 N_A_1176_466#_M1009_d N_VPWR_c_1499_n 0.00447727f $X=8.72 $Y=2.31 $X2=0
+ $Y2=0
cc_769 N_A_1176_466#_M1031_g N_VGND_c_1726_n 6.39957e-19 $X=6.535 $Y=1.075 $X2=0
+ $Y2=0
cc_770 N_A_1176_466#_M1031_g N_VGND_c_1734_n 0.00526225f $X=6.535 $Y=1.075 $X2=0
+ $Y2=0
cc_771 N_A_1176_466#_c_986_n N_VGND_c_1734_n 0.022856f $X=8.86 $Y=0.7 $X2=0
+ $Y2=0
cc_772 N_A_978_608#_M1009_g N_VPWR_c_1499_n 0.040998f $X=8.47 $Y=2.81 $X2=0
+ $Y2=0
cc_773 N_A_978_608#_M1030_d N_VPWR_c_1511_n 0.0021813f $X=4.89 $Y=3.04 $X2=0
+ $Y2=0
cc_774 N_A_978_608#_M1011_d N_VPWR_c_1511_n 0.002211f $X=7.16 $Y=3.04 $X2=0
+ $Y2=0
cc_775 N_A_978_608#_c_1088_n N_VPWR_c_1511_n 0.00724238f $X=7.3 $Y=3.225 $X2=0
+ $Y2=0
cc_776 N_A_978_608#_c_1089_n N_VPWR_c_1511_n 0.0122393f $X=5.03 $Y=3.25 $X2=0
+ $Y2=0
cc_777 N_A_978_608#_c_1079_n N_A_509_608#_c_1616_n 0.014111f $X=5.435 $Y=1.075
+ $X2=0 $Y2=0
cc_778 N_A_978_608#_c_1090_n N_A_509_608#_c_1623_n 0.00542521f $X=5.04 $Y=3
+ $X2=8.4 $Y2=0.057
cc_779 N_A_978_608#_c_1089_n N_A_509_608#_c_1624_n 0.0180684f $X=5.03 $Y=3.25
+ $X2=0 $Y2=0
cc_780 N_A_978_608#_c_1073_n N_VGND_c_1726_n 0.00995687f $X=8.47 $Y=1.395 $X2=0
+ $Y2=0
cc_781 N_A_978_608#_c_1073_n N_VGND_c_1734_n 0.0156107f $X=8.47 $Y=1.395 $X2=0
+ $Y2=0
cc_782 N_A_978_608#_c_1075_n N_VGND_c_1734_n 0.00408437f $X=6.105 $Y=1.24 $X2=0
+ $Y2=0
cc_783 N_A_978_608#_c_1079_n N_VGND_c_1734_n 0.00261152f $X=5.435 $Y=1.075 $X2=0
+ $Y2=0
cc_784 N_A_978_608#_c_1075_n A_1215_173# 0.0017778f $X=6.105 $Y=1.24 $X2=0 $Y2=0
cc_785 N_A_2122_348#_c_1218_n N_A_1900_107#_M1001_g 0.0222378f $X=12.71 $Y=1.615
+ $X2=0 $Y2=0
cc_786 N_A_2122_348#_c_1219_n N_A_1900_107#_M1001_g 0.0230619f $X=12.795 $Y=1.53
+ $X2=0 $Y2=0
cc_787 N_A_2122_348#_c_1220_n N_A_1900_107#_M1001_g 0.0137523f $X=12.91 $Y=0.745
+ $X2=0 $Y2=0
cc_788 N_A_2122_348#_c_1222_n N_A_1900_107#_M1001_g 0.00119474f $X=12.795
+ $Y=1.615 $X2=0 $Y2=0
cc_789 N_A_2122_348#_c_1256_p N_A_1900_107#_c_1305_n 0.0386626f $X=12.71
+ $Y=2.435 $X2=0.24 $Y2=0
cc_790 N_A_2122_348#_c_1226_n N_A_1900_107#_c_1305_n 0.0093702f $X=12.795
+ $Y=2.35 $X2=0.24 $Y2=0
cc_791 N_A_2122_348#_c_1227_n N_A_1900_107#_c_1305_n 0.0146366f $X=12.13
+ $Y=2.435 $X2=0.24 $Y2=0
cc_792 N_A_2122_348#_c_1226_n N_A_1900_107#_c_1295_n 0.0213052f $X=12.795
+ $Y=2.35 $X2=0 $Y2=0
cc_793 N_A_2122_348#_c_1220_n N_A_1900_107#_c_1295_n 0.00542111f $X=12.91
+ $Y=0.745 $X2=0 $Y2=0
cc_794 N_A_2122_348#_c_1222_n N_A_1900_107#_c_1295_n 0.00764841f $X=12.795
+ $Y=1.615 $X2=0 $Y2=0
cc_795 N_A_2122_348#_c_1226_n N_A_1900_107#_M1023_g 0.00228834f $X=12.795
+ $Y=2.35 $X2=0 $Y2=0
cc_796 N_A_2122_348#_c_1220_n N_A_1900_107#_M1017_g 7.96424e-19 $X=12.91
+ $Y=0.745 $X2=0 $Y2=0
cc_797 N_A_2122_348#_M1007_g N_A_1900_107#_c_1326_n 7.33647e-19 $X=11.03
+ $Y=0.745 $X2=0 $Y2=0
cc_798 N_A_2122_348#_c_1217_n N_A_1900_107#_c_1302_n 0.0152008f $X=10.945 $Y=2.2
+ $X2=0 $Y2=0
cc_799 N_A_2122_348#_c_1235_n N_A_1900_107#_c_1302_n 0.0329584f $X=11.095
+ $Y=1.395 $X2=0 $Y2=0
cc_800 N_A_2122_348#_M1007_g N_A_1900_107#_c_1302_n 0.013919f $X=11.03 $Y=0.745
+ $X2=0 $Y2=0
cc_801 N_A_2122_348#_c_1217_n N_A_1900_107#_c_1319_n 0.0305231f $X=10.945 $Y=2.2
+ $X2=0 $Y2=0
cc_802 N_A_2122_348#_c_1218_n N_A_1900_107#_c_1319_n 0.0437109f $X=12.71
+ $Y=1.615 $X2=0 $Y2=0
cc_803 N_A_2122_348#_c_1235_n N_A_1900_107#_c_1319_n 0.0232944f $X=11.095
+ $Y=1.395 $X2=0 $Y2=0
cc_804 N_A_2122_348#_c_1227_n N_A_1900_107#_c_1319_n 0.0153902f $X=12.13
+ $Y=2.435 $X2=0 $Y2=0
cc_805 N_A_2122_348#_c_1217_n N_A_1900_107#_c_1320_n 0.00832388f $X=10.945
+ $Y=2.2 $X2=0 $Y2=0
cc_806 N_A_2122_348#_c_1218_n N_A_1900_107#_c_1345_n 0.0225142f $X=12.71
+ $Y=1.615 $X2=0 $Y2=0
cc_807 N_A_2122_348#_c_1256_p N_A_1900_107#_c_1345_n 0.0158769f $X=12.71
+ $Y=2.435 $X2=0 $Y2=0
cc_808 N_A_2122_348#_c_1226_n N_A_1900_107#_c_1345_n 0.0197818f $X=12.795
+ $Y=2.35 $X2=0 $Y2=0
cc_809 N_A_2122_348#_c_1227_n N_A_1900_107#_c_1345_n 0.00464686f $X=12.13
+ $Y=2.435 $X2=0 $Y2=0
cc_810 N_A_2122_348#_c_1218_n N_A_1900_107#_c_1304_n 0.0167269f $X=12.71
+ $Y=1.615 $X2=0 $Y2=0
cc_811 N_A_2122_348#_c_1226_n N_A_1900_107#_c_1304_n 0.0174657f $X=12.795
+ $Y=2.35 $X2=0 $Y2=0
cc_812 N_A_2122_348#_c_1227_n N_A_1900_107#_c_1304_n 0.00161049f $X=12.13
+ $Y=2.435 $X2=0 $Y2=0
cc_813 N_A_2122_348#_c_1222_n N_A_1900_107#_c_1304_n 6.49734e-19 $X=12.795
+ $Y=1.615 $X2=0 $Y2=0
cc_814 N_A_2122_348#_c_1256_p N_VPWR_M1012_d 0.00411908f $X=12.71 $Y=2.435 $X2=0
+ $Y2=0
cc_815 N_A_2122_348#_c_1226_n N_VPWR_M1012_d 3.9721e-19 $X=12.795 $Y=2.35 $X2=0
+ $Y2=0
cc_816 N_A_2122_348#_c_1217_n N_VPWR_c_1502_n 0.0517066f $X=10.945 $Y=2.2 $X2=0
+ $Y2=0
cc_817 N_A_2122_348#_c_1227_n N_VPWR_c_1502_n 0.0159166f $X=12.13 $Y=2.435 $X2=0
+ $Y2=0
cc_818 N_A_2122_348#_c_1256_p N_VPWR_c_1505_n 0.0144616f $X=12.71 $Y=2.435 $X2=0
+ $Y2=0
cc_819 N_A_2122_348#_c_1226_n N_VPWR_c_1505_n 0.0139756f $X=12.795 $Y=2.35 $X2=0
+ $Y2=0
cc_820 N_A_2122_348#_c_1220_n N_VGND_c_1728_n 0.00744773f $X=12.91 $Y=0.745
+ $X2=0 $Y2=0
cc_821 N_A_2122_348#_M1007_g N_VGND_c_1728_n 0.00709087f $X=11.03 $Y=0.745 $X2=0
+ $Y2=0
cc_822 N_A_2122_348#_c_1219_n N_VGND_c_1730_n 0.0249891f $X=12.795 $Y=1.53 $X2=0
+ $Y2=0
cc_823 N_A_2122_348#_c_1220_n N_VGND_c_1730_n 0.0370573f $X=12.91 $Y=0.745 $X2=0
+ $Y2=0
cc_824 N_A_2122_348#_c_1220_n N_VGND_c_1734_n 0.0333924f $X=12.91 $Y=0.745 $X2=0
+ $Y2=0
cc_825 N_A_2122_348#_M1007_g N_VGND_c_1734_n 0.0106681f $X=11.03 $Y=0.745 $X2=0
+ $Y2=0
cc_826 N_A_1900_107#_M1033_g N_A_2937_443#_M1010_g 0.0184764f $X=15.22 $Y=2.59
+ $X2=0 $Y2=0
cc_827 N_A_1900_107#_c_1301_n N_A_2937_443#_M1010_g 0.00815685f $X=15.23 $Y=1.75
+ $X2=0 $Y2=0
cc_828 N_A_1900_107#_M1024_g N_A_2937_443#_M1021_g 0.0145305f $X=15.24 $Y=1.075
+ $X2=0 $Y2=0
cc_829 N_A_1900_107#_M1017_g N_A_2937_443#_c_1446_n 0.00155745f $X=13.87 $Y=1.08
+ $X2=16.56 $Y2=0
cc_830 N_A_1900_107#_M1024_g N_A_2937_443#_c_1446_n 0.0170445f $X=15.24 $Y=1.075
+ $X2=16.56 $Y2=0
cc_831 N_A_1900_107#_c_1301_n N_A_2937_443#_c_1446_n 0.00664239f $X=15.23
+ $Y=1.75 $X2=16.56 $Y2=0
cc_832 N_A_1900_107#_c_1298_n N_A_2937_443#_c_1453_n 0.0170695f $X=14.97
+ $Y=1.835 $X2=8.4 $Y2=0
cc_833 N_A_1900_107#_M1033_g N_A_2937_443#_c_1453_n 0.0241398f $X=15.22 $Y=2.59
+ $X2=8.4 $Y2=0
cc_834 N_A_1900_107#_c_1301_n N_A_2937_443#_c_1453_n 0.0117544f $X=15.23 $Y=1.75
+ $X2=8.4 $Y2=0
cc_835 N_A_1900_107#_c_1301_n N_A_2937_443#_c_1447_n 0.045849f $X=15.23 $Y=1.75
+ $X2=0 $Y2=0
cc_836 N_A_1900_107#_c_1301_n N_A_2937_443#_c_1448_n 0.0221341f $X=15.23 $Y=1.75
+ $X2=0 $Y2=0
cc_837 N_A_1900_107#_M1017_g N_A_2937_443#_c_1449_n 3.63305e-19 $X=13.87 $Y=1.08
+ $X2=0 $Y2=0
cc_838 N_A_1900_107#_c_1298_n N_A_2937_443#_c_1449_n 0.019537f $X=14.97 $Y=1.835
+ $X2=0 $Y2=0
cc_839 N_A_1900_107#_c_1301_n N_A_2937_443#_c_1449_n 0.00400101f $X=15.23
+ $Y=1.75 $X2=0 $Y2=0
cc_840 N_A_1900_107#_c_1319_n N_VPWR_c_1502_n 0.0560882f $X=12.2 $Y=2.085 $X2=0
+ $Y2=0
cc_841 N_A_1900_107#_c_1320_n N_VPWR_c_1502_n 0.0101077f $X=10.725 $Y=2.085
+ $X2=0 $Y2=0
cc_842 N_A_1900_107#_c_1305_n N_VPWR_c_1505_n 0.0138773f $X=12.52 $Y=2.2 $X2=0
+ $Y2=0
cc_843 N_A_1900_107#_c_1295_n N_VPWR_c_1505_n 0.0181063f $X=13.575 $Y=1.835
+ $X2=0 $Y2=0
cc_844 N_A_1900_107#_M1023_g N_VPWR_c_1505_n 0.0871826f $X=13.825 $Y=2.965 $X2=0
+ $Y2=0
cc_845 N_A_1900_107#_c_1304_n N_VPWR_c_1505_n 0.00207801f $X=12.365 $Y=1.985
+ $X2=0 $Y2=0
cc_846 N_A_1900_107#_M1033_g N_VPWR_c_1508_n 0.069435f $X=15.22 $Y=2.59 $X2=0
+ $Y2=0
cc_847 N_A_1900_107#_c_1301_n N_VPWR_c_1508_n 6.61217e-19 $X=15.23 $Y=1.75 $X2=0
+ $Y2=0
cc_848 N_A_1900_107#_c_1305_n N_VPWR_c_1511_n 0.0123644f $X=12.52 $Y=2.2 $X2=0
+ $Y2=0
cc_849 N_A_1900_107#_M1023_g N_VPWR_c_1511_n 0.00945778f $X=13.825 $Y=2.965
+ $X2=0 $Y2=0
cc_850 N_A_1900_107#_M1033_g N_VPWR_c_1511_n 0.00584154f $X=15.22 $Y=2.59 $X2=0
+ $Y2=0
cc_851 N_A_1900_107#_c_1315_n N_VPWR_c_1511_n 0.0106128f $X=9.64 $Y=2.81 $X2=0
+ $Y2=0
cc_852 N_A_1900_107#_M1017_g N_Q_N_c_1683_n 0.0113609f $X=13.87 $Y=1.08 $X2=0
+ $Y2=0
cc_853 N_A_1900_107#_c_1298_n N_Q_N_c_1683_n 0.0175826f $X=14.97 $Y=1.835 $X2=0
+ $Y2=0
cc_854 N_A_1900_107#_M1024_g N_Q_N_c_1683_n 4.15446e-19 $X=15.24 $Y=1.075 $X2=0
+ $Y2=0
cc_855 N_A_1900_107#_c_1300_n N_Q_N_c_1683_n 0.0146054f $X=13.847 $Y=1.835 $X2=0
+ $Y2=0
cc_856 N_A_1900_107#_c_1301_n N_Q_N_c_1683_n 6.74746e-19 $X=15.23 $Y=1.75 $X2=0
+ $Y2=0
cc_857 N_A_1900_107#_M1023_g N_Q_N_c_1685_n 0.00854681f $X=13.825 $Y=2.965 $X2=0
+ $Y2=0
cc_858 N_A_1900_107#_c_1298_n N_Q_N_c_1685_n 0.0320772f $X=14.97 $Y=1.835 $X2=0
+ $Y2=0
cc_859 N_A_1900_107#_M1033_g N_Q_N_c_1685_n 0.00460342f $X=15.22 $Y=2.59 $X2=0
+ $Y2=0
cc_860 N_A_1900_107#_M1017_g N_Q_N_c_1684_n 0.0183957f $X=13.87 $Y=1.08 $X2=0
+ $Y2=0
cc_861 N_A_1900_107#_M1024_g N_Q_N_c_1684_n 0.00360198f $X=15.24 $Y=1.075 $X2=0
+ $Y2=0
cc_862 N_A_1900_107#_M1001_g N_VGND_c_1728_n 0.00577968f $X=12.52 $Y=0.745 $X2=0
+ $Y2=0
cc_863 N_A_1900_107#_M1001_g N_VGND_c_1730_n 0.00582443f $X=12.52 $Y=0.745 $X2=0
+ $Y2=0
cc_864 N_A_1900_107#_c_1295_n N_VGND_c_1730_n 0.00993486f $X=13.575 $Y=1.835
+ $X2=0 $Y2=0
cc_865 N_A_1900_107#_M1017_g N_VGND_c_1730_n 0.0522527f $X=13.87 $Y=1.08 $X2=0
+ $Y2=0
cc_866 N_A_1900_107#_M1024_g N_VGND_c_1732_n 0.0476742f $X=15.24 $Y=1.075 $X2=0
+ $Y2=0
cc_867 N_A_1900_107#_M1016_d N_VGND_c_1734_n 0.00115477f $X=9.5 $Y=0.535 $X2=0
+ $Y2=0
cc_868 N_A_1900_107#_M1001_g N_VGND_c_1734_n 0.031123f $X=12.52 $Y=0.745 $X2=0
+ $Y2=0
cc_869 N_A_1900_107#_M1017_g N_VGND_c_1734_n 0.0144506f $X=13.87 $Y=1.08 $X2=0
+ $Y2=0
cc_870 N_A_1900_107#_M1024_g N_VGND_c_1734_n 0.00672879f $X=15.24 $Y=1.075 $X2=0
+ $Y2=0
cc_871 N_A_1900_107#_c_1326_n N_VGND_c_1734_n 0.035644f $X=10.555 $Y=0.7 $X2=0
+ $Y2=0
cc_872 N_A_1900_107#_c_1303_n N_VGND_c_1734_n 0.0107792f $X=9.91 $Y=0.805 $X2=0
+ $Y2=0
cc_873 N_A_1900_107#_c_1326_n A_2114_107# 4.80934e-19 $X=10.555 $Y=0.7 $X2=0
+ $Y2=0
cc_874 N_A_2937_443#_M1010_g N_VPWR_c_1508_n 0.0718832f $X=16.115 $Y=2.965 $X2=0
+ $Y2=0
cc_875 N_A_2937_443#_c_1453_n N_VPWR_c_1508_n 0.0629871f $X=14.83 $Y=2.34 $X2=0
+ $Y2=0
cc_876 N_A_2937_443#_c_1447_n N_VPWR_c_1508_n 0.0465313f $X=15.995 $Y=1.67 $X2=0
+ $Y2=0
cc_877 N_A_2937_443#_c_1448_n N_VPWR_c_1508_n 0.00137591f $X=15.995 $Y=1.67
+ $X2=0 $Y2=0
cc_878 N_A_2937_443#_M1010_g N_VPWR_c_1511_n 0.0130327f $X=16.115 $Y=2.965 $X2=0
+ $Y2=0
cc_879 N_A_2937_443#_c_1453_n N_VPWR_c_1511_n 0.0143895f $X=14.83 $Y=2.34 $X2=0
+ $Y2=0
cc_880 N_A_2937_443#_c_1446_n N_Q_N_c_1683_n 0.0132269f $X=14.85 $Y=1.075 $X2=0
+ $Y2=0
cc_881 N_A_2937_443#_c_1449_n N_Q_N_c_1683_n 0.0152792f $X=14.84 $Y=1.67 $X2=0
+ $Y2=0
cc_882 N_A_2937_443#_c_1453_n N_Q_N_c_1685_n 0.0645468f $X=14.83 $Y=2.34 $X2=0
+ $Y2=0
cc_883 N_A_2937_443#_c_1449_n N_Q_N_c_1685_n 0.00281856f $X=14.84 $Y=1.67 $X2=0
+ $Y2=0
cc_884 N_A_2937_443#_c_1446_n N_Q_N_c_1684_n 0.0318693f $X=14.85 $Y=1.075 $X2=0
+ $Y2=0
cc_885 N_A_2937_443#_M1010_g N_Q_c_1709_n 0.0476053f $X=16.115 $Y=2.965 $X2=0
+ $Y2=0
cc_886 N_A_2937_443#_M1021_g N_Q_c_1709_n 0.0239988f $X=16.135 $Y=0.91 $X2=0
+ $Y2=0
cc_887 N_A_2937_443#_c_1447_n N_Q_c_1709_n 0.0251095f $X=15.995 $Y=1.67 $X2=0
+ $Y2=0
cc_888 N_A_2937_443#_c_1448_n N_Q_c_1709_n 0.0252537f $X=15.995 $Y=1.67 $X2=0
+ $Y2=0
cc_889 N_A_2937_443#_M1021_g N_VGND_c_1732_n 0.0496278f $X=16.135 $Y=0.91 $X2=0
+ $Y2=0
cc_890 N_A_2937_443#_c_1446_n N_VGND_c_1732_n 0.0381062f $X=14.85 $Y=1.075 $X2=0
+ $Y2=0
cc_891 N_A_2937_443#_c_1447_n N_VGND_c_1732_n 0.0753947f $X=15.995 $Y=1.67 $X2=0
+ $Y2=0
cc_892 N_A_2937_443#_c_1448_n N_VGND_c_1732_n 0.00214709f $X=15.995 $Y=1.67
+ $X2=0 $Y2=0
cc_893 N_A_2937_443#_M1021_g N_VGND_c_1734_n 0.0129444f $X=16.135 $Y=0.91 $X2=0
+ $Y2=0
cc_894 N_A_2937_443#_c_1446_n N_VGND_c_1734_n 0.0192623f $X=14.85 $Y=1.075 $X2=0
+ $Y2=0
cc_895 N_VPWR_c_1511_n N_A_509_608#_M1018_s 0.00228133f $X=16.01 $Y=3.59 $X2=0
+ $Y2=0
cc_896 N_VPWR_c_1511_n N_A_509_608#_M1008_d 0.00218173f $X=16.01 $Y=3.59 $X2=0
+ $Y2=0
cc_897 N_VPWR_c_1511_n N_A_509_608#_c_1619_n 0.0121654f $X=16.01 $Y=3.59
+ $X2=0.24 $Y2=4.07
cc_898 N_VPWR_c_1511_n N_A_509_608#_c_1624_n 0.0147406f $X=16.01 $Y=3.59 $X2=0
+ $Y2=0
cc_899 N_VPWR_c_1496_n A_1134_608# 0.00285582f $X=6.575 $Y=3.59 $X2=0 $Y2=3.985
cc_900 N_VPWR_c_1511_n A_1134_608# 8.598e-19 $X=16.01 $Y=3.59 $X2=0 $Y2=3.985
cc_901 N_VPWR_c_1511_n N_Q_N_M1023_d 0.00221032f $X=16.01 $Y=3.59 $X2=0 $Y2=0
cc_902 N_VPWR_c_1505_n N_Q_N_c_1685_n 0.0677868f $X=13.435 $Y=2.34 $X2=0.24
+ $Y2=4.07
cc_903 N_VPWR_c_1511_n N_Q_N_c_1685_n 0.0381476f $X=16.01 $Y=3.59 $X2=0.24
+ $Y2=4.07
cc_904 N_VPWR_c_1508_n N_Q_c_1709_n 0.0996146f $X=15.725 $Y=2.34 $X2=8.4
+ $Y2=4.07
cc_905 N_VPWR_c_1511_n N_Q_c_1709_n 0.0452076f $X=16.01 $Y=3.59 $X2=8.4 $Y2=4.07
cc_906 N_VPWR_c_1505_n N_VGND_c_1730_n 0.0183727f $X=13.435 $Y=2.34 $X2=0 $Y2=0
cc_907 N_A_509_608#_c_1616_n N_VGND_c_1734_n 0.00248943f $X=4.49 $Y=1.075 $X2=0
+ $Y2=0
cc_908 N_Q_N_c_1683_n N_VGND_c_1730_n 0.0132956f $X=14.255 $Y=1.78 $X2=0 $Y2=0
cc_909 N_Q_N_c_1684_n N_VGND_c_1730_n 0.0445552f $X=14.26 $Y=0.83 $X2=0 $Y2=0
cc_910 N_Q_N_c_1684_n N_VGND_c_1734_n 0.0165861f $X=14.26 $Y=0.83 $X2=0 $Y2=0
cc_911 N_Q_c_1709_n N_VGND_c_1732_n 0.056224f $X=16.525 $Y=0.68 $X2=0 $Y2=0
cc_912 N_Q_c_1709_n N_VGND_c_1734_n 0.0337877f $X=16.525 $Y=0.68 $X2=0 $Y2=0
cc_913 N_VGND_c_1734_n A_2114_107# 0.00225203f $X=16.03 $Y=0.48 $X2=0 $Y2=0
cc_914 N_VGND_c_1728_n A_2412_107# 0.00682976f $X=12.09 $Y=0.48 $X2=0 $Y2=0
cc_915 N_VGND_c_1734_n A_2412_107# 0.00271077f $X=16.03 $Y=0.48 $X2=0 $Y2=0
