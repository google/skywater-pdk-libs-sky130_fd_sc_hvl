* File: sky130_fd_sc_hvl__o22a_1.pxi.spice
* Created: Wed Sep  2 09:09:06 2020
* 
x_PM_SKY130_FD_SC_HVL__O22A_1%VNB N_VNB_M1003_b VNB N_VNB_c_4_p VNB
+ PM_SKY130_FD_SC_HVL__O22A_1%VNB
x_PM_SKY130_FD_SC_HVL__O22A_1%VPB N_VPB_M1008_b VPB N_VPB_c_39_p VPB
+ PM_SKY130_FD_SC_HVL__O22A_1%VPB
x_PM_SKY130_FD_SC_HVL__O22A_1%A_87_81# N_A_87_81#_M1002_d N_A_87_81#_M1000_d
+ N_A_87_81#_c_122_p N_A_87_81#_c_85_p N_A_87_81#_c_73_n N_A_87_81#_c_87_p
+ N_A_87_81#_c_127_p N_A_87_81#_c_74_n N_A_87_81#_c_88_p N_A_87_81#_c_104_p
+ N_A_87_81#_c_77_n N_A_87_81#_c_78_n N_A_87_81#_M1003_g N_A_87_81#_M1008_g
+ PM_SKY130_FD_SC_HVL__O22A_1%A_87_81#
x_PM_SKY130_FD_SC_HVL__O22A_1%A1 N_A1_M1006_g N_A1_c_150_n N_A1_c_151_n
+ N_A1_c_152_n N_A1_c_153_n N_A1_c_154_n N_A1_c_210_p N_A1_c_155_n N_A1_c_156_n
+ A1 A1 N_A1_M1007_g N_A1_c_160_n N_A1_c_190_n A1 A1 N_A1_c_161_n
+ PM_SKY130_FD_SC_HVL__O22A_1%A1
x_PM_SKY130_FD_SC_HVL__O22A_1%B1 N_B1_M1002_g N_B1_M1009_g B1 N_B1_c_238_n
+ PM_SKY130_FD_SC_HVL__O22A_1%B1
x_PM_SKY130_FD_SC_HVL__O22A_1%B2 B2 B2 N_B2_M1004_g N_B2_M1000_g
+ PM_SKY130_FD_SC_HVL__O22A_1%B2
x_PM_SKY130_FD_SC_HVL__O22A_1%A2 A2 A2 N_A2_M1001_g N_A2_M1005_g
+ PM_SKY130_FD_SC_HVL__O22A_1%A2
x_PM_SKY130_FD_SC_HVL__O22A_1%X N_X_M1003_s N_X_M1008_s X X X X X X X
+ N_X_c_335_n PM_SKY130_FD_SC_HVL__O22A_1%X
x_PM_SKY130_FD_SC_HVL__O22A_1%VPWR N_VPWR_M1008_d N_VPWR_M1006_d VPWR
+ N_VPWR_c_349_n N_VPWR_c_352_n N_VPWR_c_355_n PM_SKY130_FD_SC_HVL__O22A_1%VPWR
x_PM_SKY130_FD_SC_HVL__O22A_1%VGND N_VGND_M1003_d N_VGND_M1001_d VGND
+ N_VGND_c_386_n N_VGND_c_388_n N_VGND_c_390_n PM_SKY130_FD_SC_HVL__O22A_1%VGND
x_PM_SKY130_FD_SC_HVL__O22A_1%A_354_107# N_A_354_107#_M1007_d
+ N_A_354_107#_M1004_d N_A_354_107#_c_434_n N_A_354_107#_c_429_n
+ N_A_354_107#_c_431_n N_A_354_107#_c_437_n
+ PM_SKY130_FD_SC_HVL__O22A_1%A_354_107#
cc_1 N_VNB_M1003_b N_A_87_81#_c_73_n 0.01603f $X=-0.33 $Y=-0.265 $X2=1.63
+ $Y2=1.51
cc_2 N_VNB_M1003_b N_A_87_81#_c_74_n 0.00131598f $X=-0.33 $Y=-0.265 $X2=1.715
+ $Y2=1.425
cc_3 N_VNB_M1003_b N_A_87_81#_M1003_g 0.091313f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=0.91
cc_4 N_VNB_c_4_p N_A_87_81#_M1003_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.685 $Y2=0.91
cc_5 N_VNB_M1003_b N_A1_c_150_n 0.00304656f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_M1003_b N_A1_c_151_n 0.00191791f $X=-0.33 $Y=-0.265 $X2=3.43
+ $Y2=2.385
cc_7 N_VNB_M1003_b N_A1_c_152_n 7.00144e-19 $X=-0.33 $Y=-0.265 $X2=0.915
+ $Y2=2.385
cc_8 N_VNB_M1003_b N_A1_c_153_n 0.00173655f $X=-0.33 $Y=-0.265 $X2=1.715
+ $Y2=1.22
cc_9 N_VNB_M1003_b N_A1_c_154_n 0.0154805f $X=-0.33 $Y=-0.265 $X2=1.715
+ $Y2=1.425
cc_10 N_VNB_M1003_b N_A1_c_155_n 0.0817952f $X=-0.33 $Y=-0.265 $X2=3.515
+ $Y2=2.755
cc_11 N_VNB_M1003_b N_A1_c_156_n 0.00442641f $X=-0.33 $Y=-0.265 $X2=3.515
+ $Y2=3.59
cc_12 N_VNB_M1003_b A1 0.00366195f $X=-0.33 $Y=-0.265 $X2=2.69 $Y2=0.917
cc_13 N_VNB_M1003_b N_A1_M1007_g 0.0871861f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.965
cc_14 N_VNB_c_4_p N_A1_M1007_g 0.00137776f $X=0.24 $Y=0 $X2=0.685 $Y2=2.965
cc_15 N_VNB_M1003_b N_A1_c_160_n 0.00504147f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_16 N_VNB_M1003_b N_A1_c_161_n 3.75344e-19 $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_17 N_VNB_M1003_b N_B1_M1002_g 0.0389595f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_18 N_VNB_M1003_b B1 0.00169403f $X=-0.33 $Y=-0.265 $X2=1.63 $Y2=1.51
cc_19 N_VNB_M1003_b N_B1_c_238_n 0.0461599f $X=-0.33 $Y=-0.265 $X2=0.915
+ $Y2=2.385
cc_20 N_VNB_M1003_b N_B2_M1004_g 0.0797841f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_21 N_VNB_M1003_b A2 0.00643091f $X=-0.33 $Y=-0.265 $X2=3.375 $Y2=2.215
cc_22 N_VNB_M1003_b N_A2_M1001_g 0.0835744f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_23 N_VNB_c_4_p N_A2_M1001_g 9.82123e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_24 N_VNB_M1003_b N_X_c_335_n 0.0670044f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_25 N_VNB_c_4_p N_X_c_335_n 5.92913e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_26 N_VNB_M1003_b N_VGND_c_386_n 0.0438029f $X=-0.33 $Y=-0.265 $X2=0.915
+ $Y2=1.51
cc_27 N_VNB_c_4_p N_VGND_c_386_n 0.00252021f $X=0.24 $Y=0 $X2=0.915 $Y2=1.51
cc_28 N_VNB_M1003_b N_VGND_c_388_n 0.118426f $X=-0.33 $Y=-0.265 $X2=3.515
+ $Y2=2.755
cc_29 N_VNB_c_4_p N_VGND_c_388_n 0.00368339f $X=0.24 $Y=0 $X2=3.515 $Y2=2.755
cc_30 N_VNB_M1003_b N_VGND_c_390_n 0.0820882f $X=-0.33 $Y=-0.265 $X2=0.75
+ $Y2=1.51
cc_31 N_VNB_c_4_p N_VGND_c_390_n 0.564092f $X=0.24 $Y=0 $X2=0.75 $Y2=1.51
cc_32 N_VNB_M1003_b N_A_354_107#_c_429_n 0.114684f $X=-0.33 $Y=-0.265 $X2=3.43
+ $Y2=2.385
cc_33 N_VNB_c_4_p N_A_354_107#_c_429_n 0.0054003f $X=0.24 $Y=0 $X2=3.43
+ $Y2=2.385
cc_34 N_VNB_M1003_b N_A_354_107#_c_431_n 0.0249724f $X=-0.33 $Y=-0.265 $X2=0.915
+ $Y2=2.385
cc_35 N_VNB_c_4_p N_A_354_107#_c_431_n 0.00109614f $X=0.24 $Y=0 $X2=0.915
+ $Y2=2.385
cc_36 N_VPB_M1008_b N_A_87_81#_c_77_n 0.00449906f $X=-0.33 $Y=1.885 $X2=3.555
+ $Y2=2.47
cc_37 N_VPB_M1008_b N_A_87_81#_c_78_n 0.00120153f $X=-0.33 $Y=1.885 $X2=3.515
+ $Y2=2.755
cc_38 VPB N_A_87_81#_c_78_n 8.01732e-19 $X=0 $Y=3.955 $X2=3.515 $Y2=2.755
cc_39 N_VPB_c_39_p N_A_87_81#_c_78_n 0.0130099f $X=5.04 $Y=4.07 $X2=3.515
+ $Y2=2.755
cc_40 N_VPB_M1008_b N_A_87_81#_M1003_g 0.0665145f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=0.91
cc_41 VPB N_A_87_81#_M1003_g 0.00970178f $X=0 $Y=3.955 $X2=0.685 $Y2=0.91
cc_42 N_VPB_c_39_p N_A_87_81#_M1003_g 0.015205f $X=5.04 $Y=4.07 $X2=0.685
+ $Y2=0.91
cc_43 N_VPB_M1008_b N_A1_M1006_g 0.0413246f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_44 VPB N_A1_M1006_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_45 N_VPB_c_39_p N_A1_M1006_g 0.013806f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_46 N_VPB_M1008_b N_A1_c_150_n 0.00296641f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_47 N_VPB_M1008_b N_A1_c_155_n 0.0263573f $X=-0.33 $Y=1.885 $X2=3.515
+ $Y2=2.755
cc_48 N_VPB_M1008_b N_A1_M1007_g 0.0304308f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.965
cc_49 N_VPB_M1008_b N_B1_M1009_g 0.0417072f $X=-0.33 $Y=1.885 $X2=0.75 $Y2=1.595
cc_50 VPB N_B1_M1009_g 0.00970178f $X=0 $Y=3.955 $X2=0.75 $Y2=1.595
cc_51 N_VPB_c_39_p N_B1_M1009_g 0.013715f $X=5.04 $Y=4.07 $X2=0.75 $Y2=1.595
cc_52 N_VPB_M1008_b B1 0.00232351f $X=-0.33 $Y=1.885 $X2=1.63 $Y2=1.51
cc_53 N_VPB_M1008_b N_B1_c_238_n 0.0213848f $X=-0.33 $Y=1.885 $X2=0.915
+ $Y2=2.385
cc_54 N_VPB_M1008_b N_B2_M1004_g 0.0528469f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_55 VPB N_B2_M1004_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_56 N_VPB_c_39_p N_B2_M1004_g 0.015205f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_57 N_VPB_M1008_b A2 0.00266475f $X=-0.33 $Y=1.885 $X2=3.375 $Y2=2.215
cc_58 N_VPB_M1008_b N_A2_M1001_g 0.0520888f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_59 VPB N_A2_M1001_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_60 N_VPB_c_39_p N_A2_M1001_g 0.0159377f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_61 N_VPB_M1008_b N_X_c_335_n 0.0684039f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_62 VPB N_X_c_335_n 7.75439e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_63 N_VPB_c_39_p N_X_c_335_n 0.0133691f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_64 N_VPB_M1008_b N_VPWR_c_349_n 0.00770895f $X=-0.33 $Y=1.885 $X2=3.555
+ $Y2=2.47
cc_65 VPB N_VPWR_c_349_n 0.0104029f $X=0 $Y=3.955 $X2=3.555 $Y2=2.47
cc_66 N_VPB_c_39_p N_VPWR_c_349_n 0.136585f $X=5.04 $Y=4.07 $X2=3.555 $Y2=2.47
cc_67 N_VPB_M1008_b N_VPWR_c_352_n 0.0781261f $X=-0.33 $Y=1.885 $X2=3.515
+ $Y2=3.59
cc_68 VPB N_VPWR_c_352_n 0.00532377f $X=0 $Y=3.955 $X2=3.515 $Y2=3.59
cc_69 N_VPB_c_39_p N_VPWR_c_352_n 0.0603963f $X=5.04 $Y=4.07 $X2=3.515 $Y2=3.59
cc_70 N_VPB_M1008_b N_VPWR_c_355_n 0.04924f $X=-0.33 $Y=1.885 $X2=3.515 $Y2=2.34
cc_71 VPB N_VPWR_c_355_n 0.560211f $X=0 $Y=3.955 $X2=3.515 $Y2=2.34
cc_72 N_VPB_c_39_p N_VPWR_c_355_n 0.0213197f $X=5.04 $Y=4.07 $X2=3.515 $Y2=2.34
cc_73 N_A_87_81#_c_78_n N_A1_M1006_g 5.56805e-19 $X=3.515 $Y=2.755 $X2=0 $Y2=0
cc_74 N_A_87_81#_c_85_p N_A1_c_150_n 0.00909816f $X=0.75 $Y=2.3 $X2=-0.33
+ $Y2=-0.265
cc_75 N_A_87_81#_c_73_n N_A1_c_150_n 0.0269403f $X=1.63 $Y=1.51 $X2=-0.33
+ $Y2=-0.265
cc_76 N_A_87_81#_c_87_p N_A1_c_150_n 0.0408729f $X=3.43 $Y=2.385 $X2=-0.33
+ $Y2=-0.265
cc_77 N_A_87_81#_c_88_p N_A1_c_150_n 0.00550377f $X=2.255 $Y=1.135 $X2=-0.33
+ $Y2=-0.265
cc_78 N_A_87_81#_M1003_g N_A1_c_150_n 9.79445e-19 $X=0.685 $Y=0.91 $X2=-0.33
+ $Y2=-0.265
cc_79 N_A_87_81#_c_73_n N_A1_c_151_n 0.00199069f $X=1.63 $Y=1.51 $X2=0.24 $Y2=0
cc_80 N_A_87_81#_c_88_p N_A1_c_152_n 0.0245104f $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_81 N_A_87_81#_c_73_n N_A1_c_153_n 0.0129574f $X=1.63 $Y=1.51 $X2=0 $Y2=0
cc_82 N_A_87_81#_c_74_n N_A1_c_153_n 0.00197712f $X=1.715 $Y=1.425 $X2=0 $Y2=0
cc_83 N_A_87_81#_c_88_p N_A1_c_153_n 0.0108241f $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_84 N_A_87_81#_M1002_d N_A1_c_156_n 0.00195711f $X=2.55 $Y=0.535 $X2=2.64
+ $Y2=0
cc_85 N_A_87_81#_c_88_p N_A1_c_156_n 0.0128983f $X=2.255 $Y=1.135 $X2=2.64 $Y2=0
cc_86 N_A_87_81#_M1002_d A1 5.94823e-19 $X=2.55 $Y=0.535 $X2=0 $Y2=0
cc_87 N_A_87_81#_c_88_p A1 0.00314976f $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_88 N_A_87_81#_c_85_p N_A1_M1007_g 0.00259662f $X=0.75 $Y=2.3 $X2=0 $Y2=0
cc_89 N_A_87_81#_c_73_n N_A1_M1007_g 0.0326273f $X=1.63 $Y=1.51 $X2=0 $Y2=0
cc_90 N_A_87_81#_c_87_p N_A1_M1007_g 0.0148039f $X=3.43 $Y=2.385 $X2=0 $Y2=0
cc_91 N_A_87_81#_c_74_n N_A1_M1007_g 0.00738152f $X=1.715 $Y=1.425 $X2=0 $Y2=0
cc_92 N_A_87_81#_c_88_p N_A1_M1007_g 7.27355e-19 $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_93 N_A_87_81#_c_104_p N_A1_M1007_g 0.00968422f $X=1.8 $Y=1.135 $X2=0 $Y2=0
cc_94 N_A_87_81#_M1003_g N_A1_M1007_g 0.0411388f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_95 N_A_87_81#_c_88_p N_A1_c_190_n 2.62416e-19 $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_96 N_A_87_81#_c_74_n N_B1_M1002_g 0.00255676f $X=1.715 $Y=1.425 $X2=0 $Y2=0
cc_97 N_A_87_81#_c_88_p N_B1_M1002_g 0.0457447f $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_98 N_A_87_81#_c_87_p N_B1_M1009_g 0.0326935f $X=3.43 $Y=2.385 $X2=0 $Y2=0
cc_99 N_A_87_81#_c_87_p B1 0.0278741f $X=3.43 $Y=2.385 $X2=0 $Y2=0
cc_100 N_A_87_81#_c_73_n N_B1_c_238_n 5.87499e-19 $X=1.63 $Y=1.51 $X2=0 $Y2=0
cc_101 N_A_87_81#_c_87_p N_B1_c_238_n 0.00280983f $X=3.43 $Y=2.385 $X2=0 $Y2=0
cc_102 N_A_87_81#_c_88_p N_B1_c_238_n 2.84686e-19 $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_103 N_A_87_81#_c_87_p B2 0.0209073f $X=3.43 $Y=2.385 $X2=0 $Y2=0
cc_104 N_A_87_81#_c_87_p N_B2_M1004_g 0.0334279f $X=3.43 $Y=2.385 $X2=0 $Y2=0
cc_105 N_A_87_81#_c_88_p N_B2_M1004_g 0.00124004f $X=2.255 $Y=1.135 $X2=0 $Y2=0
cc_106 N_A_87_81#_c_77_n N_B2_M1004_g 0.00106231f $X=3.555 $Y=2.47 $X2=0 $Y2=0
cc_107 N_A_87_81#_c_78_n N_B2_M1004_g 0.0010792f $X=3.515 $Y=2.755 $X2=0 $Y2=0
cc_108 N_A_87_81#_c_77_n A2 0.0124239f $X=3.555 $Y=2.47 $X2=0 $Y2=0
cc_109 N_A_87_81#_c_77_n N_A2_M1001_g 0.00585535f $X=3.555 $Y=2.47 $X2=0 $Y2=0
cc_110 N_A_87_81#_c_78_n N_A2_M1001_g 0.0203738f $X=3.515 $Y=2.755 $X2=0 $Y2=0
cc_111 N_A_87_81#_c_122_p N_X_c_335_n 0.0121432f $X=0.75 $Y=1.595 $X2=0 $Y2=0
cc_112 N_A_87_81#_c_85_p N_X_c_335_n 0.044421f $X=0.75 $Y=2.3 $X2=0 $Y2=0
cc_113 N_A_87_81#_M1003_g N_X_c_335_n 0.0363039f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_114 N_A_87_81#_c_87_p N_VPWR_M1008_d 0.0402229f $X=3.43 $Y=2.385 $X2=0 $Y2=0
cc_115 N_A_87_81#_c_87_p N_VPWR_c_349_n 0.158832f $X=3.43 $Y=2.385 $X2=5.04
+ $Y2=0
cc_116 N_A_87_81#_c_127_p N_VPWR_c_349_n 0.0265491f $X=0.915 $Y=2.385 $X2=5.04
+ $Y2=0
cc_117 N_A_87_81#_c_78_n N_VPWR_c_349_n 0.0473994f $X=3.515 $Y=2.755 $X2=5.04
+ $Y2=0
cc_118 N_A_87_81#_M1003_g N_VPWR_c_349_n 0.0582262f $X=0.685 $Y=0.91 $X2=5.04
+ $Y2=0
cc_119 N_A_87_81#_c_77_n N_VPWR_c_352_n 0.0215277f $X=3.555 $Y=2.47 $X2=2.64
+ $Y2=0
cc_120 N_A_87_81#_c_78_n N_VPWR_c_352_n 0.0902913f $X=3.515 $Y=2.755 $X2=2.64
+ $Y2=0
cc_121 N_A_87_81#_M1000_d N_VPWR_c_355_n 0.00221032f $X=3.375 $Y=2.215 $X2=0
+ $Y2=0
cc_122 N_A_87_81#_c_78_n N_VPWR_c_355_n 0.0308536f $X=3.515 $Y=2.755 $X2=0 $Y2=0
cc_123 N_A_87_81#_M1003_g N_VPWR_c_355_n 0.00912737f $X=0.685 $Y=0.91 $X2=0
+ $Y2=0
cc_124 N_A_87_81#_c_87_p A_533_443# 0.0038117f $X=3.43 $Y=2.385 $X2=0 $Y2=0
cc_125 N_A_87_81#_c_122_p N_VGND_c_386_n 0.0266685f $X=0.75 $Y=1.595 $X2=0.24
+ $Y2=0
cc_126 N_A_87_81#_c_73_n N_VGND_c_386_n 0.036029f $X=1.63 $Y=1.51 $X2=0.24 $Y2=0
cc_127 N_A_87_81#_c_74_n N_VGND_c_386_n 0.00177809f $X=1.715 $Y=1.425 $X2=0.24
+ $Y2=0
cc_128 N_A_87_81#_c_104_p N_VGND_c_386_n 0.0136768f $X=1.8 $Y=1.135 $X2=0.24
+ $Y2=0
cc_129 N_A_87_81#_M1003_g N_VGND_c_386_n 0.0525695f $X=0.685 $Y=0.91 $X2=0.24
+ $Y2=0
cc_130 N_A_87_81#_M1002_d N_VGND_c_390_n 2.74258e-19 $X=2.55 $Y=0.535 $X2=2.64
+ $Y2=0.057
cc_131 N_A_87_81#_c_88_p N_VGND_c_390_n 0.025857f $X=2.255 $Y=1.135 $X2=2.64
+ $Y2=0.057
cc_132 N_A_87_81#_c_104_p N_VGND_c_390_n 0.00443f $X=1.8 $Y=1.135 $X2=2.64
+ $Y2=0.057
cc_133 N_A_87_81#_M1003_g N_VGND_c_390_n 0.00871294f $X=0.685 $Y=0.91 $X2=2.64
+ $Y2=0.057
cc_134 N_A_87_81#_c_88_p N_A_354_107#_M1007_d 0.00480998f $X=2.255 $Y=1.135
+ $X2=0 $Y2=0
cc_135 N_A_87_81#_c_88_p N_A_354_107#_c_434_n 0.0223869f $X=2.255 $Y=1.135 $X2=0
+ $Y2=0
cc_136 N_A_87_81#_c_104_p N_A_354_107#_c_434_n 0.00175421f $X=1.8 $Y=1.135 $X2=0
+ $Y2=0
cc_137 N_A_87_81#_c_88_p N_A_354_107#_c_429_n 0.0271869f $X=2.255 $Y=1.135
+ $X2=0.24 $Y2=0
cc_138 N_A_87_81#_c_88_p N_A_354_107#_c_437_n 0.00650991f $X=2.255 $Y=1.135
+ $X2=0 $Y2=0
cc_139 N_A1_c_152_n N_B1_M1002_g 0.00695268f $X=2.605 $Y=1.485 $X2=0 $Y2=0
cc_140 N_A1_c_153_n N_B1_M1002_g 0.00169559f $X=2.15 $Y=1.485 $X2=0 $Y2=0
cc_141 N_A1_c_156_n N_B1_M1002_g 0.0033676f $X=2.69 $Y=1.315 $X2=0 $Y2=0
cc_142 N_A1_M1007_g N_B1_M1002_g 0.0596802f $X=1.52 $Y=0.91 $X2=0 $Y2=0
cc_143 N_A1_c_150_n B1 0.0218469f $X=1.98 $Y=1.915 $X2=0 $Y2=0
cc_144 N_A1_c_151_n B1 0.00164667f $X=2.065 $Y=1.775 $X2=0 $Y2=0
cc_145 N_A1_c_152_n B1 0.0189327f $X=2.605 $Y=1.485 $X2=0 $Y2=0
cc_146 N_A1_c_156_n B1 0.0116066f $X=2.69 $Y=1.315 $X2=0 $Y2=0
cc_147 N_A1_M1007_g B1 2.33422e-19 $X=1.52 $Y=0.91 $X2=0 $Y2=0
cc_148 N_A1_c_150_n N_B1_c_238_n 0.0109123f $X=1.98 $Y=1.915 $X2=0 $Y2=0
cc_149 N_A1_c_151_n N_B1_c_238_n 0.0108061f $X=2.065 $Y=1.775 $X2=0 $Y2=0
cc_150 N_A1_c_152_n N_B1_c_238_n 0.019573f $X=2.605 $Y=1.485 $X2=0 $Y2=0
cc_151 N_A1_c_153_n N_B1_c_238_n 0.00226722f $X=2.15 $Y=1.485 $X2=0 $Y2=0
cc_152 N_A1_c_156_n N_B1_c_238_n 0.00398118f $X=2.69 $Y=1.315 $X2=0 $Y2=0
cc_153 A1 B2 0.0209618f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A1_c_156_n N_B2_M1004_g 0.00415828f $X=2.69 $Y=1.315 $X2=0 $Y2=0
cc_155 A1 N_B2_M1004_g 0.012245f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A1_c_160_n N_B2_M1004_g 0.0195216f $X=3.615 $Y=1.305 $X2=0 $Y2=0
cc_157 N_A1_c_190_n N_B2_M1004_g 0.00566809f $X=3.13 $Y=1.305 $X2=0 $Y2=0
cc_158 N_A1_c_210_p A2 0.0160417f $X=4.715 $Y=1.545 $X2=0 $Y2=0
cc_159 N_A1_c_155_n A2 0.00306325f $X=4.715 $Y=1.545 $X2=0 $Y2=0
cc_160 N_A1_c_160_n A2 0.0501655f $X=3.615 $Y=1.305 $X2=0 $Y2=0
cc_161 N_A1_c_154_n N_A2_M1001_g 0.0249171f $X=4.55 $Y=1.315 $X2=0 $Y2=0
cc_162 N_A1_c_210_p N_A2_M1001_g 0.00172903f $X=4.715 $Y=1.545 $X2=0 $Y2=0
cc_163 N_A1_c_155_n N_A2_M1001_g 0.168003f $X=4.715 $Y=1.545 $X2=0 $Y2=0
cc_164 N_A1_c_161_n N_A2_M1001_g 0.00596899f $X=3.71 $Y=1.305 $X2=0 $Y2=0
cc_165 N_A1_M1006_g N_VPWR_c_352_n 0.105089f $X=4.615 $Y=2.965 $X2=2.64 $Y2=0
cc_166 N_A1_c_210_p N_VPWR_c_352_n 0.0265705f $X=4.715 $Y=1.545 $X2=2.64 $Y2=0
cc_167 N_A1_c_155_n N_VPWR_c_352_n 0.00149654f $X=4.715 $Y=1.545 $X2=2.64 $Y2=0
cc_168 N_A1_M1006_g N_VPWR_c_355_n 0.0026592f $X=4.615 $Y=2.965 $X2=0 $Y2=0
cc_169 N_A1_c_154_n N_VGND_M1001_d 0.00244953f $X=4.55 $Y=1.315 $X2=0 $Y2=0
cc_170 N_A1_M1007_g N_VGND_c_386_n 0.0367292f $X=1.52 $Y=0.91 $X2=0.24 $Y2=0
cc_171 N_A1_c_154_n N_VGND_c_388_n 0.0736297f $X=4.55 $Y=1.315 $X2=0 $Y2=0
cc_172 N_A1_c_155_n N_VGND_c_388_n 0.00376999f $X=4.715 $Y=1.545 $X2=0 $Y2=0
cc_173 N_A1_c_154_n N_VGND_c_390_n 0.00803105f $X=4.55 $Y=1.315 $X2=2.64
+ $Y2=0.057
cc_174 N_A1_c_156_n N_VGND_c_390_n 5.83379e-19 $X=2.69 $Y=1.315 $X2=2.64
+ $Y2=0.057
cc_175 A1 N_VGND_c_390_n 0.00509078f $X=3.035 $Y=1.21 $X2=2.64 $Y2=0.057
cc_176 N_A1_M1007_g N_VGND_c_390_n 0.0137638f $X=1.52 $Y=0.91 $X2=2.64 $Y2=0.057
cc_177 N_A1_c_160_n N_VGND_c_390_n 0.00109866f $X=3.615 $Y=1.305 $X2=2.64
+ $Y2=0.057
cc_178 N_A1_c_190_n N_VGND_c_390_n 0.00853992f $X=3.13 $Y=1.305 $X2=2.64
+ $Y2=0.057
cc_179 N_A1_c_161_n N_VGND_c_390_n 8.39007e-19 $X=3.71 $Y=1.305 $X2=2.64
+ $Y2=0.057
cc_180 N_A1_c_160_n N_A_354_107#_M1004_d 0.00178683f $X=3.615 $Y=1.305 $X2=0
+ $Y2=0
cc_181 N_A1_M1007_g N_A_354_107#_c_434_n 0.00946918f $X=1.52 $Y=0.91 $X2=0 $Y2=0
cc_182 N_A1_M1007_g N_A_354_107#_c_431_n 0.00122863f $X=1.52 $Y=0.91 $X2=0 $Y2=0
cc_183 N_A1_c_160_n N_A_354_107#_c_437_n 0.0161083f $X=3.615 $Y=1.305 $X2=0
+ $Y2=0
cc_184 B1 B2 0.0262162f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_185 N_B1_c_238_n B2 0.00141934f $X=2.495 $Y=1.89 $X2=0 $Y2=0
cc_186 N_B1_M1002_g N_B2_M1004_g 0.0257392f $X=2.3 $Y=0.91 $X2=0 $Y2=0
cc_187 B1 N_B2_M1004_g 0.00265741f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_188 N_B1_c_238_n N_B2_M1004_g 0.165372f $X=2.495 $Y=1.89 $X2=0 $Y2=0
cc_189 N_B1_M1009_g N_VPWR_c_349_n 0.0992216f $X=2.415 $Y=2.965 $X2=5.04 $Y2=0
cc_190 N_B1_M1009_g N_VPWR_c_355_n 0.00250239f $X=2.415 $Y=2.965 $X2=0 $Y2=0
cc_191 N_B1_M1002_g N_VGND_c_386_n 9.68292e-19 $X=2.3 $Y=0.91 $X2=0.24 $Y2=0
cc_192 N_B1_M1002_g N_VGND_c_390_n 0.00764436f $X=2.3 $Y=0.91 $X2=2.64 $Y2=0.057
cc_193 N_B1_M1002_g N_A_354_107#_c_434_n 0.0125995f $X=2.3 $Y=0.91 $X2=0 $Y2=0
cc_194 N_B1_M1002_g N_A_354_107#_c_429_n 0.0179559f $X=2.3 $Y=0.91 $X2=0.24
+ $Y2=0
cc_195 N_B1_M1002_g N_A_354_107#_c_431_n 8.55986e-19 $X=2.3 $Y=0.91 $X2=0 $Y2=0
cc_196 B2 A2 0.0216273f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_197 N_B2_M1004_g A2 0.00313929f $X=3.125 $Y=0.91 $X2=0 $Y2=0
cc_198 B2 N_A2_M1001_g 0.00144427f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_199 N_B2_M1004_g N_A2_M1001_g 0.0828163f $X=3.125 $Y=0.91 $X2=0 $Y2=0
cc_200 N_B2_M1004_g N_VPWR_c_349_n 0.0642653f $X=3.125 $Y=0.91 $X2=5.04 $Y2=0
cc_201 N_B2_M1004_g N_VPWR_c_355_n 0.00770765f $X=3.125 $Y=0.91 $X2=0 $Y2=0
cc_202 N_B2_M1004_g N_VGND_c_388_n 4.16979e-19 $X=3.125 $Y=0.91 $X2=0 $Y2=0
cc_203 N_B2_M1004_g N_VGND_c_390_n 0.0102125f $X=3.125 $Y=0.91 $X2=2.64
+ $Y2=0.057
cc_204 N_B2_M1004_g N_A_354_107#_c_429_n 0.0220558f $X=3.125 $Y=0.91 $X2=0.24
+ $Y2=0
cc_205 N_B2_M1004_g N_A_354_107#_c_437_n 0.017362f $X=3.125 $Y=0.91 $X2=0 $Y2=0
cc_206 N_A2_M1001_g N_VPWR_c_349_n 5.00981e-19 $X=3.905 $Y=0.91 $X2=5.04 $Y2=0
cc_207 A2 N_VPWR_c_352_n 0.0179666f $X=3.995 $Y=1.58 $X2=2.64 $Y2=0
cc_208 N_A2_M1001_g N_VPWR_c_352_n 0.0840153f $X=3.905 $Y=0.91 $X2=2.64 $Y2=0
cc_209 N_A2_M1001_g N_VPWR_c_355_n 0.0101542f $X=3.905 $Y=0.91 $X2=0 $Y2=0
cc_210 N_A2_M1001_g N_VGND_c_388_n 0.0388882f $X=3.905 $Y=0.91 $X2=0 $Y2=0
cc_211 N_A2_M1001_g N_VGND_c_390_n 0.0057771f $X=3.905 $Y=0.91 $X2=2.64
+ $Y2=0.057
cc_212 N_A2_M1001_g N_A_354_107#_c_429_n 0.00113335f $X=3.905 $Y=0.91 $X2=0.24
+ $Y2=0
cc_213 N_A2_M1001_g N_A_354_107#_c_437_n 0.0122264f $X=3.905 $Y=0.91 $X2=0 $Y2=0
cc_214 N_X_c_335_n N_VPWR_c_349_n 0.047403f $X=0.295 $Y=0.66 $X2=5.04 $Y2=0
cc_215 N_X_M1008_s N_VPWR_c_355_n 0.00221032f $X=0.15 $Y=2.215 $X2=0 $Y2=0
cc_216 N_X_c_335_n N_VPWR_c_355_n 0.0358265f $X=0.295 $Y=0.66 $X2=0 $Y2=0
cc_217 N_X_c_335_n N_VGND_c_386_n 0.0316846f $X=0.295 $Y=0.66 $X2=0.24 $Y2=0
cc_218 N_X_M1003_s N_VGND_c_390_n 0.00221032f $X=0.15 $Y=0.535 $X2=2.64
+ $Y2=0.057
cc_219 N_X_c_335_n N_VGND_c_390_n 0.0267838f $X=0.295 $Y=0.66 $X2=2.64 $Y2=0.057
cc_220 N_VPWR_c_349_n A_533_443# 0.00109358f $X=3.165 $Y=3.59 $X2=0 $Y2=3.985
cc_221 N_VGND_c_386_n N_A_354_107#_c_434_n 0.019114f $X=0.645 $Y=0.48 $X2=0
+ $Y2=0
cc_222 N_VGND_c_390_n N_A_354_107#_c_434_n 0.0203334f $X=5.08 $Y=0.48 $X2=0
+ $Y2=0
cc_223 N_VGND_c_388_n N_A_354_107#_c_429_n 0.00397098f $X=4 $Y=0.48 $X2=0.24
+ $Y2=0
cc_224 N_VGND_c_390_n N_A_354_107#_c_429_n 0.0564486f $X=5.08 $Y=0.48 $X2=0.24
+ $Y2=0
cc_225 N_VGND_c_386_n N_A_354_107#_c_431_n 0.00277036f $X=0.645 $Y=0.48 $X2=0
+ $Y2=0
cc_226 N_VGND_c_390_n N_A_354_107#_c_431_n 0.0114444f $X=5.08 $Y=0.48 $X2=0
+ $Y2=0
cc_227 N_VGND_c_388_n N_A_354_107#_c_437_n 0.0369819f $X=4 $Y=0.48 $X2=0 $Y2=0
cc_228 N_VGND_c_390_n N_A_354_107#_c_437_n 0.0209946f $X=5.08 $Y=0.48 $X2=0
+ $Y2=0
