* File: sky130_fd_sc_hvl__buf_1.spice
* Created: Fri Aug 28 09:32:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__buf_1.pex.spice"
.subckt sky130_fd_sc_hvl__buf_1  VNB VPB A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_84_81#_M1001_g N_X_M1001_s N_VNB_M1001_b NHV L=0.5
+ W=0.75 AD=0.194904 AS=0.19875 PD=1.60256 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1002 N_A_84_81#_M1002_d N_A_M1002_g N_VGND_M1001_d N_VNB_M1001_b NHV L=0.5
+ W=0.42 AD=0.1197 AS=0.109146 PD=1.41 PS=0.897436 NRD=0 NRS=59.7132 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1000 N_VPWR_M1000_d N_A_84_81#_M1000_g N_X_M1000_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.34 AS=0.4275 PD=2.52667 PS=3.57 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
MM1003 N_A_84_81#_M1003_d N_A_M1003_g N_VPWR_M1000_d N_VPB_M1000_b PHV L=0.5
+ W=0.75 AD=0.21375 AS=0.17 PD=2.07 PS=1.26333 NRD=0 NRS=29.2803 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
DX4_noxref N_VNB_M1001_b N_VPB_M1000_b NWDIODE A=7.956 P=11.32
*
.include "sky130_fd_sc_hvl__buf_1.pxi.spice"
*
.ends
*
*
