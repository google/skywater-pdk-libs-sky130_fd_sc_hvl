* NGSPICE file created from sky130_fd_sc_hvl__inv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__inv_2 A VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB phv w=1.5e+06u l=500000u
+  ad=8.55e+11p pd=7.14e+06u as=4.2e+11p ps=3.56e+06u
M1001 Y A VGND VNB nhv w=750000u l=500000u
+  ad=2.1e+11p pd=2.06e+06u as=4.275e+11p ps=4.14e+06u
M1002 Y A VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A Y VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends

