* File: sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1.spice
* Created: Wed Sep  2 09:08:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1.pex.spice"
.subckt sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1  VNB VPB LVPWR A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* LVPWR	LVPWR
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_A_M1015_g N_A_573_897#_M1015_s N_VNB_M1015_b NSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2478 PD=1.12 PS=2.27 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1016 N_A_772_151#_M1016_d N_A_573_897#_M1016_g N_VGND_M1015_d N_VNB_M1015_b
+ NSHORT L=0.15 W=0.84 AD=0.2478 AS=0.1176 PD=2.27 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A_573_897#_M1001_g N_A_816_1221#_M1001_s N_VNB_M1015_b
+ NHV L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 M=1 R=3
+ SA=250000 SB=250001 A=0.75 P=4 MULT=1
MM1004 N_VGND_M1004_d N_A_573_897#_M1004_g N_A_816_1221#_M1001_s N_VNB_M1015_b
+ NHV L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 M=1 R=3
+ SA=250001 SB=250000 A=0.75 P=4 MULT=1
MM1000 N_A_1197_107#_M1000_d N_A_772_151#_M1000_g N_VGND_M1000_s N_VNB_M1015_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 M=1 R=3
+ SA=250000 SB=250001 A=0.75 P=4 MULT=1
MM1012 N_A_1197_107#_M1000_d N_A_772_151#_M1012_g N_VGND_M1012_s N_VNB_M1015_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 M=1 R=3
+ SA=250001 SB=250000 A=0.75 P=4 MULT=1
MM1010 N_A_1197_107#_M1010_d N_A_1406_429#_M1010_g N_A_1400_777#_M1010_s
+ N_VNB_M1015_b NHV L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0
+ M=1 R=3 SA=250000 SB=250001 A=0.75 P=4 MULT=1
MM1018 N_A_1197_107#_M1018_d N_A_1406_429#_M1018_g N_A_1400_777#_M1010_s
+ N_VNB_M1015_b NHV L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0
+ M=1 R=3 SA=250001 SB=250000 A=0.75 P=4 MULT=1
MM1011 N_VGND_M1011_d N_A_816_1221#_M1011_g N_A_1406_429#_M1011_s N_VNB_M1015_b
+ NHV L=0.5 W=0.75 AD=0.121875 AS=0.19875 PD=1.075 PS=2.03 NRD=6.8286 NRS=0 M=1
+ R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1007 N_X_M1007_d N_A_1406_429#_M1007_g N_VGND_M1011_d N_VNB_M1015_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.121875 PD=2.03 PS=1.075 NRD=0 NRS=0 M=1 R=1.5 SA=250001
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1005 N_LVPWR_M1005_d N_A_M1005_g N_A_573_897#_M1005_s N_LVPWR_M1005_b PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2478 PD=1.12 PS=2.27 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1017 N_A_772_151#_M1017_d N_A_573_897#_M1017_g N_LVPWR_M1005_d N_LVPWR_M1005_b
+ PHIGHVT L=0.15 W=0.84 AD=0.2478 AS=0.1176 PD=2.27 PS=1.12 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_A_1400_777#_M1008_g N_A_816_1221#_M1008_s N_VPB_M1008_b
+ PHV L=0.5 W=1.5 AD=0.24375 AS=0.3975 PD=1.825 PS=3.53 NRD=5.7109 NRS=0 M=1 R=3
+ SA=250000 SB=250001 A=0.75 P=4 MULT=1
MM13_noxref N_VPWR_M13_noxref_d N_A_1406_429#_M13_noxref_g
+ N_A_816_1221#_M13_noxref_s N_VPB_M1008_b PHV L=1 W=0.42 AD=0.12285 AS=0.2142
+ PD=1.07 PS=1.99 NRD=37.5124 NRS=37.5124 M=1 R=0.42 SA=500000 SB=500002 A=0.42
+ P=2.84 MULT=1
MM1009 N_VPWR_M1008_d N_A_1400_777#_M1009_g N_A_816_1221#_M1009_s N_VPB_M1008_b
+ PHV L=0.5 W=1.5 AD=0.24375 AS=0.3975 PD=1.825 PS=3.53 NRD=0 NRS=0 M=1 R=3
+ SA=250001 SB=250000 A=0.75 P=4 MULT=1
MM15_noxref N_A_1400_777#_M15_noxref_d N_A_816_1221#_M15_noxref_g
+ N_VPWR_M13_noxref_d N_VPB_M1008_b PHV L=1 W=0.42 AD=0.12285 AS=0.12285 PD=1.07
+ PS=1.07 NRD=37.5124 NRS=37.5124 M=1 R=0.42 SA=500001 SB=500001 A=0.42 P=2.84
+ MULT=1
MM1013 N_VPWR_M1013_d N_A_816_1221#_M1013_g N_A_1406_429#_M1013_s N_VPB_M1008_b
+ PHV L=0.5 W=1.5 AD=0.24375 AS=0.3975 PD=1.825 PS=3.53 NRD=5.7109 NRS=0 M=1 R=3
+ SA=250000 SB=250001 A=0.75 P=4 MULT=1
MM17_noxref N_VPWR_M17_noxref_d N_A_1406_429#_M17_noxref_g
+ N_A_1400_777#_M15_noxref_d N_VPB_M1008_b PHV L=0.5 W=0.42 AD=0.2142 AS=0.12285
+ PD=1.99 PS=1.07 NRD=37.5124 NRS=37.5124 M=1 R=0.84 SA=250003 SB=250000 A=0.21
+ P=1.84 MULT=1
MM1014 N_X_M1014_d N_A_1406_429#_M1014_g N_VPWR_M1013_d N_VPB_M1008_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.24375 PD=3.53 PS=1.825 NRD=0 NRS=0 M=1 R=3 SA=250001
+ SB=250000 A=0.75 P=4 MULT=1
DX19_noxref N_VNB_M1015_b N_VPB_X19_noxref_D1 NWDIODE A=4.9381 P=11
DX20_noxref N_VNB_M1015_b N_LVPWR_M1005_b NWDIODE A=3.54585 P=7.69
DX21_noxref N_VNB_M1015_b N_VPB_M1008_b NWDIODE A=19.9932 P=18.81
*
.include "sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1.pxi.spice"
*
.ends
*
*
