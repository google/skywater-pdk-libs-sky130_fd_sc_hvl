# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__a22oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__a22oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.505000 2.755000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.940000 1.505000 3.715000 1.750000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.505000 1.795000 1.750000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.505000 0.835000 1.835000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.630000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.925000 2.175000 1.285000 3.455000 ;
        RECT 1.085000 0.810000 1.955000 0.980000 ;
        RECT 1.085000 0.980000 1.285000 2.175000 ;
        RECT 1.705000 0.495000 1.955000 0.810000 ;
        RECT 1.705000 0.980000 1.955000 1.325000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.840000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.840000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.840000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.840000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.985000 3.840000 4.155000 ;
      RECT 0.090000  0.365000 0.680000 1.325000 ;
      RECT 0.145000  2.175000 0.475000 3.635000 ;
      RECT 0.145000  3.635000 1.955000 3.805000 ;
      RECT 1.705000  1.930000 3.595000 2.100000 ;
      RECT 1.705000  2.100000 1.955000 3.635000 ;
      RECT 2.135000  0.365000 3.750000 1.325000 ;
      RECT 2.135000  2.280000 3.085000 3.755000 ;
      RECT 3.265000  2.100000 3.595000 3.755000 ;
    LAYER mcon ;
      RECT 0.120000  0.395000 0.290000 0.565000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.480000  0.395000 0.650000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.135000  0.395000 2.305000 0.565000 ;
      RECT 2.165000  3.505000 2.335000 3.675000 ;
      RECT 2.495000  0.395000 2.665000 0.565000 ;
      RECT 2.525000  3.505000 2.695000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.855000  0.395000 3.025000 0.565000 ;
      RECT 2.885000  3.505000 3.055000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.215000  0.395000 3.385000 0.565000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.575000  0.395000 3.745000 0.565000 ;
  END
END sky130_fd_sc_hvl__a22oi_1
END LIBRARY
