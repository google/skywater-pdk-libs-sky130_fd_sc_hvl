* File: sky130_fd_sc_hvl__dfsbp_1.pex.spice
* Created: Wed Sep  2 09:05:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%VNB 5 7 11
c129 5 0 8.57047e-20 $X=-0.33 $Y=-0.265
r130 7 11 0.000401182 $w=1.776e-05 $l=5.7e-08 $layer=MET1_cond $X=8.88 $Y=0.057
+ $X2=8.88 $Y2=0
r131 5 11 0.502703 $w=1.7e-07 $l=3.145e-06 $layer=mcon $count=18 $X=17.52 $Y=0
+ $X2=17.52 $Y2=0
r132 5 11 0.502703 $w=1.7e-07 $l=3.145e-06 $layer=mcon $count=18 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%VPB 4 6 14
r148 10 14 0.502703 $w=1.7e-07 $l=3.145e-06 $layer=mcon $count=18 $X=17.52
+ $Y=4.07 $X2=17.52 $Y2=4.07
r149 9 14 1127.36 $w=1.68e-07 $l=1.728e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=17.52 $Y2=4.07
r150 9 10 0.502703 $w=1.7e-07 $l=3.145e-06 $layer=mcon $count=18 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r151 6 10 0.000401182 $w=1.776e-05 $l=5.7e-08 $layer=MET1_cond $X=8.88 $Y=4.013
+ $X2=8.88 $Y2=4.07
r152 4 14 9.83784 $w=1.7e-07 $l=1.75624e-05 $layer=licon1_NTAP_notbjt $count=18
+ $X=0 $Y=3.985 $X2=17.52 $Y2=4.07
r153 4 9 9.83784 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=18
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%CLK 3 7 9 10 11 16
r30 16 19 54.0174 $w=5.2e-07 $l=5.25e-07 $layer=POLY_cond $X=0.675 $Y=1.795
+ $X2=0.675 $Y2=2.32
r31 16 18 19.0347 $w=5.2e-07 $l=1.85e-07 $layer=POLY_cond $X=0.675 $Y=1.795
+ $X2=0.675 $Y2=1.61
r32 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.725
+ $Y=1.795 $X2=0.725 $Y2=1.795
r33 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.725 $Y=2.035
+ $X2=0.725 $Y2=2.405
r34 10 17 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.725 $Y=2.035
+ $X2=0.725 $Y2=1.795
r35 9 17 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.725 $Y=1.665
+ $X2=0.725 $Y2=1.795
r36 7 19 76.5092 $w=5e-07 $l=7.15e-07 $layer=POLY_cond $X=0.685 $Y=3.035
+ $X2=0.685 $Y2=2.32
r37 3 18 89.8849 $w=5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.665 $Y=0.77 $X2=0.665
+ $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%A_30_112# 1 2 9 13 17 18 20 23 27 30 34 36
+ 38 39 41 42 43 45 46 47 49 50 51 54 55 58 59 60 61 64 65 66 68 69 70 72 73 74
+ 77 78 80 83 88 97 103
c266 65 0 1.25957e-19 $X=6.425 $Y=2.64
c267 55 0 1.42106e-19 $X=3.64 $Y=1.27
r268 92 93 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.695
+ $Y=2.39 $X2=4.695 $Y2=2.39
r269 85 87 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.64 $Y=2.31
+ $X2=3.81 $Y2=2.31
r270 83 101 54.0174 $w=5.2e-07 $l=5.25e-07 $layer=POLY_cond $X=1.455 $Y=1.365
+ $X2=1.455 $Y2=1.89
r271 83 100 26.237 $w=5.2e-07 $l=2.55e-07 $layer=POLY_cond $X=1.455 $Y=1.365
+ $X2=1.455 $Y2=1.11
r272 82 83 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.425
+ $Y=1.365 $X2=1.425 $Y2=1.365
r273 78 97 124.662 $w=5e-07 $l=1.165e-06 $layer=POLY_cond $X=9.12 $Y=2.05
+ $X2=9.12 $Y2=3.215
r274 77 78 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.035
+ $Y=2.05 $X2=9.035 $Y2=2.05
r275 75 77 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=8.995 $Y=2.545
+ $X2=8.995 $Y2=2.05
r276 73 75 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.87 $Y=2.63
+ $X2=8.995 $Y2=2.545
r277 73 74 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=8.87 $Y=2.63
+ $X2=7.675 $Y2=2.63
r278 71 74 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.59 $Y=2.715
+ $X2=7.675 $Y2=2.63
r279 71 72 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=7.59 $Y=2.715
+ $X2=7.59 $Y2=3.355
r280 69 72 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.505 $Y=3.44
+ $X2=7.59 $Y2=3.355
r281 69 70 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=7.505 $Y=3.44
+ $X2=6.595 $Y2=3.44
r282 68 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.51 $Y=3.355
+ $X2=6.595 $Y2=3.44
r283 67 68 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=6.51 $Y=2.725
+ $X2=6.51 $Y2=3.355
r284 65 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.425 $Y=2.64
+ $X2=6.51 $Y2=2.725
r285 65 66 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=6.425 $Y=2.64
+ $X2=5.5 $Y2=2.64
r286 63 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.415 $Y=2.725
+ $X2=5.5 $Y2=2.64
r287 63 64 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.415 $Y=2.725
+ $X2=5.415 $Y2=3.355
r288 62 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=3.44
+ $X2=3.81 $Y2=3.44
r289 61 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.33 $Y=3.44
+ $X2=5.415 $Y2=3.355
r290 61 62 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=5.33 $Y=3.44
+ $X2=3.895 $Y2=3.44
r291 60 87 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=2.31
+ $X2=3.81 $Y2=2.31
r292 59 92 4.28816 $w=2.13e-07 $l=8e-08 $layer=LI1_cond $X=4.692 $Y=2.31
+ $X2=4.692 $Y2=2.39
r293 59 60 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.585 $Y=2.31
+ $X2=3.895 $Y2=2.31
r294 58 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=3.355
+ $X2=3.81 $Y2=3.44
r295 57 87 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=2.395
+ $X2=3.81 $Y2=2.31
r296 57 58 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.81 $Y=2.395
+ $X2=3.81 $Y2=3.355
r297 55 103 19.0347 $w=5.2e-07 $l=1.85e-07 $layer=POLY_cond $X=3.565 $Y=1.27
+ $X2=3.565 $Y2=1.085
r298 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.64
+ $Y=1.27 $X2=3.64 $Y2=1.27
r299 52 85 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=2.225
+ $X2=3.64 $Y2=2.31
r300 52 54 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.64 $Y=2.225
+ $X2=3.64 $Y2=1.27
r301 50 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=3.44
+ $X2=3.81 $Y2=3.44
r302 50 51 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.725 $Y=3.44
+ $X2=3.025 $Y2=3.44
r303 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.94 $Y=3.355
+ $X2=3.025 $Y2=3.44
r304 48 49 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.94 $Y=2.495
+ $X2=2.94 $Y2=3.355
r305 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.855 $Y=2.41
+ $X2=2.94 $Y2=2.495
r306 46 47 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.855 $Y=2.41
+ $X2=2.29 $Y2=2.41
r307 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.205 $Y=2.495
+ $X2=2.29 $Y2=2.41
r308 44 45 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=2.205 $Y=2.495
+ $X2=2.205 $Y2=3.63
r309 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.12 $Y=3.715
+ $X2=2.205 $Y2=3.63
r310 42 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.12 $Y=3.715
+ $X2=1.59 $Y2=3.715
r311 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=3.63
+ $X2=1.59 $Y2=3.715
r312 41 84 114.824 $w=1.68e-07 $l=1.76e-06 $layer=LI1_cond $X=1.505 $Y=3.63
+ $X2=1.505 $Y2=1.87
r313 39 84 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=1.705
+ $X2=1.425 $Y2=1.87
r314 38 82 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.425 $Y=1.37
+ $X2=1.425 $Y2=1.285
r315 38 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.425 $Y=1.37
+ $X2=1.425 $Y2=1.705
r316 37 80 2.90867 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.38 $Y=1.285
+ $X2=0.245 $Y2=1.285
r317 36 82 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.26 $Y=1.285
+ $X2=1.425 $Y2=1.285
r318 36 37 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=1.26 $Y=1.285
+ $X2=0.38 $Y2=1.285
r319 32 80 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=1.37
+ $X2=0.245 $Y2=1.285
r320 32 34 60.3965 $w=2.68e-07 $l=1.415e-06 $layer=LI1_cond $X=0.245 $Y=1.37
+ $X2=0.245 $Y2=2.785
r321 28 80 3.58051 $w=2.6e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.235 $Y=1.2
+ $X2=0.245 $Y2=1.285
r322 28 30 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.235 $Y=1.2
+ $X2=0.235 $Y2=0.77
r323 27 78 25.1464 $w=5e-07 $l=2.35e-07 $layer=POLY_cond $X=9.12 $Y=1.815
+ $X2=9.12 $Y2=2.05
r324 26 27 37.2588 $w=6.9e-07 $l=5e-07 $layer=POLY_cond $X=9.215 $Y=1.315
+ $X2=9.215 $Y2=1.815
r325 23 26 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=9.31 $Y=0.975 $X2=9.31
+ $Y2=1.315
r326 18 93 26.3136 $w=5e-07 $l=2.65e-07 $layer=POLY_cond $X=4.63 $Y=2.655
+ $X2=4.63 $Y2=2.39
r327 18 20 26.028 $w=5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.63 $Y=2.655 $X2=4.63
+ $Y2=2.925
r328 17 103 31.812 $w=5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.555 $Y=0.755
+ $X2=3.555 $Y2=1.085
r329 13 101 122.522 $w=5e-07 $l=1.145e-06 $layer=POLY_cond $X=1.465 $Y=3.035
+ $X2=1.465 $Y2=1.89
r330 9 100 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.445 $Y=0.77
+ $X2=1.445 $Y2=1.11
r331 2 34 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.66 $X2=0.295 $Y2=2.785
r332 1 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.56 $X2=0.275 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%D 3 8 10 11 15
r42 15 18 96.8403 $w=5e-07 $l=9.05e-07 $layer=POLY_cond $X=2.775 $Y=0.755
+ $X2=2.775 $Y2=1.66
r43 10 11 12.3476 $w=3.48e-07 $l=3.75e-07 $layer=LI1_cond $X=2.7 $Y=1.66 $X2=2.7
+ $Y2=2.035
r44 10 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.71
+ $Y=1.66 $X2=2.71 $Y2=1.66
r45 6 18 45.4775 $w=5e-07 $l=4.25e-07 $layer=POLY_cond $X=2.775 $Y=2.085
+ $X2=2.775 $Y2=1.66
r46 5 8 31.5667 $w=5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.775 $Y=2.335 $X2=3.07
+ $Y2=2.335
r47 5 6 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.775 $Y=2.335 $X2=2.775
+ $Y2=2.085
r48 1 8 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.07 $Y=2.585 $X2=3.07
+ $Y2=2.335
r49 1 3 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.07 $Y=2.585 $X2=3.07
+ $Y2=2.925
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%A_339_112# 1 2 7 9 13 17 23 26 28 31 32 33
+ 38 39 41 43 45 48 50 52 54 56 59 65
c180 54 0 8.42554e-20 $X=10.02 $Y=2.39
c181 32 0 2.67476e-20 $X=4.29 $Y=0.35
c182 28 0 1.42106e-19 $X=2.65 $Y=1.25
c183 9 0 3.21706e-20 $X=3.85 $Y=2.925
r184 55 65 32.1018 $w=5e-07 $l=3e-07 $layer=POLY_cond $X=10.02 $Y=2.335
+ $X2=10.32 $Y2=2.335
r185 55 62 0.535029 $w=5e-07 $l=5e-09 $layer=POLY_cond $X=10.02 $Y=2.335
+ $X2=10.015 $Y2=2.335
r186 54 56 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=10.02 $Y=2.43
+ $X2=9.855 $Y2=2.43
r187 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.02
+ $Y=2.39 $X2=10.02 $Y2=2.39
r188 51 59 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.335 $Y=1.24
+ $X2=4.335 $Y2=0.755
r189 50 52 7.4145 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=4.42 $Y=1.24
+ $X2=4.42 $Y2=1.105
r190 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.42
+ $Y=1.24 $X2=4.42 $Y2=1.24
r191 45 47 9.10257 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.835 $Y=0.77
+ $X2=1.835 $Y2=1
r192 43 56 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.47 $Y=2.39
+ $X2=9.855 $Y2=2.39
r193 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.385 $Y=2.305
+ $X2=9.47 $Y2=2.39
r194 40 41 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=9.385 $Y=1.675
+ $X2=9.385 $Y2=2.305
r195 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.3 $Y=1.59
+ $X2=9.385 $Y2=1.675
r196 38 39 307.61 $w=1.68e-07 $l=4.715e-06 $layer=LI1_cond $X=9.3 $Y=1.59
+ $X2=4.585 $Y2=1.59
r197 36 52 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.375 $Y=0.435
+ $X2=4.375 $Y2=1.105
r198 35 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.42 $Y=1.505
+ $X2=4.585 $Y2=1.59
r199 34 50 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=4.42 $Y=1.27 $X2=4.42
+ $Y2=1.24
r200 34 35 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.42 $Y=1.27
+ $X2=4.42 $Y2=1.505
r201 32 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.29 $Y=0.35
+ $X2=4.375 $Y2=0.435
r202 32 33 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=4.29 $Y=0.35
+ $X2=2.82 $Y2=0.35
r203 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.735 $Y=0.435
+ $X2=2.82 $Y2=0.35
r204 30 31 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.735 $Y=0.435
+ $X2=2.735 $Y2=1.165
r205 29 48 1.93381 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2 $Y=1.25 $X2=1.885
+ $Y2=1.25
r206 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.65 $Y=1.25
+ $X2=2.735 $Y2=1.165
r207 28 29 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.65 $Y=1.25 $X2=2
+ $Y2=1.25
r208 24 48 4.50329 $w=2e-07 $l=9.88686e-08 $layer=LI1_cond $X=1.855 $Y=1.335
+ $X2=1.885 $Y2=1.25
r209 24 26 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=1.855 $Y=1.335
+ $X2=1.855 $Y2=2.785
r210 23 48 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.885 $Y=1.165
+ $X2=1.885 $Y2=1.25
r211 23 47 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=1.165
+ $X2=1.885 $Y2=1
r212 21 51 24.0763 $w=5e-07 $l=2.25e-07 $layer=POLY_cond $X=4.335 $Y=1.465
+ $X2=4.335 $Y2=1.24
r213 15 65 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=10.32 $Y=2.085
+ $X2=10.32 $Y2=2.335
r214 15 17 101.121 $w=5e-07 $l=9.45e-07 $layer=POLY_cond $X=10.32 $Y=2.085
+ $X2=10.32 $Y2=1.14
r215 11 62 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=10.015 $Y=2.585
+ $X2=10.015 $Y2=2.335
r216 11 13 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=10.015 $Y=2.585
+ $X2=10.015 $Y2=2.925
r217 7 21 53.3721 $w=4.38e-07 $l=6.42067e-07 $layer=POLY_cond $X=3.85 $Y=2.195
+ $X2=4.335 $Y2=1.83
r218 7 9 78.1143 $w=5e-07 $l=7.3e-07 $layer=POLY_cond $X=3.85 $Y=2.195 $X2=3.85
+ $Y2=2.925
r219 2 26 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.715
+ $Y=2.66 $X2=1.855 $Y2=2.785
r220 1 45 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.56 $X2=1.835 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%A_959_83# 1 2 7 9 14 16 21 24 28 32 37 40
c78 32 0 8.57047e-20 $X=6.86 $Y=2.925
c79 7 0 2.67476e-20 $X=5.045 $Y=1.075
r80 30 32 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=6.9 $Y=2.375 $X2=6.9
+ $Y2=2.925
r81 26 28 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.985 $Y=1.085
+ $X2=5.985 $Y2=0.745
r82 24 41 28.1508 $w=5.9e-07 $l=2.95e-07 $layer=POLY_cond $X=5.385 $Y=2.29
+ $X2=5.385 $Y2=2.585
r83 24 40 19.9893 $w=5.9e-07 $l=2.05e-07 $layer=POLY_cond $X=5.385 $Y=2.29
+ $X2=5.385 $Y2=2.085
r84 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.495
+ $Y=2.29 $X2=5.495 $Y2=2.29
r85 21 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.775 $Y=2.29
+ $X2=6.9 $Y2=2.375
r86 21 23 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=6.775 $Y=2.29
+ $X2=5.495 $Y2=2.29
r87 19 37 24.6114 $w=5e-07 $l=2.3e-07 $layer=POLY_cond $X=5.11 $Y=1.325 $X2=5.34
+ $Y2=1.325
r88 19 34 6.95538 $w=5e-07 $l=6.5e-08 $layer=POLY_cond $X=5.11 $Y=1.325
+ $X2=5.045 $Y2=1.325
r89 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.11
+ $Y=1.24 $X2=5.11 $Y2=1.24
r90 16 26 7.03987 $w=2.4e-07 $l=2.16852e-07 $layer=LI1_cond $X=5.82 $Y=1.205
+ $X2=5.985 $Y2=1.085
r91 16 18 34.0931 $w=2.38e-07 $l=7.1e-07 $layer=LI1_cond $X=5.82 $Y=1.205
+ $X2=5.11 $Y2=1.205
r92 14 41 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.34 $Y=2.925 $X2=5.34
+ $Y2=2.585
r93 10 37 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.34 $Y=1.575 $X2=5.34
+ $Y2=1.325
r94 10 40 54.573 $w=5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.34 $Y=1.575 $X2=5.34
+ $Y2=2.085
r95 7 34 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.045 $Y=1.075
+ $X2=5.045 $Y2=1.325
r96 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.045 $Y=1.075 $X2=5.045
+ $Y2=0.755
r97 2 32 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.72
+ $Y=2.715 $X2=6.86 $Y2=2.925
r98 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.86
+ $Y=0.535 $X2=5.985 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%A_761_109# 1 2 9 13 17 21 24 25 26 27 30 31
+ 35 36 38 42 46 50 60
c139 27 0 3.21706e-20 $X=4.98 $Y=3.09
r140 59 60 27.8768 $w=8.3e-07 $l=4.5e-07 $layer=POLY_cond $X=7.96 $Y=2.17
+ $X2=8.41 $Y2=2.17
r141 53 59 4.02665 $w=8.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.895 $Y=2.17
+ $X2=7.96 $Y2=2.17
r142 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.895
+ $Y=1.94 $X2=7.895 $Y2=1.94
r143 46 48 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.24 $Y=2.925
+ $X2=4.24 $Y2=3.09
r144 42 44 8.11295 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.945 $Y=0.77
+ $X2=3.945 $Y2=0.925
r145 38 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.895
+ $Y=2.28 $X2=7.895 $Y2=2.28
r146 36 52 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.895 $Y=2.025
+ $X2=7.895 $Y2=1.94
r147 36 38 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.895 $Y=2.025
+ $X2=7.895 $Y2=2.28
r148 35 56 29.8454 $w=5.95e-07 $l=3.15e-07 $layer=POLY_cond $X=6.422 $Y=1.94
+ $X2=6.422 $Y2=2.255
r149 35 55 18.1557 $w=5.95e-07 $l=1.85e-07 $layer=POLY_cond $X=6.422 $Y=1.94
+ $X2=6.422 $Y2=1.755
r150 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.31
+ $Y=1.94 $X2=6.31 $Y2=1.94
r151 32 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=1.94
+ $X2=5.065 $Y2=1.94
r152 32 34 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=5.15 $Y=1.94
+ $X2=6.31 $Y2=1.94
r153 31 52 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.73 $Y=1.94
+ $X2=7.895 $Y2=1.94
r154 31 34 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=7.73 $Y=1.94
+ $X2=6.31 $Y2=1.94
r155 29 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=2.025
+ $X2=5.065 $Y2=1.94
r156 29 30 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=5.065 $Y=2.025
+ $X2=5.065 $Y2=3.005
r157 28 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=3.09
+ $X2=4.24 $Y2=3.09
r158 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.98 $Y=3.09
+ $X2=5.065 $Y2=3.005
r159 27 28 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.98 $Y=3.09
+ $X2=4.405 $Y2=3.09
r160 25 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=1.94
+ $X2=5.065 $Y2=1.94
r161 25 26 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=4.98 $Y=1.94
+ $X2=4.075 $Y2=1.94
r162 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.99 $Y=1.855
+ $X2=4.075 $Y2=1.94
r163 24 44 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.99 $Y=1.855
+ $X2=3.99 $Y2=0.925
r164 19 60 14.627 $w=5e-07 $l=4.15e-07 $layer=POLY_cond $X=8.41 $Y=2.585
+ $X2=8.41 $Y2=2.17
r165 19 21 67.4137 $w=5e-07 $l=6.3e-07 $layer=POLY_cond $X=8.41 $Y=2.585
+ $X2=8.41 $Y2=3.215
r166 15 59 14.627 $w=5e-07 $l=4.15e-07 $layer=POLY_cond $X=7.96 $Y=1.755
+ $X2=7.96 $Y2=2.17
r167 15 17 90.42 $w=5e-07 $l=8.45e-07 $layer=POLY_cond $X=7.96 $Y=1.755 $X2=7.96
+ $Y2=0.91
r168 13 56 71.6939 $w=5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.47 $Y=2.925
+ $X2=6.47 $Y2=2.255
r169 9 55 108.076 $w=5e-07 $l=1.01e-06 $layer=POLY_cond $X=6.375 $Y=0.745
+ $X2=6.375 $Y2=1.755
r170 2 46 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.1
+ $Y=2.715 $X2=4.24 $Y2=2.925
r171 1 42 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=3.805
+ $Y=0.545 $X2=3.945 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%SET_B 1 3 4 5 8 11 13 16 19 25 26 27 29 31
+ 32 33 37 44
c114 13 0 1.25957e-19 $X=7.215 $Y=2.605
r115 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.53
+ $Y=1.68 $X2=12.53 $Y2=1.68
r116 37 40 100.051 $w=5e-07 $l=9.35e-07 $layer=POLY_cond $X=12.595 $Y=0.745
+ $X2=12.595 $Y2=1.68
r117 33 41 3.85178 $w=5.88e-07 $l=1.9e-07 $layer=LI1_cond $X=12.72 $Y=1.85
+ $X2=12.53 $Y2=1.85
r118 32 41 5.87903 $w=5.88e-07 $l=2.9e-07 $layer=LI1_cond $X=12.24 $Y=1.85
+ $X2=12.53 $Y2=1.85
r119 32 44 8.57049 $w=5.88e-07 $l=9e-08 $layer=LI1_cond $X=12.24 $Y=1.85
+ $X2=12.15 $Y2=1.85
r120 31 44 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=10.885 $Y=2.06
+ $X2=12.15 $Y2=2.06
r121 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.8 $Y=1.975
+ $X2=10.885 $Y2=2.06
r122 28 29 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=10.8 $Y=1.775
+ $X2=10.8 $Y2=1.975
r123 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.715 $Y=1.69
+ $X2=10.8 $Y2=1.775
r124 26 27 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.715 $Y=1.69
+ $X2=10.33 $Y2=1.69
r125 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.245 $Y=1.605
+ $X2=10.33 $Y2=1.69
r126 24 25 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.245 $Y=1.325
+ $X2=10.245 $Y2=1.605
r127 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.15
+ $Y=1.24 $X2=7.15 $Y2=1.24
r128 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.16 $Y=1.24
+ $X2=10.245 $Y2=1.325
r129 19 21 196.374 $w=1.68e-07 $l=3.01e-06 $layer=LI1_cond $X=10.16 $Y=1.24
+ $X2=7.15 $Y2=1.24
r130 17 40 43.3374 $w=5e-07 $l=4.05e-07 $layer=POLY_cond $X=12.595 $Y=2.085
+ $X2=12.595 $Y2=1.68
r131 16 17 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=12.595 $Y=2.335
+ $X2=12.595 $Y2=2.085
r132 14 16 83.9996 $w=5e-07 $l=7.85e-07 $layer=POLY_cond $X=11.81 $Y=2.335
+ $X2=12.595 $Y2=2.335
r133 9 14 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=11.81 $Y=2.585
+ $X2=11.81 $Y2=2.335
r134 9 11 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=11.81 $Y=2.585
+ $X2=11.81 $Y2=2.925
r135 8 13 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.25 $Y=2.925 $X2=7.25
+ $Y2=2.605
r136 5 13 27.696 $w=5.7e-07 $l=2.85e-07 $layer=POLY_cond $X=7.215 $Y=2.32
+ $X2=7.215 $Y2=2.605
r137 4 22 49.8912 $w=5.7e-07 $l=6.13531e-07 $layer=POLY_cond $X=7.215 $Y=1.83
+ $X2=7.167 $Y2=1.24
r138 4 5 45.9938 $w=5.7e-07 $l=4.9e-07 $layer=POLY_cond $X=7.215 $Y=1.83
+ $X2=7.215 $Y2=2.32
r139 1 22 15.8546 $w=5.48e-07 $l=2.12073e-07 $layer=POLY_cond $X=7.085 $Y=1.065
+ $X2=7.167 $Y2=1.24
r140 1 3 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.085 $Y=1.065 $X2=7.085
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%A_2156_417# 1 2 9 13 15 17 18 21 25 29 31
+ 32 33 36 38 40
c98 18 0 1.2513e-19 $X=11.065 $Y=2.585
c99 17 0 8.21585e-20 $X=11.065 $Y=2.085
r100 39 41 38.5111 $w=7.45e-07 $l=5.58e-07 $layer=POLY_cond $X=11.805 $Y=1.457
+ $X2=11.247 $Y2=1.457
r101 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.805
+ $Y=1.305 $X2=11.805 $Y2=1.305
r102 35 36 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=14.31 $Y=1.375
+ $X2=14.31 $Y2=1.905
r103 34 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.72 $Y=1.29
+ $X2=13.555 $Y2=1.29
r104 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.225 $Y=1.29
+ $X2=14.31 $Y2=1.375
r105 33 34 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=14.225 $Y=1.29
+ $X2=13.72 $Y2=1.29
r106 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.225 $Y=1.99
+ $X2=14.31 $Y2=1.905
r107 31 32 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=14.225 $Y=1.99
+ $X2=13.69 $Y2=1.99
r108 27 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.555 $Y=1.205
+ $X2=13.555 $Y2=1.29
r109 27 29 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=13.555 $Y=1.205
+ $X2=13.555 $Y2=1.075
r110 23 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.525 $Y=2.075
+ $X2=13.69 $Y2=1.99
r111 23 25 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=13.525 $Y=2.075
+ $X2=13.525 $Y2=2.425
r112 22 38 4.91858 $w=1.7e-07 $l=1.77059e-07 $layer=LI1_cond $X=11.97 $Y=1.29
+ $X2=11.805 $Y2=1.265
r113 21 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.39 $Y=1.29
+ $X2=13.555 $Y2=1.29
r114 21 22 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=13.39 $Y=1.29
+ $X2=11.97 $Y2=1.29
r115 17 18 72.6564 $w=5e-07 $l=5e-07 $layer=POLY_cond $X=11.065 $Y=2.085
+ $X2=11.065 $Y2=2.585
r116 13 39 5.52131 $w=7.45e-07 $l=8e-08 $layer=POLY_cond $X=11.885 $Y=1.457
+ $X2=11.805 $Y2=1.457
r117 13 15 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=11.885 $Y=1.085
+ $X2=11.885 $Y2=0.745
r118 11 41 33.6369 $w=2.05e-07 $l=3.73e-07 $layer=POLY_cond $X=11.247 $Y=1.83
+ $X2=11.247 $Y2=1.457
r119 11 17 82.4899 $w=2.05e-07 $l=2.55e-07 $layer=POLY_cond $X=11.247 $Y=1.83
+ $X2=11.247 $Y2=2.085
r120 9 18 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=11.03 $Y=2.925
+ $X2=11.03 $Y2=2.585
r121 2 25 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=13.38
+ $Y=2.215 $X2=13.525 $Y2=2.425
r122 1 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=13.41
+ $Y=0.865 $X2=13.555 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%A_1874_543# 1 2 3 12 16 20 24 26 27 30 34
+ 36 41 47 49 50 51 52 54 56 59 60 62 63 65 68 71
c164 51 0 1.23033e-19 $X=10.365 $Y=2.04
r165 76 77 1.07006 $w=5e-07 $l=1e-08 $layer=POLY_cond $X=14.81 $Y=1.665
+ $X2=14.82 $Y2=1.665
r166 75 76 92.5601 $w=5e-07 $l=8.65e-07 $layer=POLY_cond $X=13.945 $Y=1.665
+ $X2=14.81 $Y2=1.665
r167 74 75 3.21018 $w=5e-07 $l=3e-08 $layer=POLY_cond $X=13.915 $Y=1.665
+ $X2=13.945 $Y2=1.665
r168 70 71 11.9721 $w=8.48e-07 $l=1.65e-07 $layer=LI1_cond $X=12.2 $Y=2.75
+ $X2=12.035 $Y2=2.75
r169 66 74 3.74521 $w=5e-07 $l=3.5e-08 $layer=POLY_cond $X=13.88 $Y=1.665
+ $X2=13.915 $Y2=1.665
r170 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.88
+ $Y=1.64 $X2=13.88 $Y2=1.64
r171 63 65 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=13.18 $Y=1.64
+ $X2=13.88 $Y2=1.64
r172 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.095 $Y=1.725
+ $X2=13.18 $Y2=1.64
r173 61 62 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=13.095 $Y=1.725
+ $X2=13.095 $Y2=2.325
r174 60 70 3.73176 $w=8.48e-07 $l=2.6e-07 $layer=LI1_cond $X=12.46 $Y=2.75
+ $X2=12.2 $Y2=2.75
r175 59 62 11.8367 $w=8.5e-07 $l=4.65564e-07 $layer=LI1_cond $X=13.01 $Y=2.75
+ $X2=13.095 $Y2=2.325
r176 59 60 7.89412 $w=8.48e-07 $l=5.5e-07 $layer=LI1_cond $X=13.01 $Y=2.75
+ $X2=12.46 $Y2=2.75
r177 58 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.535 $Y=2.41
+ $X2=10.45 $Y2=2.41
r178 58 71 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=10.535 $Y=2.41
+ $X2=12.035 $Y2=2.41
r179 55 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.45 $Y=2.495
+ $X2=10.45 $Y2=2.41
r180 55 56 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=10.45 $Y=2.495
+ $X2=10.45 $Y2=3.585
r181 54 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.45 $Y=2.325
+ $X2=10.45 $Y2=2.41
r182 53 54 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=10.45 $Y=2.125
+ $X2=10.45 $Y2=2.325
r183 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.365 $Y=2.04
+ $X2=10.45 $Y2=2.125
r184 51 52 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.365 $Y=2.04
+ $X2=9.98 $Y2=2.04
r185 49 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.365 $Y=3.67
+ $X2=10.45 $Y2=3.585
r186 49 50 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.365 $Y=3.67
+ $X2=9.675 $Y2=3.67
r187 45 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.815 $Y=1.955
+ $X2=9.98 $Y2=2.04
r188 45 47 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=9.815 $Y=1.955
+ $X2=9.815 $Y2=1.59
r189 41 44 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=9.51 $Y=2.84
+ $X2=9.51 $Y2=3.215
r190 39 50 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.51 $Y=3.585
+ $X2=9.675 $Y2=3.67
r191 39 44 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.51 $Y=3.585
+ $X2=9.51 $Y2=3.215
r192 36 38 61.7342 $w=5.2e-07 $l=6e-07 $layer=POLY_cond $X=16.19 $Y=1.665
+ $X2=16.19 $Y2=2.265
r193 36 37 25.7226 $w=5.2e-07 $l=2.5e-07 $layer=POLY_cond $X=16.19 $Y=1.665
+ $X2=16.19 $Y2=1.415
r194 34 37 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=16.2 $Y=1.075 $X2=16.2
+ $Y2=1.415
r195 30 38 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=16.18 $Y=2.77
+ $X2=16.18 $Y2=2.265
r196 27 77 26.7515 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=15.07 $Y=1.665
+ $X2=14.82 $Y2=1.665
r197 26 36 3.77112 $w=5e-07 $l=2.6e-07 $layer=POLY_cond $X=15.93 $Y=1.665
+ $X2=16.19 $Y2=1.665
r198 26 27 92.0251 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=15.93 $Y=1.665
+ $X2=15.07 $Y2=1.665
r199 22 77 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=14.82 $Y=1.415
+ $X2=14.82 $Y2=1.665
r200 22 24 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=14.82 $Y=1.415
+ $X2=14.82 $Y2=0.91
r201 18 76 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=14.81 $Y=1.915
+ $X2=14.81 $Y2=1.665
r202 18 20 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=14.81 $Y=1.915
+ $X2=14.81 $Y2=2.965
r203 14 75 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=13.945 $Y=1.415
+ $X2=13.945 $Y2=1.665
r204 14 16 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=13.945 $Y=1.415
+ $X2=13.945 $Y2=1.075
r205 10 74 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=13.915 $Y=1.915
+ $X2=13.915 $Y2=1.665
r206 10 12 54.573 $w=5e-07 $l=5.1e-07 $layer=POLY_cond $X=13.915 $Y=1.915
+ $X2=13.915 $Y2=2.425
r207 3 70 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=12.06
+ $Y=2.715 $X2=12.2 $Y2=2.925
r208 2 44 300 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_PDIFF $count=2 $X=9.37
+ $Y=2.715 $X2=9.51 $Y2=3.215
r209 2 41 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=9.37
+ $Y=2.715 $X2=9.51 $Y2=2.84
r210 1 47 182 $w=1.7e-07 $l=9.43928e-07 $layer=licon1_NDIFF $count=1 $X=9.56
+ $Y=0.765 $X2=9.815 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%A_3129_479# 1 2 9 13 15 19 21 24 28
r41 22 28 131.082 $w=5e-07 $l=1.225e-06 $layer=POLY_cond $X=17.075 $Y=1.67
+ $X2=17.075 $Y2=2.895
r42 22 24 81.3245 $w=5e-07 $l=7.6e-07 $layer=POLY_cond $X=17.075 $Y=1.67
+ $X2=17.075 $Y2=0.91
r43 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=17.01
+ $Y=1.67 $X2=17.01 $Y2=1.67
r44 16 19 3.9231 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=15.975 $Y=1.59
+ $X2=15.8 $Y2=1.59
r45 15 21 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.845 $Y=1.59
+ $X2=17.01 $Y2=1.59
r46 15 16 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=16.845 $Y=1.59
+ $X2=15.975 $Y2=1.59
r47 11 19 2.80976 $w=3.4e-07 $l=8.9861e-08 $layer=LI1_cond $X=15.79 $Y=1.675
+ $X2=15.8 $Y2=1.59
r48 11 13 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=15.79 $Y=1.675
+ $X2=15.79 $Y2=2.52
r49 7 19 2.80976 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=15.8 $Y=1.505 $X2=15.8
+ $Y2=1.59
r50 7 9 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=15.8 $Y=1.505 $X2=15.8
+ $Y2=1.075
r51 2 13 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=15.645
+ $Y=2.395 $X2=15.79 $Y2=2.52
r52 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=15.665
+ $Y=0.865 $X2=15.81 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%VPWR 1 2 3 4 5 6 7 22 25 32 39 46 55 64 76
+ 84
r113 82 84 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=16.25 $Y=3.63
+ $X2=16.97 $Y2=3.63
r114 81 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.97 $Y=3.59
+ $X2=16.97 $Y2=3.59
r115 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.25 $Y=3.59
+ $X2=16.25 $Y2=3.59
r116 79 81 4.10947 $w=9.48e-07 $l=3.2e-07 $layer=LI1_cond $X=16.61 $Y=3.27
+ $X2=16.61 $Y2=3.59
r117 76 79 9.63158 $w=9.48e-07 $l=7.5e-07 $layer=LI1_cond $X=16.61 $Y=2.52
+ $X2=16.61 $Y2=3.27
r118 73 82 0.593134 $w=3.7e-07 $l=1.545e-06 $layer=MET1_cond $X=14.705 $Y=3.63
+ $X2=16.25 $Y2=3.63
r119 70 73 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=13.985 $Y=3.63
+ $X2=14.705 $Y2=3.63
r120 69 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.705 $Y=3.59
+ $X2=14.705 $Y2=3.59
r121 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.985 $Y=3.59
+ $X2=13.985 $Y2=3.59
r122 67 69 10.7232 $w=9.48e-07 $l=8.35e-07 $layer=LI1_cond $X=14.345 $Y=2.755
+ $X2=14.345 $Y2=3.59
r123 64 67 5.32947 $w=9.48e-07 $l=4.15e-07 $layer=LI1_cond $X=14.345 $Y=2.34
+ $X2=14.345 $Y2=2.755
r124 61 70 0.93481 $w=3.7e-07 $l=2.435e-06 $layer=MET1_cond $X=11.55 $Y=3.63
+ $X2=13.985 $Y2=3.63
r125 59 61 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.83 $Y=3.63
+ $X2=11.55 $Y2=3.63
r126 58 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.55 $Y=3.59
+ $X2=11.55 $Y2=3.59
r127 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.83 $Y=3.59
+ $X2=10.83 $Y2=3.59
r128 55 58 8.54 $w=9.48e-07 $l=6.65e-07 $layer=LI1_cond $X=11.19 $Y=2.925
+ $X2=11.19 $Y2=3.59
r129 50 52 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.97 $Y=3.63
+ $X2=8.69 $Y2=3.63
r130 49 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.69 $Y=3.59
+ $X2=8.69 $Y2=3.59
r131 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.97 $Y=3.59
+ $X2=7.97 $Y2=3.59
r132 46 49 7.64105 $w=9.48e-07 $l=5.95e-07 $layer=LI1_cond $X=8.33 $Y=2.995
+ $X2=8.33 $Y2=3.59
r133 43 50 0.702547 $w=3.7e-07 $l=1.83e-06 $layer=MET1_cond $X=6.14 $Y=3.63
+ $X2=7.97 $Y2=3.63
r134 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.14 $Y=3.59
+ $X2=6.14 $Y2=3.59
r135 39 42 12.49 $w=5.63e-07 $l=5.9e-07 $layer=LI1_cond $X=5.962 $Y=3 $X2=5.962
+ $Y2=3.59
r136 36 43 1.36862 $w=3.7e-07 $l=3.565e-06 $layer=MET1_cond $X=2.575 $Y=3.63
+ $X2=6.14 $Y2=3.63
r137 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.575 $Y=3.59
+ $X2=2.575 $Y2=3.59
r138 32 35 35.9778 $w=2.03e-07 $l=6.65e-07 $layer=LI1_cond $X=2.572 $Y=2.925
+ $X2=2.572 $Y2=3.59
r139 29 36 0.556663 $w=3.7e-07 $l=1.45e-06 $layer=MET1_cond $X=1.125 $Y=3.63
+ $X2=2.575 $Y2=3.63
r140 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.125 $Y=3.59
+ $X2=1.125 $Y2=3.59
r141 25 28 16.3194 $w=5.88e-07 $l=8.05e-07 $layer=LI1_cond $X=0.945 $Y=2.785
+ $X2=0.945 $Y2=3.59
r142 22 59 0.748616 $w=3.7e-07 $l=1.95e-06 $layer=MET1_cond $X=8.88 $Y=3.63
+ $X2=10.83 $Y2=3.63
r143 22 52 0.072942 $w=3.7e-07 $l=1.9e-07 $layer=MET1_cond $X=8.88 $Y=3.63
+ $X2=8.69 $Y2=3.63
r144 7 79 600 $w=1.7e-07 $l=9.94359e-07 $layer=licon1_PDIFF $count=1 $X=16.43
+ $Y=2.395 $X2=16.685 $Y2=3.27
r145 7 76 300 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=2 $X=16.43
+ $Y=2.395 $X2=16.685 $Y2=2.52
r146 6 69 400 $w=1.7e-07 $l=1.49708e-06 $layer=licon1_PDIFF $count=1 $X=14.165
+ $Y=2.215 $X2=14.42 $Y2=3.59
r147 6 67 400 $w=1.7e-07 $l=6.5521e-07 $layer=licon1_PDIFF $count=1 $X=14.165
+ $Y=2.215 $X2=14.42 $Y2=2.755
r148 6 64 600 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=1 $X=14.165
+ $Y=2.215 $X2=14.42 $Y2=2.34
r149 5 55 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.28
+ $Y=2.715 $X2=11.42 $Y2=2.925
r150 4 46 600 $w=1.7e-07 $l=6.44981e-07 $layer=licon1_PDIFF $count=1 $X=7.5
+ $Y=2.715 $X2=8.02 $Y2=2.995
r151 3 39 600 $w=1.7e-07 $l=3.92301e-07 $layer=licon1_PDIFF $count=1 $X=5.59
+ $Y=2.715 $X2=5.845 $Y2=3
r152 2 32 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=2.715 $X2=2.59 $Y2=2.925
r153 1 25 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.935
+ $Y=2.66 $X2=1.075 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%A_605_109# 1 2 8 10 16
r32 13 16 4.06667 $w=4.98e-07 $l=1.7e-07 $layer=LI1_cond $X=3.29 $Y=2.925
+ $X2=3.46 $Y2=2.925
r33 10 12 10.7057 $w=3.73e-07 $l=2.35e-07 $layer=LI1_cond $X=3.187 $Y=0.77
+ $X2=3.187 $Y2=1.005
r34 8 13 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=3.29 $Y=2.675 $X2=3.29
+ $Y2=2.925
r35 8 12 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=3.29 $Y=2.675
+ $X2=3.29 $Y2=1.005
r36 2 16 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=2.715 $X2=3.46 $Y2=2.925
r37 1 10 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.545 $X2=3.165 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%Q_N 1 2 7 8 9 10 11 12 13 22
r22 13 40 14.2455 $w=3.58e-07 $l=4.45e-07 $layer=LI1_cond $X=15.195 $Y=3.145
+ $X2=15.195 $Y2=3.59
r23 12 13 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=15.195 $Y=2.775
+ $X2=15.195 $Y2=3.145
r24 11 12 13.9254 $w=3.58e-07 $l=4.35e-07 $layer=LI1_cond $X=15.195 $Y=2.34
+ $X2=15.195 $Y2=2.775
r25 10 11 9.76375 $w=3.58e-07 $l=3.05e-07 $layer=LI1_cond $X=15.195 $Y=2.035
+ $X2=15.195 $Y2=2.34
r26 9 10 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=15.195 $Y=1.665
+ $X2=15.195 $Y2=2.035
r27 8 9 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=15.195 $Y=1.295
+ $X2=15.195 $Y2=1.665
r28 7 8 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=15.195 $Y=0.925
+ $X2=15.195 $Y2=1.295
r29 7 22 8.48326 $w=3.58e-07 $l=2.65e-07 $layer=LI1_cond $X=15.195 $Y=0.925
+ $X2=15.195 $Y2=0.66
r30 2 40 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=15.06
+ $Y=2.215 $X2=15.2 $Y2=3.59
r31 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=15.06
+ $Y=2.215 $X2=15.2 $Y2=2.34
r32 1 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=15.07
+ $Y=0.535 $X2=15.21 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%Q 1 2 7 8 9 10 11 12 13 25 47 50
r16 50 51 2.86126 $w=3.33e-07 $l=5e-08 $layer=LI1_cond $X=17.467 $Y=2.405
+ $X2=17.467 $Y2=2.355
r17 47 48 2.17324 $w=3.33e-07 $l=3e-08 $layer=LI1_cond $X=17.467 $Y=1.295
+ $X2=17.467 $Y2=1.325
r18 37 54 0.0688026 $w=3.33e-07 $l=2e-09 $layer=LI1_cond $X=17.467 $Y=2.522
+ $X2=17.467 $Y2=2.52
r19 13 43 4.30016 $w=3.33e-07 $l=1.25e-07 $layer=LI1_cond $X=17.467 $Y=3.145
+ $X2=17.467 $Y2=3.27
r20 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=17.467 $Y=2.775
+ $X2=17.467 $Y2=3.145
r21 12 37 8.70352 $w=3.33e-07 $l=2.53e-07 $layer=LI1_cond $X=17.467 $Y=2.775
+ $X2=17.467 $Y2=2.522
r22 11 54 3.37133 $w=3.33e-07 $l=9.8e-08 $layer=LI1_cond $X=17.467 $Y=2.422
+ $X2=17.467 $Y2=2.52
r23 11 50 0.584822 $w=3.33e-07 $l=1.7e-08 $layer=LI1_cond $X=17.467 $Y=2.422
+ $X2=17.467 $Y2=2.405
r24 11 51 0.901912 $w=2.28e-07 $l=1.8e-08 $layer=LI1_cond $X=17.52 $Y=2.337
+ $X2=17.52 $Y2=2.355
r25 10 11 15.1321 $w=2.28e-07 $l=3.02e-07 $layer=LI1_cond $X=17.52 $Y=2.035
+ $X2=17.52 $Y2=2.337
r26 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=17.52 $Y=1.665
+ $X2=17.52 $Y2=2.035
r27 8 47 0.963236 $w=3.33e-07 $l=2.8e-08 $layer=LI1_cond $X=17.467 $Y=1.267
+ $X2=17.467 $Y2=1.295
r28 8 23 3.74974 $w=3.33e-07 $l=1.09e-07 $layer=LI1_cond $X=17.467 $Y=1.267
+ $X2=17.467 $Y2=1.158
r29 8 9 15.6832 $w=2.28e-07 $l=3.13e-07 $layer=LI1_cond $X=17.52 $Y=1.352
+ $X2=17.52 $Y2=1.665
r30 8 48 1.35287 $w=2.28e-07 $l=2.7e-08 $layer=LI1_cond $X=17.52 $Y=1.352
+ $X2=17.52 $Y2=1.325
r31 7 23 8.0155 $w=3.33e-07 $l=2.33e-07 $layer=LI1_cond $X=17.467 $Y=0.925
+ $X2=17.467 $Y2=1.158
r32 7 25 9.11634 $w=3.33e-07 $l=2.65e-07 $layer=LI1_cond $X=17.467 $Y=0.925
+ $X2=17.467 $Y2=0.66
r33 2 54 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=17.325
+ $Y=2.395 $X2=17.465 $Y2=2.52
r34 2 43 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=17.325
+ $Y=2.395 $X2=17.465 $Y2=3.27
r35 1 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=17.325
+ $Y=0.535 $X2=17.465 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%VGND 1 2 3 4 5 6 7 22 25 34 47 57 67 71 80
+ 84
r118 86 88 5.90737 $w=9.48e-07 $l=4.6e-07 $layer=LI1_cond $X=16.63 $Y=0.68
+ $X2=16.63 $Y2=1.14
r119 81 84 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=16.27 $Y=0.44
+ $X2=16.99 $Y2=0.44
r120 80 86 2.56842 $w=9.48e-07 $l=2e-07 $layer=LI1_cond $X=16.63 $Y=0.48
+ $X2=16.63 $Y2=0.68
r121 80 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.99 $Y=0.48
+ $X2=16.99 $Y2=0.48
r122 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.27 $Y=0.48
+ $X2=16.27 $Y2=0.48
r123 75 81 0.593134 $w=3.7e-07 $l=1.545e-06 $layer=MET1_cond $X=14.725 $Y=0.44
+ $X2=16.27 $Y2=0.44
r124 72 75 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=14.005 $Y=0.44
+ $X2=14.725 $Y2=0.44
r125 71 77 4.30588 $w=9.33e-07 $l=3.3e-07 $layer=LI1_cond $X=14.367 $Y=0.48
+ $X2=14.367 $Y2=0.81
r126 71 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.725 $Y=0.48
+ $X2=14.725 $Y2=0.48
r127 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.005 $Y=0.48
+ $X2=14.005 $Y2=0.48
r128 68 72 0.372388 $w=3.7e-07 $l=9.7e-07 $layer=MET1_cond $X=13.035 $Y=0.44
+ $X2=14.005 $Y2=0.44
r129 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.035 $Y=0.48
+ $X2=13.035 $Y2=0.48
r130 65 67 0.980392 $w=6.08e-07 $l=5e-08 $layer=LI1_cond $X=12.985 $Y=0.67
+ $X2=13.035 $Y2=0.67
r131 62 68 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=12.315 $Y=0.44
+ $X2=13.035 $Y2=0.44
r132 61 65 13.1373 $w=6.08e-07 $l=6.7e-07 $layer=LI1_cond $X=12.315 $Y=0.67
+ $X2=12.985 $Y2=0.67
r133 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.315 $Y=0.48
+ $X2=12.315 $Y2=0.48
r134 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.62 $Y=0.48
+ $X2=7.62 $Y2=0.48
r135 55 57 0.980392 $w=6.08e-07 $l=5e-08 $layer=LI1_cond $X=7.57 $Y=0.67
+ $X2=7.62 $Y2=0.67
r136 52 58 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=6.9 $Y=0.44
+ $X2=7.62 $Y2=0.44
r137 51 55 13.1373 $w=6.08e-07 $l=6.7e-07 $layer=LI1_cond $X=6.9 $Y=0.67
+ $X2=7.57 $Y2=0.67
r138 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.9 $Y=0.48
+ $X2=6.9 $Y2=0.48
r139 48 52 0.543226 $w=3.7e-07 $l=1.415e-06 $layer=MET1_cond $X=5.485 $Y=0.44
+ $X2=6.9 $Y2=0.44
r140 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.485 $Y=0.48
+ $X2=5.485 $Y2=0.48
r141 45 47 1.10748 $w=5.38e-07 $l=5e-08 $layer=LI1_cond $X=5.435 $Y=0.635
+ $X2=5.485 $Y2=0.635
r142 42 48 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=4.765 $Y=0.44
+ $X2=5.485 $Y2=0.44
r143 41 45 14.8402 $w=5.38e-07 $l=6.7e-07 $layer=LI1_cond $X=4.765 $Y=0.635
+ $X2=5.435 $Y2=0.635
r144 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.765 $Y=0.48
+ $X2=4.765 $Y2=0.48
r145 35 42 0.93289 $w=3.7e-07 $l=2.43e-06 $layer=MET1_cond $X=2.335 $Y=0.44
+ $X2=4.765 $Y2=0.44
r146 34 38 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=2.345 $Y=0.48
+ $X2=2.345 $Y2=0.755
r147 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.335 $Y=0.48
+ $X2=2.335 $Y2=0.48
r148 29 35 0.368549 $w=3.7e-07 $l=9.6e-07 $layer=MET1_cond $X=1.375 $Y=0.44
+ $X2=2.335 $Y2=0.44
r149 26 29 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.655 $Y=0.44
+ $X2=1.375 $Y2=0.44
r150 25 31 3.72421 $w=9.48e-07 $l=2.9e-07 $layer=LI1_cond $X=1.015 $Y=0.48
+ $X2=1.015 $Y2=0.77
r151 25 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.375 $Y=0.48
+ $X2=1.375 $Y2=0.48
r152 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.655 $Y=0.48
+ $X2=0.655 $Y2=0.48
r153 22 62 1.31872 $w=3.7e-07 $l=3.435e-06 $layer=MET1_cond $X=8.88 $Y=0.44
+ $X2=12.315 $Y2=0.44
r154 22 58 0.483721 $w=3.7e-07 $l=1.26e-06 $layer=MET1_cond $X=8.88 $Y=0.44
+ $X2=7.62 $Y2=0.44
r155 7 88 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=16.45
+ $Y=0.865 $X2=16.685 $Y2=1.14
r156 7 86 182 $w=1.7e-07 $l=3.14166e-07 $layer=licon1_NDIFF $count=1 $X=16.45
+ $Y=0.865 $X2=16.685 $Y2=0.68
r157 6 77 182 $w=1.7e-07 $l=2.61056e-07 $layer=licon1_NDIFF $count=1 $X=14.195
+ $Y=0.865 $X2=14.43 $Y2=0.81
r158 5 65 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.845
+ $Y=0.535 $X2=12.985 $Y2=0.745
r159 4 55 182 $w=1.7e-07 $l=3.4821e-07 $layer=licon1_NDIFF $count=1 $X=7.335
+ $Y=0.535 $X2=7.57 $Y2=0.785
r160 3 45 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.545 $X2=5.435 $Y2=0.755
r161 2 38 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.26
+ $Y=0.545 $X2=2.385 $Y2=0.755
r162 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.915
+ $Y=0.56 $X2=1.055 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%A_1642_107# 1 2 9 11 12 15
r34 13 15 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=10.985 $Y=0.545
+ $X2=10.985 $Y2=0.91
r35 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.86 $Y=0.46
+ $X2=10.985 $Y2=0.545
r36 11 12 152.989 $w=1.68e-07 $l=2.345e-06 $layer=LI1_cond $X=10.86 $Y=0.46
+ $X2=8.515 $Y2=0.46
r37 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.35 $Y=0.545
+ $X2=8.515 $Y2=0.46
r38 7 9 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=8.35 $Y=0.545 $X2=8.35
+ $Y2=0.785
r39 2 15 182 $w=1.7e-07 $l=4.41588e-07 $layer=licon1_NDIFF $count=1 $X=10.57
+ $Y=0.765 $X2=10.945 $Y2=0.91
r40 1 9 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=8.21
+ $Y=0.535 $X2=8.35 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSBP_1%A_1755_153# 1 2 7 12 13 14 16 18
r45 18 20 10.5634 $w=3.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.475 $Y=0.745
+ $X2=11.475 $Y2=0.975
r46 16 20 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=11.375 $Y=1.255
+ $X2=11.375 $Y2=0.975
r47 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.29 $Y=1.34
+ $X2=11.375 $Y2=1.255
r48 13 14 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.29 $Y=1.34
+ $X2=10.68 $Y2=1.34
r49 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.595 $Y=1.255
+ $X2=10.68 $Y2=1.34
r50 11 12 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.595 $Y=0.975
+ $X2=10.595 $Y2=1.255
r51 7 11 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.51 $Y=0.85
+ $X2=10.595 $Y2=0.975
r52 7 9 73.2954 $w=2.48e-07 $l=1.59e-06 $layer=LI1_cond $X=10.51 $Y=0.85
+ $X2=8.92 $Y2=0.85
r53 2 18 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=11.37
+ $Y=0.535 $X2=11.495 $Y2=0.745
r54 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=8.775
+ $Y=0.765 $X2=8.92 $Y2=0.89
.ends

