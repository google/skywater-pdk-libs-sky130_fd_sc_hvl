# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  8.140000 ;
  SYMMETRY X Y R90 ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.205000 1.685000 9.895000 2.015000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  7.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.730000 1.830000 5.400000 2.160000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.397500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.755000 1.315000 1.175000 1.605000 ;
        RECT 0.755000 1.605000 0.975000 2.405000 ;
        RECT 0.755000 2.405000 1.175000 2.695000 ;
        RECT 0.955000 0.895000 1.175000 1.315000 ;
        RECT 0.955000 2.695000 1.175000 3.075000 ;
    END
  END X
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 13.850000 3.305000 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 13.920000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 13.920000 8.255000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 13.920000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 13.920000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.985000  0.685000 4.155000 ;
      RECT  0.000000  8.055000 13.920000 8.225000 ;
      RECT  0.360000  4.155000  0.530000 5.280000 ;
      RECT  0.895000  4.575000  2.780000 4.795000 ;
      RECT  0.895000  4.795000  1.115000 6.055000 ;
      RECT  0.895000  6.055000  1.955000 6.275000 ;
      RECT  0.955000  6.445000  1.175000 7.625000 ;
      RECT  0.955000  7.625000  4.900000 7.845000 ;
      RECT  1.365000  5.555000  2.035000 5.665000 ;
      RECT  1.365000  5.665000  5.675000 5.885000 ;
      RECT  1.400000  0.395000  1.990000 0.625000 ;
      RECT  1.735000  6.275000  1.955000 7.455000 ;
      RECT  1.760000  0.625000  1.990000 1.565000 ;
      RECT  1.760000  2.405000  1.930000 3.445000 ;
      RECT  1.760000  3.445000  2.350000 3.735000 ;
      RECT  2.110000  4.295000  2.780000 4.575000 ;
      RECT  2.260000  0.645000  2.480000 2.860000 ;
      RECT  2.260000  2.860000  2.780000 3.085000 ;
      RECT  2.515000  6.445000  2.735000 7.625000 ;
      RECT  2.560000  3.085000  2.780000 4.295000 ;
      RECT  2.650000  1.830000  3.320000 1.940000 ;
      RECT  2.650000  1.940000  4.425000 2.160000 ;
      RECT  3.060000  3.445000  3.645000 3.735000 ;
      RECT  3.175000  0.395000  3.765000 0.625000 ;
      RECT  3.175000  4.410000  3.645000 4.630000 ;
      RECT  3.175000  4.630000  3.395000 5.405000 ;
      RECT  3.295000  5.885000  3.515000 7.455000 ;
      RECT  3.360000  0.625000  3.590000 1.655000 ;
      RECT  3.425000  2.405000  3.645000 3.445000 ;
      RECT  3.425000  3.735000  3.645000 4.410000 ;
      RECT  4.075000  6.445000  4.295000 7.625000 ;
      RECT  4.205000  0.645000  4.425000 1.940000 ;
      RECT  4.205000  2.160000  4.425000 3.755000 ;
      RECT  4.680000  6.295000  8.445000 6.515000 ;
      RECT  4.680000  6.515000  4.900000 7.625000 ;
      RECT  5.455000  4.945000  5.675000 5.665000 ;
      RECT  6.465000  1.305000  6.685000 6.295000 ;
      RECT  7.155000  0.395000  7.745000 0.625000 ;
      RECT  7.340000  0.625000  7.570000 6.055000 ;
      RECT  7.750000  7.075000  9.535000 7.405000 ;
      RECT  8.225000  1.305000  8.445000 6.295000 ;
      RECT  9.100000  3.905000 10.035000 4.235000 ;
      RECT  9.205000  4.775000  9.535000 7.075000 ;
      RECT  9.305000  0.395000  9.895000 0.625000 ;
      RECT  9.305000  3.020000  9.895000 3.365000 ;
      RECT  9.565000  0.625000  9.895000 1.515000 ;
      RECT  9.565000  2.335000  9.895000 3.020000 ;
      RECT  9.565000  3.365000  9.895000 3.905000 ;
      RECT  9.705000  4.235000 10.035000 5.805000 ;
      RECT  9.705000  6.125000 10.535000 6.455000 ;
      RECT  9.705000  6.625000 10.035000 7.520000 ;
      RECT  9.705000  7.520000 10.295000 7.750000 ;
      RECT 10.065000  0.735000 10.395000 3.035000 ;
      RECT 10.065000  3.035000 10.535000 3.365000 ;
      RECT 10.205000  3.365000 10.535000 6.125000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.155000  8.055000  0.325000 8.225000 ;
      RECT  0.515000  3.985000  0.685000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  8.055000  0.805000 8.225000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  8.055000  1.285000 8.225000 ;
      RECT  1.430000  0.425000  1.600000 0.595000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  8.055000  1.765000 8.225000 ;
      RECT  1.790000  0.425000  1.960000 0.595000 ;
      RECT  1.790000  3.505000  1.960000 3.675000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  8.055000  2.245000 8.225000 ;
      RECT  2.150000  3.505000  2.320000 3.675000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  8.055000  2.725000 8.225000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  8.055000  3.205000 8.225000 ;
      RECT  3.090000  3.505000  3.260000 3.675000 ;
      RECT  3.205000  0.425000  3.375000 0.595000 ;
      RECT  3.450000  3.505000  3.620000 3.675000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  8.055000  3.685000 8.225000 ;
      RECT  3.565000  0.425000  3.735000 0.595000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  8.055000  4.165000 8.225000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  8.055000  4.645000 8.225000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  8.055000  5.125000 8.225000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  8.055000  5.605000 8.225000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  8.055000  6.085000 8.225000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  8.055000  6.565000 8.225000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  8.055000  7.045000 8.225000 ;
      RECT  7.185000  0.425000  7.355000 0.595000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  8.055000  7.525000 8.225000 ;
      RECT  7.545000  0.425000  7.715000 0.595000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  8.055000  8.005000 8.225000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  8.055000  8.485000 8.225000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  8.055000  8.965000 8.225000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  8.055000  9.445000 8.225000 ;
      RECT  9.335000  0.425000  9.505000 0.595000 ;
      RECT  9.335000  3.080000  9.505000 3.250000 ;
      RECT  9.695000  0.425000  9.865000 0.595000 ;
      RECT  9.695000  3.080000  9.865000 3.250000 ;
      RECT  9.735000  7.550000  9.905000 7.720000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  8.055000  9.925000 8.225000 ;
      RECT 10.095000  7.550000 10.265000 7.720000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  8.055000 10.405000 8.225000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  8.055000 10.885000 8.225000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  8.055000 11.365000 8.225000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  8.055000 11.845000 8.225000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  8.055000 12.325000 8.225000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  8.055000 12.805000 8.225000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  8.055000 13.285000 8.225000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  8.055000 13.765000 8.225000 ;
    LAYER met1 ;
      RECT 0.000000 -0.115000 13.920000 0.115000 ;
      RECT 0.000000  0.255000 13.920000 0.625000 ;
      RECT 0.000000  3.445000 13.920000 3.815000 ;
  END
END sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1
END LIBRARY
