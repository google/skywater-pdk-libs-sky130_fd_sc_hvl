* File: sky130_fd_sc_hvl__einvn_1.pex.spice
* Created: Wed Sep  2 09:06:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__EINVN_1%VNB 5 7 11 25
r19 7 25 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0.058
r20 7 11 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0
r21 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r22 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVN_1%VPB 4 6 14 21
r23 10 21 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=4.07
+ $X2=1.68 $Y2=4.013
r24 10 14 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=4.07
+ $X2=3.12 $Y2=4.07
r25 9 14 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=3.12 $Y2=4.07
r26 9 10 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r27 6 21 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=4.012
+ $X2=1.68 $Y2=4.013
r28 4 14 52 $w=1.7e-07 $l=3.16221e-06 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=3.12 $Y2=4.07
r29 4 9 52 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVN_1%TE_B 3 7 9 11 13 14 15 16 26 27
c45 16 0 4.80347e-20 $X=1.68 $Y=2.035
r46 25 27 3.51593 $w=2.93e-07 $l=9e-08 $layer=LI1_cond $X=1.02 $Y=1.972 $X2=0.93
+ $Y2=1.972
r47 24 26 43.5109 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.02 $Y=1.855
+ $X2=1.185 $Y2=1.855
r48 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.02
+ $Y=1.91 $X2=1.02 $Y2=1.91
r49 22 24 27.8215 $w=5e-07 $l=2.6e-07 $layer=POLY_cond $X=0.76 $Y=1.855 $X2=1.02
+ $Y2=1.855
r50 20 22 10.1656 $w=5e-07 $l=9.5e-08 $layer=POLY_cond $X=0.665 $Y=1.855
+ $X2=0.76 $Y2=1.855
r51 15 16 18.7516 $w=2.93e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.972
+ $X2=1.68 $Y2=1.972
r52 15 25 7.03186 $w=2.93e-07 $l=1.8e-07 $layer=LI1_cond $X=1.2 $Y=1.972
+ $X2=1.02 $Y2=1.972
r53 14 27 8.81998 $w=2.95e-07 $l=2.1e-07 $layer=LI1_cond $X=0.72 $Y=1.972
+ $X2=0.93 $Y2=1.972
r54 11 13 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.815 $Y=2.105
+ $X2=1.815 $Y2=2.965
r55 9 11 36.9698 $w=1.65e-07 $l=2.88531e-07 $layer=POLY_cond $X=1.565 $Y=2.022
+ $X2=1.815 $Y2=2.105
r56 9 26 165.535 $w=1.65e-07 $l=3.8e-07 $layer=POLY_cond $X=1.565 $Y=2.022
+ $X2=1.185 $Y2=2.022
r57 5 22 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.76 $Y=2.105 $X2=0.76
+ $Y2=1.855
r58 5 7 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.76 $Y=2.105 $X2=0.76
+ $Y2=2.61
r59 1 20 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.665 $Y=1.605
+ $X2=0.665 $Y2=1.855
r60 1 3 56.7131 $w=5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.665 $Y=1.605 $X2=0.665
+ $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVN_1%A_30_173# 1 2 7 9 12 15 20 21 23 25
c42 21 0 3.79452e-20 $X=1.9 $Y=1.56
r43 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.9 $Y=1.56
+ $X2=1.9 $Y2=1.56
r44 18 23 2.51069 $w=2.2e-07 $l=1.75e-07 $layer=LI1_cond $X=0.44 $Y=1.535
+ $X2=0.265 $Y2=1.535
r45 18 20 76.4803 $w=2.18e-07 $l=1.46e-06 $layer=LI1_cond $X=0.44 $Y=1.535
+ $X2=1.9 $Y2=1.535
r46 15 25 6.65996 $w=4.19e-07 $l=2.07123e-07 $layer=LI1_cond $X=0.217 $Y=2.195
+ $X2=0.312 $Y2=2.36
r47 14 23 3.93362 $w=3.02e-07 $l=1.31833e-07 $layer=LI1_cond $X=0.217 $Y=1.645
+ $X2=0.265 $Y2=1.535
r48 14 15 24.8566 $w=2.53e-07 $l=5.5e-07 $layer=LI1_cond $X=0.217 $Y=1.645
+ $X2=0.217 $Y2=2.195
r49 10 23 3.93362 $w=3.02e-07 $l=1.1e-07 $layer=LI1_cond $X=0.265 $Y=1.425
+ $X2=0.265 $Y2=1.535
r50 10 12 11.5244 $w=3.48e-07 $l=3.5e-07 $layer=LI1_cond $X=0.265 $Y=1.425
+ $X2=0.265 $Y2=1.075
r51 7 21 5.58609 $w=3.02e-07 $l=3.5e-08 $layer=POLY_cond $X=1.935 $Y=1.562
+ $X2=1.9 $Y2=1.562
r52 7 9 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.935 $Y=1.395 $X2=1.935
+ $Y2=0.91
r53 2 25 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.225
+ $Y=2.235 $X2=0.37 $Y2=2.36
r54 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.865 $X2=0.275 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVN_1%A 3 5 6 7 8 17 23 34 37
c36 6 0 3.79452e-20 $X=2.555 $Y=1.58
c37 3 0 4.80347e-20 $X=2.645 $Y=2.965
r38 35 37 1.37371 $w=5.03e-07 $l=5.8e-08 $layer=LI1_cond $X=2.527 $Y=1.977
+ $X2=2.527 $Y2=2.035
r39 34 43 2.51442 $w=2.73e-07 $l=6e-08 $layer=LI1_cond $X=2.642 $Y=1.665
+ $X2=2.642 $Y2=1.725
r40 23 26 16.3989 $w=6.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=1.89
+ $X2=2.585 $Y2=2.055
r41 23 25 16.3989 $w=6.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=1.89
+ $X2=2.585 $Y2=1.725
r42 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.44
+ $Y=1.89 $X2=2.44 $Y2=1.89
r43 20 25 17.656 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.56
+ $X2=2.645 $Y2=1.725
r44 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.695
+ $Y=1.56 $X2=2.695 $Y2=1.56
r45 17 20 69.5538 $w=5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.645 $Y=0.91
+ $X2=2.645 $Y2=1.56
r46 7 35 0.331586 $w=5.03e-07 $l=1.4e-08 $layer=LI1_cond $X=2.527 $Y=1.963
+ $X2=2.527 $Y2=1.977
r47 7 24 1.72898 $w=5.03e-07 $l=7.3e-08 $layer=LI1_cond $X=2.527 $Y=1.963
+ $X2=2.527 $Y2=1.89
r48 7 8 8.45545 $w=5.03e-07 $l=3.57e-07 $layer=LI1_cond $X=2.527 $Y=2.048
+ $X2=2.527 $Y2=2.405
r49 7 37 0.307901 $w=5.03e-07 $l=1.3e-08 $layer=LI1_cond $X=2.527 $Y=2.048
+ $X2=2.527 $Y2=2.035
r50 6 24 3.62376 $w=5.03e-07 $l=1.53e-07 $layer=LI1_cond $X=2.527 $Y=1.737
+ $X2=2.527 $Y2=1.89
r51 6 43 2.74792 $w=5.03e-07 $l=1.2e-08 $layer=LI1_cond $X=2.527 $Y=1.737
+ $X2=2.527 $Y2=1.725
r52 6 34 0.544791 $w=2.73e-07 $l=1.3e-08 $layer=LI1_cond $X=2.642 $Y=1.652
+ $X2=2.642 $Y2=1.665
r53 6 21 3.85545 $w=2.73e-07 $l=9.2e-08 $layer=LI1_cond $X=2.642 $Y=1.652
+ $X2=2.642 $Y2=1.56
r54 5 21 11.1054 $w=2.73e-07 $l=2.65e-07 $layer=LI1_cond $X=2.642 $Y=1.295
+ $X2=2.642 $Y2=1.56
r55 3 26 97.3754 $w=5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.645 $Y=2.965
+ $X2=2.645 $Y2=2.055
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVN_1%VPWR 1 4 11 14
r25 11 14 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.655 $Y=3.59
+ $X2=2.655 $Y2=3.59
r26 11 12 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.855 $Y=3.59
+ $X2=0.855 $Y2=3.59
r27 9 11 2.64929 $w=1.842e-06 $l=4e-07 $layer=LI1_cond $X=1.755 $Y=3.19
+ $X2=1.755 $Y2=3.59
r28 7 9 5.3317 $w=1.842e-06 $l=8.05e-07 $layer=LI1_cond $X=1.755 $Y=2.385
+ $X2=1.755 $Y2=3.19
r29 4 14 0.374308 $w=3.7e-07 $l=9.75e-07 $layer=MET1_cond $X=1.68 $Y=3.63
+ $X2=2.655 $Y2=3.63
r30 4 12 0.316722 $w=3.7e-07 $l=8.25e-07 $layer=MET1_cond $X=1.68 $Y=3.63
+ $X2=0.855 $Y2=3.63
r31 1 9 300 $w=1.7e-07 $l=1.12276e-06 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=2.235 $X2=1.375 $Y2=3.19
r32 1 7 300 $w=1.7e-07 $l=4.33561e-07 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=2.235 $X2=1.375 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVN_1%Z 1 2 7 8 9 10 11 12 13 22
r13 13 40 17.9943 $w=2.83e-07 $l=4.45e-07 $layer=LI1_cond $X=3.092 $Y=3.145
+ $X2=3.092 $Y2=3.59
r14 12 13 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.092 $Y=2.775
+ $X2=3.092 $Y2=3.145
r15 11 12 17.5899 $w=2.83e-07 $l=4.35e-07 $layer=LI1_cond $X=3.092 $Y=2.34
+ $X2=3.092 $Y2=2.775
r16 10 11 12.3332 $w=2.83e-07 $l=3.05e-07 $layer=LI1_cond $X=3.092 $Y=2.035
+ $X2=3.092 $Y2=2.34
r17 9 10 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.092 $Y=1.665
+ $X2=3.092 $Y2=2.035
r18 8 9 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.092 $Y=1.295
+ $X2=3.092 $Y2=1.665
r19 7 8 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.092 $Y=0.925
+ $X2=3.092 $Y2=1.295
r20 7 22 10.7157 $w=2.83e-07 $l=2.65e-07 $layer=LI1_cond $X=3.092 $Y=0.925
+ $X2=3.092 $Y2=0.66
r21 2 40 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.895
+ $Y=2.215 $X2=3.035 $Y2=3.59
r22 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.895
+ $Y=2.215 $X2=3.035 $Y2=2.34
r23 1 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.895
+ $Y=0.535 $X2=3.035 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVN_1%VGND 1 4 10 12
r22 12 14 2.95973 $w=2.061e-06 $l=5e-07 $layer=LI1_cond $X=1.605 $Y=0.66
+ $X2=1.605 $Y2=1.16
r23 7 12 1.0655 $w=2.061e-06 $l=1.8e-07 $layer=LI1_cond $X=1.605 $Y=0.48
+ $X2=1.605 $Y2=0.66
r24 7 10 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.685 $Y=0.48
+ $X2=2.685 $Y2=0.48
r25 7 8 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.525 $Y=0.48
+ $X2=0.525 $Y2=0.48
r26 4 10 0.385825 $w=3.7e-07 $l=1.005e-06 $layer=MET1_cond $X=1.68 $Y=0.44
+ $X2=2.685 $Y2=0.44
r27 4 8 0.443411 $w=3.7e-07 $l=1.155e-06 $layer=MET1_cond $X=1.68 $Y=0.44
+ $X2=0.525 $Y2=0.44
r28 1 14 91 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=2 $X=0.915
+ $Y=0.865 $X2=1.055 $Y2=1.16
r29 1 12 91 $w=1.7e-07 $l=7.25293e-07 $layer=licon1_NDIFF $count=2 $X=0.915
+ $Y=0.865 $X2=1.545 $Y2=0.66
.ends

