* NGSPICE file created from sky130_fd_sc_hvl__lsbufhv2lv_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VNB VPB VPWR X
M1000 a_30_1337# A VPWR VPB phv w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=1.197e+11p ps=1.41e+06u
M1001 LVPWR a_389_1337# a_389_141# LVPWR phighvt w=1.12e+06u l=150000u
+  ad=6.104e+11p pd=5.57e+06u as=2.968e+11p ps=2.77e+06u
M1002 a_187_207# a_30_1337# a_30_207# VNB nhv w=420000u l=500000u
+  ad=9.54e+11p pd=8.61e+06u as=1.197e+11p ps=1.41e+06u
M1003 LVPWR a_389_141# X LVPWR phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=2.968e+11p ps=2.77e+06u
M1004 a_187_207# a_30_207# a_389_141# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=6.075e+11p ps=6.12e+06u
M1005 a_389_1337# a_30_1337# VGND VNB nhv w=750000u l=500000u
+  ad=6.075e+11p pd=6.12e+06u as=7.665e+11p ps=6.61e+06u
M1006 a_187_207# a_30_207# a_389_141# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_187_207# a_30_207# a_389_141# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_30_1337# a_389_1337# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_30_1337# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1010 a_389_141# a_30_207# a_187_207# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_187_207# a_389_141# X VNB nshort w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=1.961e+11p ps=2.01e+06u
M1012 VGND a_30_1337# a_389_1337# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_389_1337# a_389_141# LVPWR LVPWR phighvt w=1.12e+06u l=150000u
+  ad=2.968e+11p pd=2.77e+06u as=0p ps=0u
M1014 a_389_1337# a_30_1337# VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_30_207# a_30_1337# a_30_443# VPB phv w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=1.197e+11p ps=1.41e+06u
.ends

