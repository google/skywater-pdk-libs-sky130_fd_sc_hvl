* File: sky130_fd_sc_hvl__a21oi_1.spice
* Created: Wed Sep  2 09:03:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__a21oi_1.pex.spice"
.subckt sky130_fd_sc_hvl__a21oi_1  VNB VPB A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1000 A_271_107# N_A2_M1000_g N_VGND_M1000_s N_VNB_M1000_b NHV L=0.5 W=0.75
+ AD=0.07875 AS=0.21375 PD=0.96 PS=2.07 NRD=7.5924 NRS=0 M=1 R=1.5 SA=250000
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1004 N_Y_M1004_d N_A1_M1004_g A_271_107# N_VNB_M1000_b NHV L=0.5 W=0.75
+ AD=0.1425 AS=0.07875 PD=1.13 PS=0.96 NRD=15.1962 NRS=7.5924 M=1 R=1.5
+ SA=250001 SB=250001 A=0.375 P=2.5 MULT=1
MM1002 N_VGND_M1002_d N_B1_M1002_g N_Y_M1004_d N_VNB_M1000_b NHV L=0.5 W=0.75
+ AD=0.19875 AS=0.1425 PD=2.03 PS=1.13 NRD=0 NRS=0 M=1 R=1.5 SA=250002 SB=250000
+ A=0.375 P=2.5 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_56_443#_M1003_s N_VPB_M1003_b PHV L=0.5
+ W=1.5 AD=0.375 AS=0.4275 PD=2 PS=3.57 NRD=0 NRS=0 M=1 R=3 SA=250000 SB=250002
+ A=0.75 P=4 MULT=1
MM1005 N_A_56_443#_M1005_d N_A1_M1005_g N_VPWR_M1003_d N_VPB_M1003_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.375 PD=1.78 PS=2 NRD=0 NRS=28.0006 M=1 R=3 SA=250001
+ SB=250001 A=0.75 P=4 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_A_56_443#_M1005_d N_VPB_M1003_b PHV L=0.5
+ W=1.5 AD=0.5475 AS=0.21 PD=3.73 PS=1.78 NRD=10.1803 NRS=0 M=1 R=3 SA=250002
+ SB=250000 A=0.75 P=4 MULT=1
DX6_noxref N_VNB_M1000_b N_VPB_M1003_b NWDIODE A=10.452 P=13.24
*
.include "sky130_fd_sc_hvl__a21oi_1.pxi.spice"
*
.ends
*
*
