* File: sky130_fd_sc_hvl__probe_p_8.pxi.spice
* Created: Fri Aug 28 09:39:22 2020
* 
x_PM_SKY130_FD_SC_HVL__PROBE_P_8%VNB N_VNB_M1003_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__PROBE_P_8%VNB
x_PM_SKY130_FD_SC_HVL__PROBE_P_8%VPB N_VPB_M1006_b VPB N_VPB_c_44_p VPB
+ PM_SKY130_FD_SC_HVL__PROBE_P_8%VPB
x_PM_SKY130_FD_SC_HVL__PROBE_P_8%A N_A_M1006_g N_A_c_124_n N_A_M1003_g
+ N_A_c_126_n N_A_c_127_n N_A_M1008_g N_A_M1007_g N_A_c_128_n N_A_M1015_g
+ N_A_M1019_g N_A_c_129_n A A A A N_A_c_130_n PM_SKY130_FD_SC_HVL__PROBE_P_8%A
x_PM_SKY130_FD_SC_HVL__PROBE_P_8%A_45_443# N_A_45_443#_M1003_d
+ N_A_45_443#_M1008_d N_A_45_443#_M1006_s N_A_45_443#_M1007_s
+ N_A_45_443#_M1001_g N_A_45_443#_c_210_n N_A_45_443#_M1000_g
+ N_A_45_443#_M1002_g N_A_45_443#_c_213_n N_A_45_443#_M1004_g
+ N_A_45_443#_M1009_g N_A_45_443#_c_216_n N_A_45_443#_M1005_g
+ N_A_45_443#_M1013_g N_A_45_443#_c_219_n N_A_45_443#_M1010_g
+ N_A_45_443#_M1014_g N_A_45_443#_c_222_n N_A_45_443#_M1011_g
+ N_A_45_443#_M1018_g N_A_45_443#_c_225_n N_A_45_443#_M1012_g
+ N_A_45_443#_M1020_g N_A_45_443#_c_228_n N_A_45_443#_M1016_g
+ N_A_45_443#_M1021_g N_A_45_443#_c_231_n N_A_45_443#_M1017_g
+ N_A_45_443#_c_244_n N_A_45_443#_c_206_n N_A_45_443#_c_235_n
+ N_A_45_443#_c_237_n N_A_45_443#_c_252_n N_A_45_443#_c_416_p
+ N_A_45_443#_c_254_n N_A_45_443#_c_258_n N_A_45_443#_c_207_n
+ N_A_45_443#_c_208_n N_A_45_443#_c_239_n N_A_45_443#_c_240_n
+ N_A_45_443#_c_265_n N_A_45_443#_c_268_n N_A_45_443#_c_209_n
+ PM_SKY130_FD_SC_HVL__PROBE_P_8%A_45_443#
x_PM_SKY130_FD_SC_HVL__PROBE_P_8%VPWR N_VPWR_M1006_d N_VPWR_M1019_d
+ N_VPWR_M1004_s N_VPWR_M1010_s N_VPWR_M1012_s N_VPWR_M1017_s N_VPWR_c_464_n
+ N_VPWR_c_467_n N_VPWR_c_470_n N_VPWR_c_473_n N_VPWR_c_476_n N_VPWR_c_477_n
+ N_VPWR_c_478_n N_VPWR_c_481_n N_VPWR_c_484_n N_VPWR_c_487_n VPWR
+ N_VPWR_c_502_n N_VPWR_c_532_n N_VPWR_c_537_n N_VPWR_c_542_n N_VPWR_c_490_n
+ N_VPWR_c_493_n N_VPWR_c_496_n PM_SKY130_FD_SC_HVL__PROBE_P_8%VPWR
x_PM_SKY130_FD_SC_HVL__PROBE_P_8%noxref_6 N_noxref_6_M1001_d N_noxref_6_M1009_d
+ N_noxref_6_M1014_d N_noxref_6_M1020_d N_noxref_6_M1000_d N_noxref_6_M1005_d
+ N_noxref_6_M1011_d N_noxref_6_M1016_d N_noxref_6_c_615_n N_noxref_6_c_604_n
+ N_noxref_6_c_620_n N_noxref_6_c_621_n N_noxref_6_c_609_n N_noxref_6_c_626_n
+ N_noxref_6_c_629_n N_noxref_6_c_605_n N_noxref_6_c_634_n N_noxref_6_c_610_n
+ N_noxref_6_c_638_n N_noxref_6_c_606_n N_noxref_6_c_643_n N_noxref_6_c_644_n
+ N_noxref_6_c_646_n N_noxref_6_c_760_p N_noxref_6_c_607_n N_noxref_6_c_651_n
+ N_noxref_6_c_652_n N_noxref_6_c_654_n N_noxref_6_c_657_n N_noxref_6_c_658_n
+ N_noxref_6_c_661_n N_noxref_6_c_611_n N_noxref_6_c_665_n N_noxref_6_c_668_n
+ N_noxref_6_c_671_n N_noxref_6_c_673_n N_noxref_6_c_608_n N_noxref_6_c_613_n
+ N_noxref_6_c_704_n N_noxref_6_R23_noxref_pos N_noxref_6_c_705_n
+ PM_SKY130_FD_SC_HVL__PROBE_P_8%noxref_6
x_PM_SKY130_FD_SC_HVL__PROBE_P_8%VGND N_VGND_M1003_s N_VGND_M1015_s
+ N_VGND_M1002_s N_VGND_M1013_s N_VGND_M1018_s N_VGND_M1021_s N_VGND_c_772_n
+ N_VGND_c_773_n VGND N_VGND_c_774_n N_VGND_c_776_n N_VGND_c_778_n
+ N_VGND_c_780_n N_VGND_c_781_n N_VGND_c_782_n N_VGND_c_783_n N_VGND_c_784_n
+ N_VGND_c_785_n N_VGND_c_786_n N_VGND_c_787_n
+ PM_SKY130_FD_SC_HVL__PROBE_P_8%VGND
x_PM_SKY130_FD_SC_HVL__PROBE_P_8%X X N_X_R23_noxref_neg
+ PM_SKY130_FD_SC_HVL__PROBE_P_8%X
cc_1 N_VNB_M1003_b N_A_c_124_n 0.0456634f $X=-0.33 $Y=-0.265 $X2=0.78 $Y2=1.565
cc_2 N_VNB_c_2_p N_A_c_124_n 5.58874e-19 $X=0.24 $Y=0 $X2=0.78 $Y2=1.565
cc_3 N_VNB_M1003_b N_A_c_126_n 0.0274014f $X=-0.33 $Y=-0.265 $X2=1.57 $Y2=1.815
cc_4 N_VNB_M1003_b N_A_c_127_n 0.0391903f $X=-0.33 $Y=-0.265 $X2=1.82 $Y2=1.565
cc_5 N_VNB_M1003_b N_A_c_128_n 0.0378062f $X=-0.33 $Y=-0.265 $X2=2.6 $Y2=1.565
cc_6 N_VNB_M1003_b N_A_c_129_n 0.0267973f $X=-0.33 $Y=-0.265 $X2=0.77 $Y2=1.815
cc_7 N_VNB_M1003_b N_A_c_130_n 0.0506531f $X=-0.33 $Y=-0.265 $X2=2.6 $Y2=1.815
cc_8 N_VNB_M1003_b N_A_45_443#_M1001_g 0.0406558f $X=-0.33 $Y=-0.265 $X2=1.82
+ $Y2=2.965
cc_9 N_VNB_M1003_b N_A_45_443#_M1002_g 0.0399246f $X=-0.33 $Y=-0.265 $X2=2.6
+ $Y2=2.965
cc_10 N_VNB_M1003_b N_A_45_443#_M1009_g 0.0399246f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1003_b N_A_45_443#_M1013_g 0.0399246f $X=-0.33 $Y=-0.265 $X2=1.82
+ $Y2=1.815
cc_12 N_VNB_M1003_b N_A_45_443#_M1014_g 0.0403249f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1003_b N_A_45_443#_M1018_g 0.0406374f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_M1003_b N_A_45_443#_M1020_g 0.0400078f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_15 N_VNB_M1003_b N_A_45_443#_M1021_g 0.0475743f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_16 N_VNB_M1003_b N_A_45_443#_c_206_n 0.0201484f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_17 N_VNB_M1003_b N_A_45_443#_c_207_n 0.00264768f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1003_b N_A_45_443#_c_208_n 0.00132121f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_19 N_VNB_M1003_b N_A_45_443#_c_209_n 0.219325f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_20 N_VNB_M1003_b N_noxref_6_c_604_n 0.00805267f $X=-0.33 $Y=-0.265 $X2=1.735
+ $Y2=1.815
cc_21 N_VNB_M1003_b N_noxref_6_c_605_n 0.00805267f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_22 N_VNB_M1003_b N_noxref_6_c_606_n 0.00270308f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_23 N_VNB_M1003_b N_noxref_6_c_607_n 0.00201572f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_24 N_VNB_M1003_b N_noxref_6_c_608_n 0.00160124f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_25 N_VNB_M1003_b N_VGND_c_772_n 0.0113819f $X=-0.33 $Y=-0.265 $X2=2.6
+ $Y2=1.08
cc_26 N_VNB_M1003_b N_VGND_c_773_n 0.0421164f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_27 N_VNB_M1003_b N_VGND_c_774_n 0.090476f $X=-0.33 $Y=-0.265 $X2=1.68
+ $Y2=1.697
cc_28 N_VNB_c_2_p N_VGND_c_774_n 0.00538291f $X=0.24 $Y=0 $X2=1.68 $Y2=1.697
cc_29 N_VNB_M1003_b N_VGND_c_776_n 0.0421797f $X=-0.33 $Y=-0.265 $X2=2.16
+ $Y2=1.697
cc_30 N_VNB_c_2_p N_VGND_c_776_n 0.00247336f $X=0.24 $Y=0 $X2=2.16 $Y2=1.697
cc_31 N_VNB_M1003_b N_VGND_c_778_n 0.251101f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_32 N_VNB_c_2_p N_VGND_c_778_n 0.0168113f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_33 N_VNB_M1003_b N_VGND_c_780_n 0.00648157f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_34 N_VNB_M1003_b N_VGND_c_781_n 0.00846255f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_35 N_VNB_M1003_b N_VGND_c_782_n 0.00648157f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_36 N_VNB_M1003_b N_VGND_c_783_n 0.00846255f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_37 N_VNB_M1003_b N_VGND_c_784_n 0.00659769f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_38 N_VNB_M1003_b N_VGND_c_785_n 0.0125522f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_39 N_VNB_M1003_b N_VGND_c_786_n 0.00867563f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_40 N_VNB_M1003_b N_VGND_c_787_n 0.151233f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_41 N_VNB_c_2_p N_VGND_c_787_n 1.02625f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_42 N_VPB_M1006_b N_A_M1006_g 0.0429652f $X=-0.33 $Y=1.885 $X2=0.76 $Y2=2.965
cc_43 VPB N_A_M1006_g 0.00970178f $X=0 $Y=3.955 $X2=0.76 $Y2=2.965
cc_44 N_VPB_c_44_p N_A_M1006_g 0.0148199f $X=9.36 $Y=4.07 $X2=0.76 $Y2=2.965
cc_45 N_VPB_M1006_b N_A_c_126_n 0.0193995f $X=-0.33 $Y=1.885 $X2=1.57 $Y2=1.815
cc_46 N_VPB_M1006_b N_A_M1007_g 0.0378158f $X=-0.33 $Y=1.885 $X2=1.82 $Y2=2.965
cc_47 VPB N_A_M1007_g 0.00970178f $X=0 $Y=3.955 $X2=1.82 $Y2=2.965
cc_48 N_VPB_c_44_p N_A_M1007_g 0.013528f $X=9.36 $Y=4.07 $X2=1.82 $Y2=2.965
cc_49 N_VPB_M1006_b N_A_M1019_g 0.0364141f $X=-0.33 $Y=1.885 $X2=2.6 $Y2=2.965
cc_50 VPB N_A_M1019_g 0.00970178f $X=0 $Y=3.955 $X2=2.6 $Y2=2.965
cc_51 N_VPB_c_44_p N_A_M1019_g 0.0135178f $X=9.36 $Y=4.07 $X2=2.6 $Y2=2.965
cc_52 N_VPB_M1006_b N_A_c_129_n 0.0144517f $X=-0.33 $Y=1.885 $X2=0.77 $Y2=1.815
cc_53 N_VPB_M1006_b N_A_c_130_n 0.0299911f $X=-0.33 $Y=1.885 $X2=2.6 $Y2=1.815
cc_54 N_VPB_M1006_b N_A_45_443#_c_210_n 0.0328513f $X=-0.33 $Y=1.885 $X2=2.6
+ $Y2=1.565
cc_55 VPB N_A_45_443#_c_210_n 0.00970178f $X=0 $Y=3.955 $X2=2.6 $Y2=1.565
cc_56 N_VPB_c_44_p N_A_45_443#_c_210_n 0.0135156f $X=9.36 $Y=4.07 $X2=2.6
+ $Y2=1.565
cc_57 N_VPB_M1006_b N_A_45_443#_c_213_n 0.0320774f $X=-0.33 $Y=1.885 $X2=0.77
+ $Y2=1.815
cc_58 VPB N_A_45_443#_c_213_n 0.00970178f $X=0 $Y=3.955 $X2=0.77 $Y2=1.815
cc_59 N_VPB_c_44_p N_A_45_443#_c_213_n 0.0135156f $X=9.36 $Y=4.07 $X2=0.77
+ $Y2=1.815
cc_60 N_VPB_M1006_b N_A_45_443#_c_216_n 0.0320774f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_61 VPB N_A_45_443#_c_216_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_62 N_VPB_c_44_p N_A_45_443#_c_216_n 0.0135156f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_63 N_VPB_M1006_b N_A_45_443#_c_219_n 0.032061f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_64 VPB N_A_45_443#_c_219_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_65 N_VPB_c_44_p N_A_45_443#_c_219_n 0.0135156f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_66 N_VPB_M1006_b N_A_45_443#_c_222_n 0.032061f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_67 VPB N_A_45_443#_c_222_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_68 N_VPB_c_44_p N_A_45_443#_c_222_n 0.0135156f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_69 N_VPB_M1006_b N_A_45_443#_c_225_n 0.0321055f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_70 VPB N_A_45_443#_c_225_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_71 N_VPB_c_44_p N_A_45_443#_c_225_n 0.0135156f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_72 N_VPB_M1006_b N_A_45_443#_c_228_n 0.0321054f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_73 VPB N_A_45_443#_c_228_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_74 N_VPB_c_44_p N_A_45_443#_c_228_n 0.0135156f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_75 N_VPB_M1006_b N_A_45_443#_c_231_n 0.0390747f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_76 VPB N_A_45_443#_c_231_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_77 N_VPB_c_44_p N_A_45_443#_c_231_n 0.0135186f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_78 N_VPB_M1006_b N_A_45_443#_c_206_n 0.00998322f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_79 VPB N_A_45_443#_c_235_n 4.22267e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_80 N_VPB_c_44_p N_A_45_443#_c_235_n 0.00452125f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_81 N_VPB_M1006_b N_A_45_443#_c_237_n 0.00764217f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_82 N_VPB_M1006_b N_A_45_443#_c_207_n 0.00381808f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_83 N_VPB_M1006_b N_A_45_443#_c_239_n 0.00526456f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_84 N_VPB_M1006_b N_A_45_443#_c_240_n 0.00544073f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_85 N_VPB_M1006_b N_A_45_443#_c_209_n 0.17523f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_86 N_VPB_M1006_b N_VPWR_c_464_n 0.0010569f $X=-0.33 $Y=1.885 $X2=2.6 $Y2=1.08
cc_87 VPB N_VPWR_c_464_n 0.00362936f $X=0 $Y=3.955 $X2=2.6 $Y2=1.08
cc_88 N_VPB_c_44_p N_VPWR_c_464_n 0.054215f $X=9.36 $Y=4.07 $X2=2.6 $Y2=1.08
cc_89 N_VPB_M1006_b N_VPWR_c_467_n 0.0010569f $X=-0.33 $Y=1.885 $X2=2.6
+ $Y2=2.965
cc_90 VPB N_VPWR_c_467_n 0.00262607f $X=0 $Y=3.955 $X2=2.6 $Y2=2.965
cc_91 N_VPB_c_44_p N_VPWR_c_467_n 0.0405322f $X=9.36 $Y=4.07 $X2=2.6 $Y2=2.965
cc_92 N_VPB_M1006_b N_VPWR_c_470_n 0.0010569f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_470_n 0.00262607f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_94 N_VPB_c_44_p N_VPWR_c_470_n 0.0405322f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_95 N_VPB_M1006_b N_VPWR_c_473_n 0.0010569f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_96 VPB N_VPWR_c_473_n 0.00262607f $X=0 $Y=3.955 $X2=0.635 $Y2=1.58
cc_97 N_VPB_c_44_p N_VPWR_c_473_n 0.0405322f $X=9.36 $Y=4.07 $X2=0.635 $Y2=1.58
cc_98 N_VPB_M1006_b N_VPWR_c_476_n 0.00769488f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_99 N_VPB_M1006_b N_VPWR_c_477_n 0.0525239f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_100 N_VPB_M1006_b N_VPWR_c_478_n 0.00105831f $X=-0.33 $Y=1.885 $X2=1.82
+ $Y2=1.815
cc_101 VPB N_VPWR_c_478_n 0.00279423f $X=0 $Y=3.955 $X2=1.82 $Y2=1.815
cc_102 N_VPB_c_44_p N_VPWR_c_478_n 0.0413412f $X=9.36 $Y=4.07 $X2=1.82 $Y2=1.815
cc_103 N_VPB_M1006_b N_VPWR_c_481_n 0.00105831f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_481_n 0.00385318f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_105 N_VPB_c_44_p N_VPWR_c_481_n 0.0545489f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_106 N_VPB_M1006_b N_VPWR_c_484_n 0.00105831f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_484_n 0.00385318f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_108 N_VPB_c_44_p N_VPWR_c_484_n 0.0545489f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_109 N_VPB_M1006_b N_VPWR_c_487_n 0.00105831f $X=-0.33 $Y=1.885 $X2=1.2
+ $Y2=1.697
cc_110 VPB N_VPWR_c_487_n 0.00385318f $X=0 $Y=3.955 $X2=1.2 $Y2=1.697
cc_111 N_VPB_c_44_p N_VPWR_c_487_n 0.0545489f $X=9.36 $Y=4.07 $X2=1.2 $Y2=1.697
cc_112 N_VPB_M1006_b N_VPWR_c_490_n 0.00270841f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_490_n 0.00513943f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_114 N_VPB_c_44_p N_VPWR_c_490_n 0.0771568f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_115 N_VPB_M1006_b N_VPWR_c_493_n 0.0010569f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_493_n 0.00535847f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_117 N_VPB_c_44_p N_VPWR_c_493_n 0.0847751f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_118 N_VPB_M1006_b N_VPWR_c_496_n 0.0587432f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_496_n 1.01609f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_120 N_VPB_c_44_p N_VPWR_c_496_n 0.033555f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_121 N_VPB_M1006_b N_noxref_6_c_609_n 0.00173812f $X=-0.33 $Y=1.885 $X2=2.6
+ $Y2=1.815
cc_122 N_VPB_M1006_b N_noxref_6_c_610_n 9.9481e-19 $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_123 N_VPB_M1006_b N_noxref_6_c_611_n 0.00261732f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_124 N_A_c_128_n N_A_45_443#_M1001_g 0.0206085f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_125 N_A_M1019_g N_A_45_443#_c_210_n 0.0206085f $X=2.6 $Y=2.965 $X2=9.36 $Y2=0
cc_126 N_A_c_124_n N_A_45_443#_c_244_n 0.00436519f $X=0.78 $Y=1.565 $X2=0 $Y2=0
cc_127 N_A_c_124_n N_A_45_443#_c_206_n 0.00386514f $X=0.78 $Y=1.565 $X2=0 $Y2=0
cc_128 N_A_c_129_n N_A_45_443#_c_206_n 0.0206904f $X=0.77 $Y=1.815 $X2=0 $Y2=0
cc_129 A N_A_45_443#_c_206_n 0.0165919f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_130 N_A_M1006_g N_A_45_443#_c_237_n 0.0358157f $X=0.76 $Y=2.965 $X2=0 $Y2=0
cc_131 N_A_c_126_n N_A_45_443#_c_237_n 0.011632f $X=1.57 $Y=1.815 $X2=0 $Y2=0
cc_132 N_A_M1007_g N_A_45_443#_c_237_n 0.0313016f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_133 A N_A_45_443#_c_237_n 0.0678558f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_134 N_A_M1007_g N_A_45_443#_c_252_n 0.0260651f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_135 N_A_M1019_g N_A_45_443#_c_252_n 0.0458362f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_136 N_A_c_127_n N_A_45_443#_c_254_n 9.17632e-19 $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_137 N_A_c_128_n N_A_45_443#_c_254_n 0.00801446f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_138 A N_A_45_443#_c_254_n 0.00316816f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A_c_130_n N_A_45_443#_c_254_n 0.00323912f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_140 N_A_M1019_g N_A_45_443#_c_258_n 0.00130677f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_141 N_A_c_130_n N_A_45_443#_c_258_n 0.0083811f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_142 N_A_c_130_n N_A_45_443#_c_207_n 0.0311559f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_143 N_A_M1007_g N_A_45_443#_c_240_n 0.00229199f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_144 N_A_M1019_g N_A_45_443#_c_240_n 0.0125891f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_145 A N_A_45_443#_c_240_n 0.0112571f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_146 N_A_c_130_n N_A_45_443#_c_240_n 0.00355898f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_147 N_A_c_128_n N_A_45_443#_c_265_n 0.0156753f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_148 A N_A_45_443#_c_265_n 0.00887026f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_149 N_A_c_130_n N_A_45_443#_c_265_n 0.00269586f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_150 A N_A_45_443#_c_268_n 0.0152738f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A_c_130_n N_A_45_443#_c_268_n 0.0154167f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_152 N_A_c_130_n N_A_45_443#_c_209_n 0.0206085f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_153 N_A_M1007_g N_VPWR_c_464_n 0.0103088f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_154 N_A_M1019_g N_VPWR_c_464_n 0.0156302f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_155 N_A_M1019_g N_VPWR_c_478_n 0.00249815f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_156 N_A_M1007_g N_VPWR_c_502_n 7.78697e-19 $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_157 N_A_M1019_g N_VPWR_c_502_n 0.030772f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_158 N_A_M1006_g N_VPWR_c_490_n 0.0716973f $X=0.76 $Y=2.965 $X2=0 $Y2=0
cc_159 N_A_M1007_g N_VPWR_c_490_n 0.0862897f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_160 N_A_M1019_g N_VPWR_c_490_n 0.00121482f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_161 N_A_M1006_g N_VPWR_c_496_n 0.00951892f $X=0.76 $Y=2.965 $X2=0 $Y2=0
cc_162 N_A_M1007_g N_VPWR_c_496_n 0.010513f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_163 N_A_M1019_g N_VPWR_c_496_n 0.010744f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_164 N_A_c_128_n N_noxref_6_c_608_n 0.00217811f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_165 N_A_c_128_n N_noxref_6_c_613_n 0.00142024f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_166 A N_noxref_6_c_613_n 4.32971e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_167 N_A_c_127_n N_VGND_c_772_n 0.00367492f $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_168 N_A_c_128_n N_VGND_c_772_n 0.00793008f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_169 N_A_c_124_n N_VGND_c_774_n 0.0572185f $X=0.78 $Y=1.565 $X2=0 $Y2=0
cc_170 N_A_c_126_n N_VGND_c_774_n 0.00914385f $X=1.57 $Y=1.815 $X2=0 $Y2=0
cc_171 N_A_c_127_n N_VGND_c_774_n 0.0624373f $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_172 N_A_c_128_n N_VGND_c_774_n 6.48731e-19 $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_173 A N_VGND_c_774_n 0.0836537f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_174 N_A_c_127_n N_VGND_c_776_n 4.13084e-19 $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_175 N_A_c_128_n N_VGND_c_776_n 0.0408201f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_176 N_A_c_124_n N_VGND_c_787_n 0.00915616f $X=0.78 $Y=1.565 $X2=0 $Y2=0
cc_177 N_A_c_127_n N_VGND_c_787_n 0.00865748f $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_178 N_A_c_128_n N_VGND_c_787_n 0.00795556f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_179 N_A_45_443#_c_237_n N_VPWR_M1006_d 0.00539862f $X=2.045 $Y=2.18 $X2=0
+ $Y2=0
cc_180 N_A_45_443#_M1007_s N_VPWR_c_464_n 8.28689e-19 $X=2.07 $Y=2.215 $X2=0
+ $Y2=0
cc_181 N_A_45_443#_c_252_n N_VPWR_c_464_n 0.0314378f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_182 N_A_45_443#_c_210_n N_VPWR_c_467_n 0.00981852f $X=3.38 $Y=2.105 $X2=4.8
+ $Y2=0
cc_183 N_A_45_443#_c_213_n N_VPWR_c_467_n 0.00984257f $X=4.16 $Y=2.105 $X2=4.8
+ $Y2=0
cc_184 N_A_45_443#_c_216_n N_VPWR_c_470_n 0.00984257f $X=4.94 $Y=2.105 $X2=4.8
+ $Y2=0.057
cc_185 N_A_45_443#_c_219_n N_VPWR_c_470_n 0.00984257f $X=5.72 $Y=2.105 $X2=4.8
+ $Y2=0.057
cc_186 N_A_45_443#_c_222_n N_VPWR_c_473_n 0.00984257f $X=6.5 $Y=2.105 $X2=4.8
+ $Y2=0.058
cc_187 N_A_45_443#_c_225_n N_VPWR_c_473_n 0.00984257f $X=7.28 $Y=2.105 $X2=4.8
+ $Y2=0.058
cc_188 N_A_45_443#_c_228_n N_VPWR_c_476_n 7.80614e-19 $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_189 N_A_45_443#_c_231_n N_VPWR_c_476_n 0.014504f $X=8.84 $Y=2.105 $X2=0 $Y2=0
cc_190 N_A_45_443#_c_210_n N_VPWR_c_478_n 0.00656115f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_191 N_A_45_443#_c_213_n N_VPWR_c_481_n 0.00656544f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_192 N_A_45_443#_c_216_n N_VPWR_c_481_n 0.00656544f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_193 N_A_45_443#_c_219_n N_VPWR_c_484_n 0.00656544f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_194 N_A_45_443#_c_222_n N_VPWR_c_484_n 0.00656544f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_195 N_A_45_443#_c_225_n N_VPWR_c_487_n 0.00656544f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_196 N_A_45_443#_c_228_n N_VPWR_c_487_n 0.00656544f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_197 N_A_45_443#_c_210_n N_VPWR_c_502_n 0.0595501f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_198 N_A_45_443#_c_213_n N_VPWR_c_502_n 4.52391e-19 $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_199 N_A_45_443#_c_252_n N_VPWR_c_502_n 0.0873251f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_200 N_A_45_443#_c_207_n N_VPWR_c_502_n 0.0223037f $X=3.295 $Y=1.79 $X2=0
+ $Y2=0
cc_201 N_A_45_443#_c_210_n N_VPWR_c_532_n 4.54877e-19 $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_202 N_A_45_443#_c_213_n N_VPWR_c_532_n 0.0549628f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_203 N_A_45_443#_c_216_n N_VPWR_c_532_n 0.0549628f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_204 N_A_45_443#_c_219_n N_VPWR_c_532_n 4.54877e-19 $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_205 N_A_45_443#_c_209_n N_VPWR_c_532_n 5.92537e-19 $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_206 N_A_45_443#_c_216_n N_VPWR_c_537_n 4.54877e-19 $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_207 N_A_45_443#_c_219_n N_VPWR_c_537_n 0.0549628f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_208 N_A_45_443#_c_222_n N_VPWR_c_537_n 0.0567237f $X=6.5 $Y=2.105 $X2=0 $Y2=0
cc_209 N_A_45_443#_c_225_n N_VPWR_c_537_n 4.54877e-19 $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_210 N_A_45_443#_c_209_n N_VPWR_c_537_n 5.92537e-19 $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_211 N_A_45_443#_c_222_n N_VPWR_c_542_n 4.54877e-19 $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_212 N_A_45_443#_c_225_n N_VPWR_c_542_n 0.0569865f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_213 N_A_45_443#_c_228_n N_VPWR_c_542_n 0.0581256f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_214 N_A_45_443#_c_231_n N_VPWR_c_542_n 0.0011619f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_215 N_A_45_443#_c_209_n N_VPWR_c_542_n 6.12604e-19 $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_216 N_A_45_443#_c_235_n N_VPWR_c_490_n 0.0817667f $X=0.35 $Y=2.36 $X2=0 $Y2=0
cc_217 N_A_45_443#_c_237_n N_VPWR_c_490_n 0.0847738f $X=2.045 $Y=2.18 $X2=0
+ $Y2=0
cc_218 N_A_45_443#_c_252_n N_VPWR_c_490_n 0.0787997f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_219 N_A_45_443#_c_228_n N_VPWR_c_493_n 0.0098265f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_220 N_A_45_443#_c_231_n N_VPWR_c_493_n 0.0115186f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_221 N_A_45_443#_M1006_s N_VPWR_c_496_n 0.00425071f $X=0.225 $Y=2.215 $X2=0
+ $Y2=0
cc_222 N_A_45_443#_c_210_n N_VPWR_c_496_n 0.00967409f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_223 N_A_45_443#_c_213_n N_VPWR_c_496_n 0.00966853f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_224 N_A_45_443#_c_216_n N_VPWR_c_496_n 0.00966853f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_225 N_A_45_443#_c_219_n N_VPWR_c_496_n 0.00966853f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_226 N_A_45_443#_c_222_n N_VPWR_c_496_n 0.00994001f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_227 N_A_45_443#_c_225_n N_VPWR_c_496_n 0.00994001f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_228 N_A_45_443#_c_228_n N_VPWR_c_496_n 0.00989505f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_229 N_A_45_443#_c_231_n N_VPWR_c_496_n 0.0107477f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_230 N_A_45_443#_c_235_n N_VPWR_c_496_n 0.0196936f $X=0.35 $Y=2.36 $X2=0 $Y2=0
cc_231 N_A_45_443#_c_252_n N_VPWR_c_496_n 0.0205648f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_232 N_A_45_443#_c_210_n N_noxref_6_c_615_n 0.0234771f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_233 N_A_45_443#_c_213_n N_noxref_6_c_615_n 0.0234771f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_234 N_A_45_443#_M1001_g N_noxref_6_c_604_n 0.00440473f $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_235 N_A_45_443#_M1002_g N_noxref_6_c_604_n 0.00441377f $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_236 N_A_45_443#_c_209_n N_noxref_6_c_604_n 0.00432417f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_237 N_A_45_443#_c_209_n N_noxref_6_c_620_n 0.0615828f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_238 N_A_45_443#_c_207_n N_noxref_6_c_621_n 0.00900397f $X=3.295 $Y=1.79 $X2=0
+ $Y2=0
cc_239 N_A_45_443#_c_209_n N_noxref_6_c_621_n 0.00843233f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_240 N_A_45_443#_c_213_n N_noxref_6_c_609_n 0.0156902f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_241 N_A_45_443#_c_216_n N_noxref_6_c_609_n 0.0156902f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_242 N_A_45_443#_c_209_n N_noxref_6_c_609_n 0.0245717f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_243 N_A_45_443#_c_210_n N_noxref_6_c_626_n 0.00529873f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_244 N_A_45_443#_c_213_n N_noxref_6_c_626_n 0.00141551f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_245 N_A_45_443#_c_209_n N_noxref_6_c_626_n 0.01313f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_246 N_A_45_443#_c_216_n N_noxref_6_c_629_n 0.0234771f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_247 N_A_45_443#_c_219_n N_noxref_6_c_629_n 0.0232569f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_248 N_A_45_443#_M1009_g N_noxref_6_c_605_n 0.00441377f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_249 N_A_45_443#_M1013_g N_noxref_6_c_605_n 0.00441377f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_250 N_A_45_443#_c_209_n N_noxref_6_c_605_n 0.00437511f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_251 N_A_45_443#_c_209_n N_noxref_6_c_634_n 0.0644185f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_252 N_A_45_443#_c_219_n N_noxref_6_c_610_n 0.0121299f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_253 N_A_45_443#_c_222_n N_noxref_6_c_610_n 0.0120576f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_254 N_A_45_443#_c_209_n N_noxref_6_c_610_n 0.0224309f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_255 N_A_45_443#_c_222_n N_noxref_6_c_638_n 0.0250679f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_256 N_A_45_443#_c_225_n N_noxref_6_c_638_n 0.0252769f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_257 N_A_45_443#_M1014_g N_noxref_6_c_606_n 0.00400399f $X=6.5 $Y=1.08 $X2=0
+ $Y2=0
cc_258 N_A_45_443#_M1018_g N_noxref_6_c_606_n 0.00400399f $X=7.28 $Y=1.08 $X2=0
+ $Y2=0
cc_259 N_A_45_443#_c_209_n N_noxref_6_c_606_n 0.00455707f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_260 N_A_45_443#_c_209_n N_noxref_6_c_643_n 0.078465f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_261 N_A_45_443#_c_228_n N_noxref_6_c_644_n 0.0094348f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_262 N_A_45_443#_c_231_n N_noxref_6_c_644_n 0.0275957f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_263 N_A_45_443#_c_228_n N_noxref_6_c_646_n 0.0176022f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_264 N_A_45_443#_c_231_n N_noxref_6_c_646_n 0.0363847f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_265 N_A_45_443#_M1020_g N_noxref_6_c_607_n 0.00400399f $X=8.06 $Y=1.08 $X2=0
+ $Y2=0
cc_266 N_A_45_443#_M1021_g N_noxref_6_c_607_n 0.00133825f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_267 N_A_45_443#_c_209_n N_noxref_6_c_607_n 0.00399266f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_268 N_A_45_443#_M1021_g N_noxref_6_c_651_n 0.0183266f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_269 N_A_45_443#_M1021_g N_noxref_6_c_652_n 0.0291857f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_270 N_A_45_443#_c_209_n N_noxref_6_c_652_n 0.0394165f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_271 N_A_45_443#_c_216_n N_noxref_6_c_654_n 0.00141551f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_272 N_A_45_443#_c_219_n N_noxref_6_c_654_n 0.00141551f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_273 N_A_45_443#_c_209_n N_noxref_6_c_654_n 0.00854953f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_274 N_A_45_443#_c_209_n N_noxref_6_c_657_n 0.00585522f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_275 N_A_45_443#_c_222_n N_noxref_6_c_658_n 0.00141551f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_276 N_A_45_443#_c_225_n N_noxref_6_c_658_n 0.00141551f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_277 N_A_45_443#_c_209_n N_noxref_6_c_658_n 0.00807226f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_278 N_A_45_443#_c_209_n N_noxref_6_c_661_n 0.00630631f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_279 N_A_45_443#_c_225_n N_noxref_6_c_611_n 0.0133649f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_280 N_A_45_443#_c_228_n N_noxref_6_c_611_n 0.0173368f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_281 N_A_45_443#_c_209_n N_noxref_6_c_611_n 0.0268604f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_282 N_A_45_443#_c_228_n N_noxref_6_c_665_n 0.00141551f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_283 N_A_45_443#_c_231_n N_noxref_6_c_665_n 0.00911503f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_284 N_A_45_443#_c_209_n N_noxref_6_c_665_n 0.0234141f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_285 N_A_45_443#_c_222_n N_noxref_6_c_668_n 0.0119036f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_286 N_A_45_443#_c_225_n N_noxref_6_c_668_n 0.0088113f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_287 N_A_45_443#_c_209_n N_noxref_6_c_668_n 0.0160657f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_288 N_A_45_443#_c_219_n N_noxref_6_c_671_n 0.00902392f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_289 N_A_45_443#_c_209_n N_noxref_6_c_671_n 0.0103187f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_290 N_A_45_443#_c_209_n N_noxref_6_c_673_n 0.00270744f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_291 N_A_45_443#_M1001_g N_noxref_6_c_608_n 0.00360335f $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_292 N_A_45_443#_c_210_n N_noxref_6_c_608_n 0.00529116f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_293 N_A_45_443#_M1002_g N_noxref_6_c_608_n 0.00204637f $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_294 N_A_45_443#_c_213_n N_noxref_6_c_608_n 0.00234371f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_295 N_A_45_443#_M1009_g N_noxref_6_c_608_n 0.00204637f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_296 N_A_45_443#_c_216_n N_noxref_6_c_608_n 0.00234371f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_297 N_A_45_443#_M1013_g N_noxref_6_c_608_n 0.00176874f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_298 N_A_45_443#_c_219_n N_noxref_6_c_608_n 0.00206235f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_299 N_A_45_443#_M1014_g N_noxref_6_c_608_n 8.02658e-19 $X=6.5 $Y=1.08 $X2=0
+ $Y2=0
cc_300 N_A_45_443#_c_222_n N_noxref_6_c_608_n 7.33013e-19 $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_301 N_A_45_443#_c_252_n N_noxref_6_c_608_n 0.00164841f $X=2.21 $Y=2.34 $X2=0
+ $Y2=0
cc_302 N_A_45_443#_c_254_n N_noxref_6_c_608_n 0.0013506f $X=2.51 $Y=1.625 $X2=0
+ $Y2=0
cc_303 N_A_45_443#_c_258_n N_noxref_6_c_608_n 9.16329e-19 $X=2.51 $Y=2.095 $X2=0
+ $Y2=0
cc_304 N_A_45_443#_c_207_n N_noxref_6_c_608_n 0.0024863f $X=3.295 $Y=1.79 $X2=0
+ $Y2=0
cc_305 N_A_45_443#_c_240_n N_noxref_6_c_608_n 0.00162285f $X=2.32 $Y=2.18 $X2=0
+ $Y2=0
cc_306 N_A_45_443#_c_209_n N_noxref_6_c_608_n 0.00843505f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_307 N_A_45_443#_M1001_g N_noxref_6_c_613_n 0.00435634f $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_308 N_A_45_443#_c_210_n N_noxref_6_c_613_n 0.00429145f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_309 N_A_45_443#_M1002_g N_noxref_6_c_613_n 0.00191064f $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_310 N_A_45_443#_M1009_g N_noxref_6_c_613_n 0.00191064f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_311 N_A_45_443#_M1013_g N_noxref_6_c_613_n 0.00191064f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_312 N_A_45_443#_M1014_g N_noxref_6_c_613_n 0.00274535f $X=6.5 $Y=1.08 $X2=0
+ $Y2=0
cc_313 N_A_45_443#_c_222_n N_noxref_6_c_613_n 0.00254426f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_314 N_A_45_443#_c_252_n N_noxref_6_c_613_n 0.00165664f $X=2.21 $Y=2.34 $X2=0
+ $Y2=0
cc_315 N_A_45_443#_c_254_n N_noxref_6_c_613_n 0.00141076f $X=2.51 $Y=1.625 $X2=0
+ $Y2=0
cc_316 N_A_45_443#_c_258_n N_noxref_6_c_613_n 0.00102155f $X=2.51 $Y=2.095 $X2=0
+ $Y2=0
cc_317 N_A_45_443#_c_207_n N_noxref_6_c_613_n 0.00734543f $X=3.295 $Y=1.79 $X2=0
+ $Y2=0
cc_318 N_A_45_443#_c_240_n N_noxref_6_c_613_n 0.00165668f $X=2.32 $Y=2.18 $X2=0
+ $Y2=0
cc_319 N_A_45_443#_c_265_n N_noxref_6_c_613_n 3.7935e-19 $X=2.51 $Y=1.315 $X2=0
+ $Y2=0
cc_320 N_A_45_443#_c_209_n N_noxref_6_c_613_n 0.00949279f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_321 N_A_45_443#_c_209_n N_noxref_6_c_704_n 0.00660997f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_322 N_A_45_443#_c_219_n N_noxref_6_c_705_n 0.0110025f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_323 N_A_45_443#_c_209_n N_noxref_6_c_705_n 0.0205876f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_324 N_A_45_443#_c_416_p N_VGND_c_772_n 0.0122346f $X=2.21 $Y=0.895 $X2=0
+ $Y2=0
cc_325 N_A_45_443#_M1021_g N_VGND_c_773_n 0.00589056f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_326 N_A_45_443#_c_244_n N_VGND_c_774_n 0.0377885f $X=0.37 $Y=0.97 $X2=0 $Y2=0
cc_327 N_A_45_443#_M1001_g N_VGND_c_776_n 0.0552367f $X=3.38 $Y=1.08 $X2=0 $Y2=0
cc_328 N_A_45_443#_M1002_g N_VGND_c_776_n 0.00107004f $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_329 N_A_45_443#_c_254_n N_VGND_c_776_n 0.00342789f $X=2.51 $Y=1.625 $X2=0
+ $Y2=0
cc_330 N_A_45_443#_c_207_n N_VGND_c_776_n 0.0437936f $X=3.295 $Y=1.79 $X2=0
+ $Y2=0
cc_331 N_A_45_443#_c_265_n N_VGND_c_776_n 0.0138755f $X=2.51 $Y=1.315 $X2=0
+ $Y2=0
cc_332 N_A_45_443#_M1001_g N_VGND_c_778_n 0.00328808f $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_333 N_A_45_443#_M1002_g N_VGND_c_778_n 0.00328808f $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_334 N_A_45_443#_M1001_g N_VGND_c_780_n 0.00106904f $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_335 N_A_45_443#_M1002_g N_VGND_c_780_n 0.0510174f $X=4.16 $Y=1.08 $X2=0 $Y2=0
cc_336 N_A_45_443#_M1009_g N_VGND_c_780_n 0.0510174f $X=4.94 $Y=1.08 $X2=0 $Y2=0
cc_337 N_A_45_443#_M1013_g N_VGND_c_780_n 0.00106904f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_338 N_A_45_443#_c_209_n N_VGND_c_780_n 0.00244164f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_339 N_A_45_443#_M1009_g N_VGND_c_781_n 0.00328808f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_340 N_A_45_443#_M1013_g N_VGND_c_781_n 0.00328808f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_341 N_A_45_443#_M1009_g N_VGND_c_782_n 0.00106904f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_342 N_A_45_443#_M1013_g N_VGND_c_782_n 0.0510174f $X=5.72 $Y=1.08 $X2=0 $Y2=0
cc_343 N_A_45_443#_M1014_g N_VGND_c_782_n 0.0523853f $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_344 N_A_45_443#_M1018_g N_VGND_c_782_n 9.10934e-19 $X=7.28 $Y=1.08 $X2=0
+ $Y2=0
cc_345 N_A_45_443#_c_209_n N_VGND_c_782_n 0.00244164f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_346 N_A_45_443#_M1014_g N_VGND_c_783_n 0.00328808f $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_347 N_A_45_443#_M1018_g N_VGND_c_783_n 0.00328808f $X=7.28 $Y=1.08 $X2=0
+ $Y2=0
cc_348 N_A_45_443#_M1014_g N_VGND_c_784_n 9.10934e-19 $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_349 N_A_45_443#_M1018_g N_VGND_c_784_n 0.0525581f $X=7.28 $Y=1.08 $X2=0 $Y2=0
cc_350 N_A_45_443#_M1020_g N_VGND_c_784_n 0.0532979f $X=8.06 $Y=1.08 $X2=0 $Y2=0
cc_351 N_A_45_443#_M1021_g N_VGND_c_784_n 0.00130456f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_352 N_A_45_443#_c_209_n N_VGND_c_784_n 0.00257674f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_353 N_A_45_443#_M1020_g N_VGND_c_785_n 0.00520463f $X=8.06 $Y=1.08 $X2=0
+ $Y2=0
cc_354 N_A_45_443#_M1021_g N_VGND_c_785_n 0.00965248f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_355 N_A_45_443#_M1021_g N_VGND_c_786_n 0.00617584f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_356 N_A_45_443#_M1001_g N_VGND_c_787_n 0.00739524f $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_357 N_A_45_443#_M1002_g N_VGND_c_787_n 0.00739524f $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_358 N_A_45_443#_M1009_g N_VGND_c_787_n 0.00739524f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_359 N_A_45_443#_M1013_g N_VGND_c_787_n 0.00739524f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_360 N_A_45_443#_M1014_g N_VGND_c_787_n 0.00808151f $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_361 N_A_45_443#_M1018_g N_VGND_c_787_n 0.00808151f $X=7.28 $Y=1.08 $X2=0
+ $Y2=0
cc_362 N_A_45_443#_M1020_g N_VGND_c_787_n 0.00808151f $X=8.06 $Y=1.08 $X2=0
+ $Y2=0
cc_363 N_A_45_443#_M1021_g N_VGND_c_787_n 0.0148456f $X=8.84 $Y=1.08 $X2=0 $Y2=0
cc_364 N_A_45_443#_c_244_n N_VGND_c_787_n 0.0118041f $X=0.37 $Y=0.97 $X2=0 $Y2=0
cc_365 N_A_45_443#_c_416_p N_VGND_c_787_n 0.00689067f $X=2.21 $Y=0.895 $X2=0
+ $Y2=0
cc_366 N_A_45_443#_c_265_n N_VGND_c_787_n 0.00762664f $X=2.51 $Y=1.315 $X2=0
+ $Y2=0
cc_367 N_A_45_443#_c_210_n X 0.0023443f $X=3.38 $Y=2.105 $X2=0 $Y2=0
cc_368 N_A_45_443#_c_213_n X 0.0023443f $X=4.16 $Y=2.105 $X2=0 $Y2=0
cc_369 N_A_45_443#_c_216_n X 0.0023443f $X=4.94 $Y=2.105 $X2=0 $Y2=0
cc_370 N_A_45_443#_c_219_n X 0.0023443f $X=5.72 $Y=2.105 $X2=0 $Y2=0
cc_371 N_A_45_443#_c_252_n X 4.88711e-19 $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_372 N_VPWR_c_467_n N_noxref_6_M1000_d 8.28689e-19 $X=4.105 $Y=3.71 $X2=0
+ $Y2=0
cc_373 N_VPWR_c_470_n N_noxref_6_M1005_d 8.28689e-19 $X=5.665 $Y=3.71 $X2=0
+ $Y2=3.955
cc_374 N_VPWR_c_473_n N_noxref_6_M1011_d 8.28689e-19 $X=7.225 $Y=3.71 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_493_n N_noxref_6_M1016_d 8.28689e-19 $X=8.905 $Y=3.635 $X2=0.24
+ $Y2=4.07
cc_376 N_VPWR_c_467_n N_noxref_6_c_615_n 0.0178796f $X=4.105 $Y=3.71 $X2=0 $Y2=0
cc_377 N_VPWR_c_502_n N_noxref_6_c_615_n 0.0839169f $X=2.99 $Y=2.55 $X2=0 $Y2=0
cc_378 N_VPWR_c_532_n N_noxref_6_c_615_n 0.0840214f $X=4.55 $Y=2.55 $X2=0 $Y2=0
cc_379 N_VPWR_c_496_n N_noxref_6_c_615_n 0.01238f $X=9.35 $Y=3.56 $X2=0 $Y2=0
cc_380 N_VPWR_c_532_n N_noxref_6_c_609_n 0.0644067f $X=4.55 $Y=2.55 $X2=0 $Y2=0
cc_381 N_VPWR_c_470_n N_noxref_6_c_629_n 0.0178796f $X=5.665 $Y=3.71 $X2=0 $Y2=0
cc_382 N_VPWR_c_532_n N_noxref_6_c_629_n 0.0840214f $X=4.55 $Y=2.55 $X2=0 $Y2=0
cc_383 N_VPWR_c_537_n N_noxref_6_c_629_n 0.0840214f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_384 N_VPWR_c_496_n N_noxref_6_c_629_n 0.01238f $X=9.35 $Y=3.56 $X2=0 $Y2=0
cc_385 N_VPWR_c_537_n N_noxref_6_c_610_n 0.0593743f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_386 N_VPWR_c_473_n N_noxref_6_c_638_n 0.0178796f $X=7.225 $Y=3.71 $X2=0 $Y2=0
cc_387 N_VPWR_c_537_n N_noxref_6_c_638_n 0.0842143f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_388 N_VPWR_c_542_n N_noxref_6_c_638_n 0.0842143f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_389 N_VPWR_c_496_n N_noxref_6_c_638_n 0.01238f $X=9.35 $Y=3.56 $X2=0 $Y2=0
cc_390 N_VPWR_c_476_n N_noxref_6_c_644_n 0.0026211f $X=9.32 $Y=3.475 $X2=0 $Y2=0
cc_391 N_VPWR_c_542_n N_noxref_6_c_644_n 0.0462063f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_392 N_VPWR_c_493_n N_noxref_6_c_644_n 0.0292853f $X=8.905 $Y=3.635 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_496_n N_noxref_6_c_644_n 0.0232887f $X=9.35 $Y=3.56 $X2=0 $Y2=0
cc_394 N_VPWR_c_542_n N_noxref_6_c_646_n 0.0422929f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_395 N_VPWR_c_542_n N_noxref_6_c_611_n 0.0605198f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_396 N_VPWR_M1010_s N_noxref_6_c_668_n 0.00281468f $X=5.97 $Y=2.215 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_542_n N_noxref_6_c_668_n 0.00221579f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_398 N_VPWR_M1010_s N_noxref_6_c_671_n 6.57737e-19 $X=5.97 $Y=2.215 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_537_n N_noxref_6_c_671_n 0.0211813f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_400 N_VPWR_M1010_s N_noxref_6_c_673_n 0.00194331f $X=5.97 $Y=2.215 $X2=0
+ $Y2=0
cc_401 N_VPWR_M1010_s N_noxref_6_c_608_n 0.00170316f $X=5.97 $Y=2.215 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_502_n N_noxref_6_c_608_n 0.00255084f $X=2.99 $Y=2.55 $X2=0 $Y2=0
cc_403 N_VPWR_c_532_n N_noxref_6_c_608_n 0.0149797f $X=4.55 $Y=2.55 $X2=0 $Y2=0
cc_404 N_VPWR_c_537_n N_noxref_6_c_608_n 0.010022f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_405 N_VPWR_c_502_n N_noxref_6_c_613_n 0.00443935f $X=2.99 $Y=2.55 $X2=0 $Y2=0
cc_406 N_VPWR_c_532_n N_noxref_6_c_613_n 2.2199e-19 $X=4.55 $Y=2.55 $X2=0 $Y2=0
cc_407 N_VPWR_c_537_n N_noxref_6_c_613_n 0.00411589f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_408 N_VPWR_M1010_s N_noxref_6_c_705_n 0.00403395f $X=5.97 $Y=2.215 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_502_n X 0.00592951f $X=2.99 $Y=2.55 $X2=0 $Y2=3.985
cc_410 N_VPWR_c_532_n X 0.0134543f $X=4.55 $Y=2.55 $X2=0 $Y2=3.985
cc_411 N_VPWR_c_537_n X 0.0130519f $X=6.11 $Y=2.55 $X2=0 $Y2=3.985
cc_412 N_VPWR_c_496_n X 0.030685f $X=9.35 $Y=3.56 $X2=0 $Y2=3.985
cc_413 N_noxref_6_c_604_n N_VGND_c_776_n 0.0309863f $X=3.77 $Y=0.97 $X2=0 $Y2=0
cc_414 N_noxref_6_c_608_n N_VGND_c_776_n 0.00286772f $X=5.6 $Y=1.945 $X2=0 $Y2=0
cc_415 N_noxref_6_c_613_n N_VGND_c_776_n 0.00715684f $X=5.6 $Y=1.945 $X2=0 $Y2=0
cc_416 N_noxref_6_c_604_n N_VGND_c_778_n 0.0086879f $X=3.77 $Y=0.97 $X2=0 $Y2=0
cc_417 N_noxref_6_c_604_n N_VGND_c_780_n 0.0309252f $X=3.77 $Y=0.97 $X2=0 $Y2=0
cc_418 N_noxref_6_c_620_n N_VGND_c_780_n 0.0719426f $X=5.225 $Y=1.71 $X2=0 $Y2=0
cc_419 N_noxref_6_c_605_n N_VGND_c_780_n 0.0309252f $X=5.33 $Y=0.97 $X2=0 $Y2=0
cc_420 N_noxref_6_c_608_n N_VGND_c_780_n 0.014978f $X=5.6 $Y=1.945 $X2=0 $Y2=0
cc_421 N_noxref_6_c_613_n N_VGND_c_780_n 0.015949f $X=5.6 $Y=1.945 $X2=0 $Y2=0
cc_422 N_noxref_6_c_605_n N_VGND_c_781_n 0.0086879f $X=5.33 $Y=0.97 $X2=0 $Y2=0
cc_423 N_noxref_6_c_605_n N_VGND_c_782_n 0.0309252f $X=5.33 $Y=0.97 $X2=0 $Y2=0
cc_424 N_noxref_6_c_634_n N_VGND_c_782_n 0.0710502f $X=6.785 $Y=1.71 $X2=0 $Y2=0
cc_425 N_noxref_6_c_608_n N_VGND_c_782_n 0.00935962f $X=5.6 $Y=1.945 $X2=0 $Y2=0
cc_426 N_noxref_6_c_613_n N_VGND_c_782_n 0.0146975f $X=5.6 $Y=1.945 $X2=0 $Y2=0
cc_427 N_noxref_6_c_606_n N_VGND_c_783_n 0.0086879f $X=6.89 $Y=0.97 $X2=0 $Y2=0
cc_428 N_noxref_6_c_643_n N_VGND_c_784_n 0.0685594f $X=8.345 $Y=1.71 $X2=0 $Y2=0
cc_429 N_noxref_6_c_760_p N_VGND_c_785_n 0.00873551f $X=8.45 $Y=0.975 $X2=0
+ $Y2=0
cc_430 N_noxref_6_c_651_n N_VGND_c_785_n 0.0168514f $X=8.735 $Y=0.89 $X2=0 $Y2=0
cc_431 N_noxref_6_c_604_n N_VGND_c_787_n 0.00668507f $X=3.77 $Y=0.97 $X2=0 $Y2=0
cc_432 N_noxref_6_c_605_n N_VGND_c_787_n 0.00668507f $X=5.33 $Y=0.97 $X2=0 $Y2=0
cc_433 N_noxref_6_c_606_n N_VGND_c_787_n 0.00668507f $X=6.89 $Y=0.97 $X2=0 $Y2=0
cc_434 N_noxref_6_c_760_p N_VGND_c_787_n 0.00674935f $X=8.45 $Y=0.975 $X2=0
+ $Y2=0
cc_435 N_noxref_6_c_651_n N_VGND_c_787_n 0.011179f $X=8.735 $Y=0.89 $X2=0 $Y2=0
cc_436 N_noxref_6_c_608_n N_VGND_c_787_n 0.0407576f $X=5.6 $Y=1.945 $X2=0 $Y2=0
cc_437 N_noxref_6_c_613_n N_VGND_c_787_n 0.0463638f $X=5.6 $Y=1.945 $X2=0 $Y2=0
cc_438 N_noxref_6_c_615_n X 0.00515769f $X=3.77 $Y=2.34 $X2=0 $Y2=0
cc_439 N_noxref_6_c_629_n X 0.00515769f $X=5.33 $Y=2.34 $X2=0 $Y2=0
cc_440 N_noxref_6_c_638_n X 5.06817e-19 $X=6.89 $Y=2.34 $X2=0 $Y2=0
