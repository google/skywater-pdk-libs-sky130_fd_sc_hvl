* File: sky130_fd_sc_hvl__dfstp_1.pex.spice
* Created: Wed Sep  2 09:05:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%VNB 5 7 11
r102 7 11 0.000478831 $w=1.488e-05 $l=5.7e-08 $layer=MET1_cond $X=7.44 $Y=0.057
+ $X2=7.44 $Y2=0
r103 5 11 0.6 $w=1.7e-07 $l=2.635e-06 $layer=mcon $count=15 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r104 5 11 0.6 $w=1.7e-07 $l=2.635e-06 $layer=mcon $count=15 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%VPB 4 6 14
r153 10 14 0.6 $w=1.7e-07 $l=2.635e-06 $layer=mcon $count=15 $X=14.64 $Y=4.07
+ $X2=14.64 $Y2=4.07
r154 9 14 939.465 $w=1.68e-07 $l=1.44e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=14.64 $Y2=4.07
r155 9 10 0.6 $w=1.7e-07 $l=2.635e-06 $layer=mcon $count=15 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r156 6 10 0.000478831 $w=1.488e-05 $l=5.7e-08 $layer=MET1_cond $X=7.44 $Y=4.013
+ $X2=7.44 $Y2=4.07
r157 4 14 11.7419 $w=1.7e-07 $l=1.46824e-05 $layer=licon1_NTAP_notbjt $count=15
+ $X=0 $Y=3.985 $X2=14.64 $Y2=4.07
r158 4 9 11.7419 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=15
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%CLK 3 7 9 12
r27 12 15 21.8167 $w=5.15e-07 $l=2.1e-07 $layer=POLY_cond $X=0.677 $Y=2.24
+ $X2=0.677 $Y2=2.45
r28 12 14 30.1279 $w=5.15e-07 $l=2.9e-07 $layer=POLY_cond $X=0.677 $Y=2.24
+ $X2=0.677 $Y2=1.95
r29 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.71
+ $Y=2.24 $X2=0.71 $Y2=2.24
r30 9 13 0.178519 $w=6.68e-07 $l=1e-08 $layer=LI1_cond $X=0.72 $Y=2.41 $X2=0.71
+ $Y2=2.41
r31 7 14 116.101 $w=5e-07 $l=1.085e-06 $layer=POLY_cond $X=0.685 $Y=0.865
+ $X2=0.685 $Y2=1.95
r32 3 15 95.2352 $w=5e-07 $l=8.9e-07 $layer=POLY_cond $X=0.67 $Y=3.34 $X2=0.67
+ $Y2=2.45
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%A_30_131# 1 2 9 13 17 18 20 23 27 31 33 38
+ 39 40 42 43 44 46 47 48 51 54 58 60 61 62 63 65 67 68 69 70 75 76 81 89
c240 89 0 1.48283e-19 $X=4.645 $Y=3.175
c241 76 0 1.92639e-19 $X=8.795 $Y=2.25
c242 51 0 3.85523e-20 $X=3.8 $Y=1.25
c243 39 0 1.1261e-19 $X=2.12 $Y=0.35
r244 76 93 92.4947 $w=4.69e-07 $l=9e-07 $layer=POLY_cond $X=8.795 $Y=2.12
+ $X2=9.695 $Y2=2.12
r245 76 91 7.19403 $w=4.69e-07 $l=7e-08 $layer=POLY_cond $X=8.795 $Y=2.12
+ $X2=8.725 $Y2=2.12
r246 75 78 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=8.795 $Y=2.25
+ $X2=8.795 $Y2=2.41
r247 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.795
+ $Y=2.25 $X2=8.795 $Y2=2.25
r248 70 72 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.55 $Y=2.24
+ $X2=6.55 $Y2=2.41
r249 68 87 51.252 $w=5.55e-07 $l=5.25e-07 $layer=POLY_cond $X=1.437 $Y=1.425
+ $X2=1.437 $Y2=1.95
r250 68 86 21.8495 $w=5.55e-07 $l=2.2e-07 $layer=POLY_cond $X=1.437 $Y=1.425
+ $X2=1.437 $Y2=1.205
r251 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.345
+ $Y=1.425 $X2=1.345 $Y2=1.425
r252 64 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.635 $Y=2.41
+ $X2=6.55 $Y2=2.41
r253 63 78 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.63 $Y=2.41
+ $X2=8.795 $Y2=2.41
r254 63 64 130.155 $w=1.68e-07 $l=1.995e-06 $layer=LI1_cond $X=8.63 $Y=2.41
+ $X2=6.635 $Y2=2.41
r255 61 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.465 $Y=2.24
+ $X2=6.55 $Y2=2.24
r256 61 62 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=6.465 $Y=2.24
+ $X2=5.005 $Y2=2.24
r257 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.92 $Y=2.325
+ $X2=5.005 $Y2=2.24
r258 59 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.92 $Y=2.325
+ $X2=4.92 $Y2=3.285
r259 58 89 27.761 $w=5.3e-07 $l=2.75e-07 $layer=POLY_cond $X=4.645 $Y=3.45
+ $X2=4.645 $Y2=3.175
r260 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.565
+ $Y=3.45 $X2=4.565 $Y2=3.45
r261 55 69 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.885 $Y=3.45
+ $X2=3.8 $Y2=3.45
r262 55 57 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.885 $Y=3.45
+ $X2=4.565 $Y2=3.45
r263 54 60 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.835 $Y=3.45
+ $X2=4.92 $Y2=3.285
r264 54 57 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=4.835 $Y=3.45
+ $X2=4.565 $Y2=3.45
r265 52 81 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.74 $Y=1.25 $X2=3.74
+ $Y2=0.745
r266 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.8
+ $Y=1.25 $X2=3.8 $Y2=1.25
r267 49 69 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=3.285
+ $X2=3.8 $Y2=3.45
r268 49 51 132.765 $w=1.68e-07 $l=2.035e-06 $layer=LI1_cond $X=3.8 $Y=3.285
+ $X2=3.8 $Y2=1.25
r269 47 69 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.715 $Y=3.45
+ $X2=3.8 $Y2=3.45
r270 47 48 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.715 $Y=3.45
+ $X2=3.185 $Y2=3.45
r271 46 48 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.1 $Y=3.285
+ $X2=3.185 $Y2=3.45
r272 45 46 126.567 $w=1.68e-07 $l=1.94e-06 $layer=LI1_cond $X=3.1 $Y=1.345
+ $X2=3.1 $Y2=3.285
r273 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.015 $Y=1.26
+ $X2=3.1 $Y2=1.345
r274 43 44 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.015 $Y=1.26
+ $X2=2.29 $Y2=1.26
r275 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.205 $Y=1.175
+ $X2=2.29 $Y2=1.26
r276 41 42 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.205 $Y=0.435
+ $X2=2.205 $Y2=1.175
r277 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.12 $Y=0.35
+ $X2=2.205 $Y2=0.435
r278 39 40 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.12 $Y=0.35
+ $X2=1.51 $Y2=0.35
r279 38 67 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.425 $Y=1.295
+ $X2=1.345 $Y2=1.38
r280 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.425 $Y=0.435
+ $X2=1.51 $Y2=0.35
r281 37 38 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.425 $Y=0.435
+ $X2=1.425 $Y2=1.295
r282 34 65 2.87242 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=0.38 $Y=1.38
+ $X2=0.247 $Y2=1.38
r283 33 67 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.18 $Y=1.38
+ $X2=1.345 $Y2=1.38
r284 33 34 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.18 $Y=1.38 $X2=0.38
+ $Y2=1.38
r285 29 65 3.6114 $w=2.57e-07 $l=8.84308e-08 $layer=LI1_cond $X=0.24 $Y=1.465
+ $X2=0.247 $Y2=1.38
r286 29 31 75.8307 $w=2.48e-07 $l=1.645e-06 $layer=LI1_cond $X=0.24 $Y=1.465
+ $X2=0.24 $Y2=3.11
r287 25 65 3.6114 $w=2.57e-07 $l=8.5e-08 $layer=LI1_cond $X=0.247 $Y=1.295
+ $X2=0.247 $Y2=1.38
r288 25 27 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=0.247 $Y=1.295
+ $X2=0.247 $Y2=0.865
r289 21 93 1.27363 $w=5e-07 $l=3.45e-07 $layer=POLY_cond $X=9.695 $Y=1.775
+ $X2=9.695 $Y2=2.12
r290 21 23 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=9.695 $Y=1.775
+ $X2=9.695 $Y2=1.225
r291 18 91 1.27363 $w=5e-07 $l=3.45e-07 $layer=POLY_cond $X=8.725 $Y=2.465
+ $X2=8.725 $Y2=2.12
r292 18 20 58.804 $w=5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.725 $Y=2.465
+ $X2=8.725 $Y2=3.075
r293 17 89 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.66 $Y=2.855 $X2=4.66
+ $Y2=3.175
r294 13 86 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.465 $Y=0.865
+ $X2=1.465 $Y2=1.205
r295 9 87 148.738 $w=5e-07 $l=1.39e-06 $layer=POLY_cond $X=1.45 $Y=3.34 $X2=1.45
+ $Y2=1.95
r296 2 31 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.155
+ $Y=2.965 $X2=0.28 $Y2=3.11
r297 1 27 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.655 $X2=0.295 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%D 3 5 7 9
c33 3 0 1.1261e-19 $X=2.96 $Y=0.745
r34 9 12 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.67 $Y=1.64
+ $X2=2.67 $Y2=1.64
r35 5 12 62.8564 $w=7.25e-07 $l=9.53021e-07 $layer=POLY_cond $X=3.06 $Y=2.515
+ $X2=2.897 $Y2=1.64
r36 5 7 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.06 $Y=2.515 $X2=3.06
+ $Y2=2.855
r37 1 12 27.6206 $w=7.25e-07 $l=3.7518e-07 $layer=POLY_cond $X=2.96 $Y=1.295
+ $X2=2.897 $Y2=1.64
r38 1 3 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.96 $Y=1.295 $X2=2.96
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%A_340_593# 1 2 10 13 15 17 18 21 25 29 33
+ 36 38 39 41 43 46 48 49 51 52 53 55 59 60 61 65 74 76 80
c212 76 0 1.92639e-19 $X=8.785 $Y=1.71
c213 46 0 1.62708e-19 $X=8.45 $Y=1.71
c214 36 0 6.88421e-21 $X=4.535 $Y=1.805
c215 15 0 1.85301e-19 $X=8.685 $Y=1.315
c216 13 0 3.85523e-20 $X=4.54 $Y=0.745
r217 74 76 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.62 $Y=1.71
+ $X2=8.785 $Y2=1.71
r218 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.62
+ $Y=1.71 $X2=8.62 $Y2=1.71
r219 65 67 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.9 $Y=1.89 $X2=6.9
+ $Y2=2.06
r220 58 59 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=9.225 $Y=1.875
+ $X2=9.225 $Y2=2.675
r221 56 80 95.7703 $w=5e-07 $l=8.95e-07 $layer=POLY_cond $X=9.695 $Y=3.68
+ $X2=9.695 $Y2=2.785
r222 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.66
+ $Y=3.68 $X2=9.66 $Y2=3.68
r223 53 55 41.987 $w=2.08e-07 $l=7.95e-07 $layer=LI1_cond $X=8.865 $Y=3.7
+ $X2=9.66 $Y2=3.7
r224 51 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.14 $Y=2.76
+ $X2=9.225 $Y2=2.675
r225 51 52 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.14 $Y=2.76
+ $X2=8.865 $Y2=2.76
r226 49 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.14 $Y=1.79
+ $X2=9.225 $Y2=1.875
r227 49 76 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.14 $Y=1.79
+ $X2=8.785 $Y2=1.79
r228 48 53 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.78 $Y=3.595
+ $X2=8.865 $Y2=3.7
r229 47 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.78 $Y=2.845
+ $X2=8.865 $Y2=2.76
r230 47 48 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=8.78 $Y=2.845
+ $X2=8.78 $Y2=3.595
r231 46 71 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.365 $Y=1.71
+ $X2=8.365 $Y2=2.06
r232 46 74 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=8.45 $Y=1.71
+ $X2=8.62 $Y2=1.71
r233 44 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=2.06
+ $X2=6.9 $Y2=2.06
r234 43 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.28 $Y=2.06
+ $X2=8.365 $Y2=2.06
r235 43 44 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=8.28 $Y=2.06
+ $X2=6.985 $Y2=2.06
r236 42 63 3.85266 $w=1.7e-07 $l=1.60624e-07 $layer=LI1_cond $X=4.655 $Y=1.89
+ $X2=4.535 $Y2=1.985
r237 41 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.815 $Y=1.89
+ $X2=6.9 $Y2=1.89
r238 41 42 140.92 $w=1.68e-07 $l=2.16e-06 $layer=LI1_cond $X=6.815 $Y=1.89
+ $X2=4.655 $Y2=1.89
r239 39 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.535
+ $Y=2 $X2=4.535 $Y2=2
r240 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.535
+ $Y=1.66 $X2=4.535 $Y2=1.66
r241 36 63 3.22548 $w=2.4e-07 $l=1.8e-07 $layer=LI1_cond $X=4.535 $Y=1.805
+ $X2=4.535 $Y2=1.985
r242 36 38 6.96268 $w=2.38e-07 $l=1.45e-07 $layer=LI1_cond $X=4.535 $Y=1.805
+ $X2=4.535 $Y2=1.66
r243 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.75
+ $Y=3.59 $X2=2.75 $Y2=3.59
r244 31 33 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=2.75 $Y=2.445
+ $X2=2.75 $Y2=3.59
r245 30 61 3.22099 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.005 $Y=2.36
+ $X2=1.847 $Y2=2.36
r246 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.665 $Y=2.36
+ $X2=2.75 $Y2=2.445
r247 29 30 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.665 $Y=2.36
+ $X2=2.005 $Y2=2.36
r248 27 61 3.32435 $w=2.82e-07 $l=8.5e-08 $layer=LI1_cond $X=1.847 $Y=2.445
+ $X2=1.847 $Y2=2.36
r249 27 60 18.2927 $w=3.13e-07 $l=5e-07 $layer=LI1_cond $X=1.847 $Y=2.445
+ $X2=1.847 $Y2=2.945
r250 23 61 3.32435 $w=2.82e-07 $l=9.97246e-08 $layer=LI1_cond $X=1.815 $Y=2.275
+ $X2=1.847 $Y2=2.36
r251 23 25 64.9978 $w=2.48e-07 $l=1.41e-06 $layer=LI1_cond $X=1.815 $Y=2.275
+ $X2=1.815 $Y2=0.865
r252 21 60 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.84 $Y=3.11
+ $X2=1.84 $Y2=2.945
r253 18 34 89.8849 $w=5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.59 $Y=3.655
+ $X2=2.75 $Y2=3.655
r254 15 75 39.5806 $w=5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.685 $Y=1.315
+ $X2=8.685 $Y2=1.71
r255 15 17 24.582 $w=5e-07 $l=2.55e-07 $layer=POLY_cond $X=8.685 $Y=1.315
+ $X2=8.685 $Y2=1.06
r256 11 39 0.392508 $w=6.14e-07 $l=5e-09 $layer=POLY_cond $X=4.54 $Y=1.755
+ $X2=4.535 $Y2=1.755
r257 11 13 78.1143 $w=5e-07 $l=7.3e-07 $layer=POLY_cond $X=4.54 $Y=1.475
+ $X2=4.54 $Y2=0.745
r258 8 18 26.9307 $w=5e-07 $l=3.53553e-07 $layer=POLY_cond $X=3.84 $Y=3.405
+ $X2=3.59 $Y2=3.655
r259 8 10 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.84 $Y=3.405 $X2=3.84
+ $Y2=2.855
r260 7 39 54.5586 $w=6.14e-07 $l=1.07261e-06 $layer=POLY_cond $X=3.84 $Y=2.535
+ $X2=4.535 $Y2=1.755
r261 7 10 34.2419 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.84 $Y=2.535 $X2=3.84
+ $Y2=2.855
r262 2 21 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.7
+ $Y=2.965 $X2=1.84 $Y2=3.11
r263 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.715
+ $Y=0.655 $X2=1.855 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%A_1000_81# 1 2 9 13 14 17 20 24 27 28 29 31
+ 35 41
c73 28 0 1.48283e-19 $X=5.425 $Y=2.59
c74 13 0 6.88421e-21 $X=5.37 $Y=2.285
r75 35 38 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=6.73 $Y=2.76
+ $X2=6.73 $Y2=2.855
r76 31 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.2 $Y=2.59 $X2=6.2
+ $Y2=2.76
r77 30 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.285 $Y=2.76
+ $X2=6.2 $Y2=2.76
r78 29 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.565 $Y=2.76
+ $X2=6.73 $Y2=2.76
r79 29 30 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.565 $Y=2.76
+ $X2=6.285 $Y2=2.76
r80 27 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.115 $Y=2.59
+ $X2=6.2 $Y2=2.59
r81 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.115 $Y=2.59
+ $X2=5.425 $Y2=2.59
r82 25 41 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=5.37 $Y=3.39 $X2=5.37
+ $Y2=2.855
r83 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.305
+ $Y=3.39 $X2=5.305 $Y2=3.39
r84 22 28 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=5.305 $Y=2.675
+ $X2=5.425 $Y2=2.59
r85 22 24 34.3332 $w=2.38e-07 $l=7.15e-07 $layer=LI1_cond $X=5.305 $Y=2.675
+ $X2=5.305 $Y2=3.39
r86 17 45 23.0071 $w=5e-07 $l=1.85e-07 $layer=POLY_cond $X=5.25 $Y=1.47 $X2=5.25
+ $Y2=1.655
r87 16 20 14.8702 $w=3.08e-07 $l=4e-07 $layer=LI1_cond $X=5.3 $Y=1.47 $X2=5.7
+ $Y2=1.47
r88 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.3
+ $Y=1.47 $X2=5.3 $Y2=1.47
r89 14 45 55.6154 $w=3.8e-07 $l=3.8e-07 $layer=POLY_cond $X=5.31 $Y=2.035
+ $X2=5.31 $Y2=1.655
r90 13 41 60.9934 $w=5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.37 $Y=2.285 $X2=5.37
+ $Y2=2.855
r91 13 14 29.9625 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.37 $Y=2.285 $X2=5.37
+ $Y2=2.035
r92 7 17 6.95538 $w=5e-07 $l=6.5e-08 $layer=POLY_cond $X=5.25 $Y=1.405 $X2=5.25
+ $Y2=1.47
r93 7 9 70.6239 $w=5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.25 $Y=1.405 $X2=5.25
+ $Y2=0.745
r94 2 38 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.59
+ $Y=2.645 $X2=6.73 $Y2=2.855
r95 1 20 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=1.255 $X2=5.7 $Y2=1.465
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%SET_B 3 6 8 9 12 16 17 20 23 25 26 27 28 29
+ 30 31 40 41 44 46 49 61
c94 46 0 2.65827e-19 $X=7.182 $Y=1.545
c95 41 0 8.88678e-20 $X=11.05 $Y=0.72
c96 17 0 2.22527e-19 $X=7.93 $Y=1.675
r97 40 44 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=11.115 $Y=0.72
+ $X2=11.115 $Y2=1.225
r98 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.05
+ $Y=0.72 $X2=11.05 $Y2=0.72
r99 31 41 3.78945 $w=6.23e-07 $l=1.65e-07 $layer=LI1_cond $X=10.885 $Y=0.797
+ $X2=11.05 $Y2=0.797
r100 30 31 12.618 $w=4.53e-07 $l=4.8e-07 $layer=LI1_cond $X=10.32 $Y=0.782
+ $X2=10.8 $Y2=0.782
r101 29 30 12.618 $w=4.53e-07 $l=4.8e-07 $layer=LI1_cond $X=9.84 $Y=0.782
+ $X2=10.32 $Y2=0.782
r102 28 29 12.618 $w=4.53e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=0.782
+ $X2=9.84 $Y2=0.782
r103 27 28 12.618 $w=4.53e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=0.782
+ $X2=9.36 $Y2=0.782
r104 27 49 9.67378 $w=4.53e-07 $l=3.68e-07 $layer=LI1_cond $X=8.88 $Y=0.782
+ $X2=8.512 $Y2=0.782
r105 26 49 2.94419 $w=4.53e-07 $l=1.12e-07 $layer=LI1_cond $X=8.4 $Y=0.782
+ $X2=8.512 $Y2=0.782
r106 26 61 7.93754 $w=4.53e-07 $l=1.15e-07 $layer=LI1_cond $X=8.4 $Y=0.782
+ $X2=8.285 $Y2=0.782
r107 25 61 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.1 $Y=0.925
+ $X2=8.285 $Y2=0.925
r108 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.015 $Y=1.01
+ $X2=8.1 $Y2=0.925
r109 22 23 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=8.015 $Y=1.01
+ $X2=8.015 $Y2=1.555
r110 20 47 30.3683 $w=6.65e-07 $l=3.35e-07 $layer=POLY_cond $X=7.182 $Y=1.71
+ $X2=7.182 $Y2=2.045
r111 20 46 16.6909 $w=6.65e-07 $l=1.65e-07 $layer=POLY_cond $X=7.182 $Y=1.71
+ $X2=7.182 $Y2=1.545
r112 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.33
+ $Y=1.71 $X2=7.33 $Y2=1.71
r113 17 23 7.07814 $w=2.4e-07 $l=1.56844e-07 $layer=LI1_cond $X=7.93 $Y=1.675
+ $X2=8.015 $Y2=1.555
r114 17 19 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=7.93 $Y=1.675
+ $X2=7.33 $Y2=1.675
r115 15 44 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=11.115 $Y=1.565
+ $X2=11.115 $Y2=1.225
r116 12 16 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=11.185 $Y=2.785
+ $X2=11.185 $Y2=2.445
r117 9 16 27.696 $w=5.7e-07 $l=2.85e-07 $layer=POLY_cond $X=11.15 $Y=2.16
+ $X2=11.15 $Y2=2.445
r118 8 15 27.696 $w=5.7e-07 $l=2.85e-07 $layer=POLY_cond $X=11.15 $Y=1.85
+ $X2=11.15 $Y2=1.565
r119 8 9 29.0981 $w=5.7e-07 $l=3.1e-07 $layer=POLY_cond $X=11.15 $Y=1.85
+ $X2=11.15 $Y2=2.16
r120 6 47 86.6748 $w=5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.12 $Y=2.855 $X2=7.12
+ $Y2=2.045
r121 3 46 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.1 $Y=1.225 $X2=7.1
+ $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%A_798_107# 1 2 7 10 13 15 20 23 25 27 30 34
+ 36 38 42 45 46
c120 42 0 8.51819e-20 $X=6.15 $Y=0.43
c121 38 0 1.80645e-19 $X=5.985 $Y=1.05
c122 27 0 1.62708e-19 $X=7.995 $Y=2.465
c123 25 0 3.72258e-20 $X=6.215 $Y=2.515
r124 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.15
+ $Y=0.43 $X2=6.15 $Y2=0.43
r125 40 42 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=6.15 $Y=0.965
+ $X2=6.15 $Y2=0.43
r126 39 45 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.315 $Y=1.05
+ $X2=4.19 $Y2=1.05
r127 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.985 $Y=1.05
+ $X2=6.15 $Y2=0.965
r128 38 39 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=5.985 $Y=1.05
+ $X2=4.315 $Y2=1.05
r129 34 46 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.23 $Y=2.77
+ $X2=4.23 $Y2=2.605
r130 34 36 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.23 $Y=2.77
+ $X2=4.23 $Y2=2.855
r131 32 45 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.15 $Y=1.135
+ $X2=4.19 $Y2=1.05
r132 32 46 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=4.15 $Y=1.135
+ $X2=4.15 $Y2=2.605
r133 28 45 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.19 $Y=0.965
+ $X2=4.19 $Y2=1.05
r134 28 30 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=4.19 $Y=0.965
+ $X2=4.19 $Y2=0.745
r135 26 27 37.6502 $w=5.4e-07 $l=3.8e-07 $layer=POLY_cond $X=7.995 $Y=2.085
+ $X2=7.995 $Y2=2.465
r136 24 25 50.046 $w=7.5e-07 $l=7.3e-07 $layer=POLY_cond $X=6.215 $Y=1.785
+ $X2=6.215 $Y2=2.515
r137 23 27 58.804 $w=5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.015 $Y=3.075
+ $X2=8.015 $Y2=2.465
r138 20 26 109.681 $w=5e-07 $l=1.025e-06 $layer=POLY_cond $X=7.975 $Y=1.06
+ $X2=7.975 $Y2=2.085
r139 17 20 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.975 $Y=0.575
+ $X2=7.975 $Y2=1.06
r140 16 43 14.4767 $w=4.35e-07 $l=2.5e-07 $layer=POLY_cond $X=6.34 $Y=0.357
+ $X2=6.09 $Y2=0.357
r141 15 17 27.1004 $w=4.35e-07 $l=3.42053e-07 $layer=POLY_cond $X=7.725 $Y=0.357
+ $X2=7.975 $Y2=0.575
r142 15 16 177.074 $w=4.35e-07 $l=1.385e-06 $layer=POLY_cond $X=7.725 $Y=0.357
+ $X2=6.34 $Y2=0.357
r143 13 25 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.34 $Y=2.855 $X2=6.34
+ $Y2=2.515
r144 10 24 34.2419 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.09 $Y=1.465
+ $X2=6.09 $Y2=1.785
r145 7 43 12.6237 $w=5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.09 $Y=0.575
+ $X2=6.09 $Y2=0.357
r146 7 10 95.2352 $w=5e-07 $l=8.9e-07 $layer=POLY_cond $X=6.09 $Y=0.575 $X2=6.09
+ $Y2=1.465
r147 2 36 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.09
+ $Y=2.645 $X2=4.23 $Y2=2.855
r148 1 30 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.535 $X2=4.15 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%A_2031_177# 1 2 7 9 11 13 17 20 22 28 30 34
c74 30 0 6.97556e-20 $X=10.405 $Y=1.225
c75 13 0 1.25177e-19 $X=12.39 $Y=3.09
c76 9 0 1.57837e-19 $X=11.425 $Y=3.38
r77 23 34 115.031 $w=5e-07 $l=1.075e-06 $layer=POLY_cond $X=10.405 $Y=1.71
+ $X2=10.405 $Y2=2.785
r78 23 30 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=10.405 $Y=1.71
+ $X2=10.405 $Y2=1.225
r79 22 25 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=10.47 $Y=1.71
+ $X2=10.47 $Y2=1.74
r80 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.47
+ $Y=1.71 $X2=10.47 $Y2=1.71
r81 19 28 3.70735 $w=2.5e-07 $l=1.72337e-07 $layer=LI1_cond $X=12.475 $Y=1.825
+ $X2=12.34 $Y2=1.74
r82 19 20 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=12.475 $Y=1.825
+ $X2=12.475 $Y2=3.005
r83 15 28 3.70735 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=12.285 $Y=1.655
+ $X2=12.34 $Y2=1.74
r84 15 17 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.285 $Y=1.655
+ $X2=12.285 $Y2=1.225
r85 14 27 1.57051 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.55 $Y=3.09
+ $X2=11.425 $Y2=3.09
r86 13 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.39 $Y=3.09
+ $X2=12.475 $Y2=3.005
r87 13 14 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=12.39 $Y=3.09
+ $X2=11.55 $Y2=3.09
r88 9 27 14.7546 $w=2.5e-07 $l=2.9e-07 $layer=LI1_cond $X=11.425 $Y=3.38
+ $X2=11.425 $Y2=3.09
r89 9 11 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=11.425 $Y=3.38
+ $X2=11.425 $Y2=3.505
r90 8 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.635 $Y=1.74
+ $X2=10.47 $Y2=1.74
r91 7 28 2.76166 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=12.12 $Y=1.74
+ $X2=12.34 $Y2=1.74
r92 7 8 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=12.12 $Y=1.74
+ $X2=10.635 $Y2=1.74
r93 2 11 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=11.32
+ $Y=3.295 $X2=11.465 $Y2=3.505
r94 1 17 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.145
+ $Y=1.015 $X2=12.285 $Y2=1.225
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%A_1787_137# 1 2 3 12 16 19 23 25 27 28 29
+ 30 31 35 40 42 43 45 48 49
c125 35 0 6.97556e-20 $X=9.49 $Y=3.22
c126 29 0 1.57837e-19 $X=12.027 $Y=3.185
c127 19 0 1.25177e-19 $X=13.05 $Y=2.235
c128 12 0 8.88678e-20 $X=11.895 $Y=1.225
r129 49 51 7.28358 $w=5.36e-07 $l=4.21426e-07 $layer=LI1_cond $X=11.81 $Y=2.4
+ $X2=11.575 $Y2=2.72
r130 47 49 5.23507 $w=5.36e-07 $l=3.30568e-07 $layer=LI1_cond $X=12.045 $Y=2.17
+ $X2=11.81 $Y2=2.4
r131 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.045
+ $Y=2.17 $X2=12.045 $Y2=2.17
r132 44 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=2.4
+ $X2=9.575 $Y2=2.4
r133 43 49 7.59541 $w=1.7e-07 $l=4e-07 $layer=LI1_cond $X=11.41 $Y=2.4 $X2=11.81
+ $Y2=2.4
r134 43 44 114.171 $w=1.68e-07 $l=1.75e-06 $layer=LI1_cond $X=11.41 $Y=2.4
+ $X2=9.66 $Y2=2.4
r135 41 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.575 $Y=2.485
+ $X2=9.575 $Y2=2.4
r136 41 42 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=9.575 $Y=2.485
+ $X2=9.575 $Y2=3.025
r137 40 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.575 $Y=2.315
+ $X2=9.575 $Y2=2.4
r138 39 40 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=9.575 $Y=1.475
+ $X2=9.575 $Y2=2.315
r139 35 42 8.28377 $w=3.9e-07 $l=2.33666e-07 $layer=LI1_cond $X=9.49 $Y=3.22
+ $X2=9.575 $Y2=3.025
r140 35 37 8.27395 $w=3.88e-07 $l=2.8e-07 $layer=LI1_cond $X=9.49 $Y=3.22
+ $X2=9.21 $Y2=3.22
r141 31 39 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=9.49 $Y=1.332
+ $X2=9.575 $Y2=1.475
r142 31 33 12.131 $w=2.83e-07 $l=3e-07 $layer=LI1_cond $X=9.49 $Y=1.332 $X2=9.19
+ $Y2=1.332
r143 28 29 22.5012 $w=5.35e-07 $l=2.25e-07 $layer=POLY_cond $X=12.027 $Y=2.96
+ $X2=12.027 $Y2=3.185
r144 25 30 20.4101 $w=5e-07 $l=2.59808e-07 $layer=POLY_cond $X=13.34 $Y=2.485
+ $X2=13.32 $Y2=2.235
r145 25 27 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=13.34 $Y=2.485
+ $X2=13.34 $Y2=2.97
r146 21 30 20.4101 $w=5e-07 $l=2.59808e-07 $layer=POLY_cond $X=13.3 $Y=1.985
+ $X2=13.32 $Y2=2.235
r147 21 23 81.3245 $w=5e-07 $l=7.6e-07 $layer=POLY_cond $X=13.3 $Y=1.985
+ $X2=13.3 $Y2=1.225
r148 20 48 5.30422 $w=5e-07 $l=3.25e-07 $layer=POLY_cond $X=12.295 $Y=2.235
+ $X2=11.97 $Y2=2.235
r149 19 30 5.30422 $w=5e-07 $l=2.7e-07 $layer=POLY_cond $X=13.05 $Y=2.235
+ $X2=13.32 $Y2=2.235
r150 19 20 80.7895 $w=5e-07 $l=7.55e-07 $layer=POLY_cond $X=13.05 $Y=2.235
+ $X2=12.295 $Y2=2.235
r151 17 48 20.4101 $w=5e-07 $l=2.85044e-07 $layer=POLY_cond $X=12.045 $Y=2.485
+ $X2=11.97 $Y2=2.235
r152 17 28 50.8278 $w=5e-07 $l=4.75e-07 $layer=POLY_cond $X=12.045 $Y=2.485
+ $X2=12.045 $Y2=2.96
r153 16 29 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=12.01 $Y=3.505
+ $X2=12.01 $Y2=3.185
r154 10 48 20.4101 $w=5e-07 $l=2.85044e-07 $layer=POLY_cond $X=11.895 $Y=1.985
+ $X2=11.97 $Y2=2.235
r155 10 12 81.3245 $w=5e-07 $l=7.6e-07 $layer=POLY_cond $X=11.895 $Y=1.985
+ $X2=11.895 $Y2=1.225
r156 3 51 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.435
+ $Y=2.575 $X2=11.575 $Y2=2.72
r157 2 37 600 $w=1.7e-07 $l=7.53392e-07 $layer=licon1_PDIFF $count=1 $X=8.975
+ $Y=2.575 $X2=9.21 $Y2=3.22
r158 1 33 182 $w=1.7e-07 $l=7.21318e-07 $layer=licon1_NDIFF $count=1 $X=8.935
+ $Y=0.685 $X2=9.19 $Y2=1.29
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%A_2553_203# 1 2 9 13 15 18 21 24 27 29 33
+ 34 36 37
r63 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.075
+ $Y=1.89 $X2=14.075 $Y2=1.89
r64 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=14.075 $Y=2.225
+ $X2=14.075 $Y2=1.89
r65 30 37 2.45049 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.115 $Y=2.31
+ $X2=12.99 $Y2=2.31
r66 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.91 $Y=2.31
+ $X2=14.075 $Y2=2.225
r67 29 30 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=13.91 $Y=2.31
+ $X2=13.115 $Y2=2.31
r68 25 37 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.99 $Y=2.395
+ $X2=12.99 $Y2=2.31
r69 25 27 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=12.99 $Y=2.395
+ $X2=12.99 $Y2=2.74
r70 24 37 3.98977 $w=2.3e-07 $l=9.44722e-08 $layer=LI1_cond $X=12.97 $Y=2.225
+ $X2=12.99 $Y2=2.31
r71 24 36 39.6104 $w=2.08e-07 $l=7.5e-07 $layer=LI1_cond $X=12.97 $Y=2.225
+ $X2=12.97 $Y2=1.475
r72 19 36 7.28026 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.91 $Y=1.31
+ $X2=12.91 $Y2=1.475
r73 19 21 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=12.91 $Y=1.31
+ $X2=12.91 $Y2=1.225
r74 17 34 26.798 $w=5.75e-07 $l=2.88e-07 $layer=POLY_cond $X=14.177 $Y=2.178
+ $X2=14.177 $Y2=1.89
r75 17 18 27.7583 $w=5.75e-07 $l=2.87e-07 $layer=POLY_cond $X=14.177 $Y=2.178
+ $X2=14.177 $Y2=2.465
r76 15 34 3.53585 $w=5.75e-07 $l=3.8e-08 $layer=POLY_cond $X=14.177 $Y=1.852
+ $X2=14.177 $Y2=1.89
r77 15 16 27.4041 $w=5.75e-07 $l=2.87e-07 $layer=POLY_cond $X=14.177 $Y=1.852
+ $X2=14.177 $Y2=1.565
r78 13 18 67.4137 $w=5e-07 $l=6.3e-07 $layer=POLY_cond $X=14.215 $Y=3.095
+ $X2=14.215 $Y2=2.465
r79 9 16 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=14.195 $Y=1.06
+ $X2=14.195 $Y2=1.565
r80 2 27 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=12.825
+ $Y=2.595 $X2=12.95 $Y2=2.74
r81 1 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=12.765
+ $Y=1.015 $X2=12.91 $Y2=1.225
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%VPWR 1 2 3 4 5 6 7 22 25 34 41 48 59 72 77
+ 85
r121 83 85 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=13.405 $Y=3.63
+ $X2=14.125 $Y2=3.63
r122 82 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.125 $Y=3.59
+ $X2=14.125 $Y2=3.59
r123 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.405 $Y=3.59
+ $X2=13.405 $Y2=3.59
r124 80 82 1.80741 $w=9.43e-07 $l=1.4e-07 $layer=LI1_cond $X=13.767 $Y=3.45
+ $X2=13.767 $Y2=3.59
r125 77 80 9.16614 $w=9.43e-07 $l=7.1e-07 $layer=LI1_cond $X=13.767 $Y=2.74
+ $X2=13.767 $Y2=3.45
r126 74 83 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=12.565 $Y=3.63
+ $X2=13.405 $Y2=3.63
r127 72 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.565 $Y=3.59
+ $X2=12.565 $Y2=3.59
r128 69 74 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=11.845 $Y=3.63
+ $X2=12.565 $Y2=3.63
r129 68 72 16.8317 $w=3.78e-07 $l=5.55e-07 $layer=LI1_cond $X=11.845 $Y=3.545
+ $X2=12.4 $Y2=3.545
r130 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.845 $Y=3.59
+ $X2=11.845 $Y2=3.59
r131 65 69 0.383905 $w=3.7e-07 $l=1e-06 $layer=MET1_cond $X=10.845 $Y=3.63
+ $X2=11.845 $Y2=3.63
r132 63 65 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.125 $Y=3.63
+ $X2=10.845 $Y2=3.63
r133 62 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.845 $Y=3.59
+ $X2=10.845 $Y2=3.59
r134 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.125 $Y=3.59
+ $X2=10.125 $Y2=3.59
r135 59 62 10.0168 $w=9.48e-07 $l=7.8e-07 $layer=LI1_cond $X=10.485 $Y=2.81
+ $X2=10.485 $Y2=3.59
r136 56 63 0.85035 $w=3.7e-07 $l=2.215e-06 $layer=MET1_cond $X=7.91 $Y=3.63
+ $X2=10.125 $Y2=3.63
r137 53 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.91 $Y=3.59
+ $X2=7.91 $Y2=3.59
r138 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.19 $Y=3.59
+ $X2=7.19 $Y2=3.59
r139 51 53 6.22842 $w=9.48e-07 $l=4.85e-07 $layer=LI1_cond $X=7.55 $Y=3.105
+ $X2=7.55 $Y2=3.59
r140 48 51 4.43053 $w=9.48e-07 $l=3.45e-07 $layer=LI1_cond $X=7.55 $Y=2.76
+ $X2=7.55 $Y2=3.105
r141 45 54 0.564341 $w=3.7e-07 $l=1.47e-06 $layer=MET1_cond $X=5.72 $Y=3.63
+ $X2=7.19 $Y2=3.63
r142 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.72 $Y=3.59
+ $X2=5.72 $Y2=3.59
r143 41 44 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=5.77 $Y=2.94
+ $X2=5.77 $Y2=3.59
r144 38 45 1.29376 $w=3.7e-07 $l=3.37e-06 $layer=MET1_cond $X=2.35 $Y=3.63
+ $X2=5.72 $Y2=3.63
r145 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.35 $Y=3.59
+ $X2=2.35 $Y2=3.59
r146 34 37 33.8818 $w=2.48e-07 $l=7.35e-07 $layer=LI1_cond $X=2.36 $Y=2.855
+ $X2=2.36 $Y2=3.59
r147 31 38 0.372388 $w=3.7e-07 $l=9.7e-07 $layer=MET1_cond $X=1.38 $Y=3.63
+ $X2=2.35 $Y2=3.63
r148 29 31 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.66 $Y=3.63
+ $X2=1.38 $Y2=3.63
r149 28 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.38 $Y=3.59
+ $X2=1.38 $Y2=3.59
r150 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.66 $Y=3.59
+ $X2=0.66 $Y2=3.59
r151 25 28 6.42105 $w=9.48e-07 $l=5e-07 $layer=LI1_cond $X=1.02 $Y=3.09 $X2=1.02
+ $Y2=3.59
r152 22 56 0.180436 $w=3.7e-07 $l=4.7e-07 $layer=MET1_cond $X=7.44 $Y=3.63
+ $X2=7.91 $Y2=3.63
r153 22 54 0.0959764 $w=3.7e-07 $l=2.5e-07 $layer=MET1_cond $X=7.44 $Y=3.63
+ $X2=7.19 $Y2=3.63
r154 7 80 600 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=13.59
+ $Y=2.595 $X2=13.825 $Y2=3.45
r155 7 77 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=13.59
+ $Y=2.595 $X2=13.825 $Y2=2.74
r156 6 72 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=12.26
+ $Y=3.295 $X2=12.4 $Y2=3.505
r157 5 59 600 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=10.655
+ $Y=2.575 $X2=10.795 $Y2=2.81
r158 4 51 300 $w=1.7e-07 $l=5.73498e-07 $layer=licon1_PDIFF $count=2 $X=7.37
+ $Y=2.645 $X2=7.625 $Y2=3.105
r159 4 48 600 $w=1.7e-07 $l=3.07164e-07 $layer=licon1_PDIFF $count=1 $X=7.37
+ $Y=2.645 $X2=7.625 $Y2=2.76
r160 3 41 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=5.62
+ $Y=2.645 $X2=5.77 $Y2=2.94
r161 2 34 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=2.645 $X2=2.4 $Y2=2.855
r162 1 25 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.92
+ $Y=2.965 $X2=1.06 $Y2=3.09
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%A_642_107# 1 2 9 12
r20 12 14 11.2873 $w=3.48e-07 $l=2.5e-07 $layer=LI1_cond $X=3.36 $Y=0.745
+ $X2=3.36 $Y2=0.995
r21 9 14 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=3.45 $Y=2.855
+ $X2=3.45 $Y2=0.995
r22 2 9 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.31
+ $Y=2.645 $X2=3.45 $Y2=2.855
r23 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.21
+ $Y=0.535 $X2=3.35 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%Q 1 2 7 8 9 10 11 12 13 22
r15 13 40 10.0427 $w=3.48e-07 $l=3.05e-07 $layer=LI1_cond $X=14.595 $Y=3.145
+ $X2=14.595 $Y2=3.45
r16 12 13 13.3354 $w=3.48e-07 $l=4.05e-07 $layer=LI1_cond $X=14.595 $Y=2.74
+ $X2=14.595 $Y2=3.145
r17 11 12 11.0305 $w=3.48e-07 $l=3.35e-07 $layer=LI1_cond $X=14.595 $Y=2.405
+ $X2=14.595 $Y2=2.74
r18 10 11 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=14.595 $Y=2.035
+ $X2=14.595 $Y2=2.405
r19 9 10 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=14.595 $Y=1.665
+ $X2=14.595 $Y2=2.035
r20 8 9 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=14.595 $Y=1.295
+ $X2=14.595 $Y2=1.665
r21 7 8 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=14.595 $Y=0.925
+ $X2=14.595 $Y2=1.295
r22 7 22 3.7866 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=14.595 $Y=0.925
+ $X2=14.595 $Y2=0.81
r23 2 40 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=14.465
+ $Y=2.595 $X2=14.605 $Y2=3.45
r24 2 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=14.465
+ $Y=2.595 $X2=14.605 $Y2=2.74
r25 1 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=14.445
+ $Y=0.685 $X2=14.585 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HVL__DFSTP_1%VGND 1 2 3 4 5 6 19 22 29 42 46 57 64 68
r100 70 72 6.42105 $w=9.48e-07 $l=5e-07 $layer=LI1_cond $X=13.73 $Y=0.81
+ $X2=13.73 $Y2=1.31
r101 65 68 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=13.37 $Y=0.44
+ $X2=14.09 $Y2=0.44
r102 64 70 4.23789 $w=9.48e-07 $l=3.3e-07 $layer=LI1_cond $X=13.73 $Y=0.48
+ $X2=13.73 $Y2=0.81
r103 64 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.09 $Y=0.48
+ $X2=14.09 $Y2=0.48
r104 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.37 $Y=0.48
+ $X2=13.37 $Y2=0.48
r105 58 65 0.596973 $w=3.7e-07 $l=1.555e-06 $layer=MET1_cond $X=11.815 $Y=0.44
+ $X2=13.37 $Y2=0.44
r106 57 61 15.103 $w=5.88e-07 $l=7.45e-07 $layer=LI1_cond $X=11.635 $Y=0.48
+ $X2=11.635 $Y2=1.225
r107 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.815 $Y=0.48
+ $X2=11.815 $Y2=0.48
r108 52 54 5.90737 $w=9.48e-07 $l=4.6e-07 $layer=LI1_cond $X=7.275 $Y=0.83
+ $X2=7.275 $Y2=1.29
r109 50 58 1.60472 $w=3.7e-07 $l=4.18e-06 $layer=MET1_cond $X=7.635 $Y=0.44
+ $X2=11.815 $Y2=0.44
r110 46 52 4.49474 $w=9.48e-07 $l=3.5e-07 $layer=LI1_cond $X=7.275 $Y=0.48
+ $X2=7.275 $Y2=0.83
r111 46 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.635 $Y=0.48
+ $X2=7.635 $Y2=0.48
r112 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.915 $Y=0.48
+ $X2=6.915 $Y2=0.48
r113 43 47 0.470284 $w=3.7e-07 $l=1.225e-06 $layer=MET1_cond $X=5.69 $Y=0.44
+ $X2=6.915 $Y2=0.44
r114 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.69 $Y=0.48
+ $X2=5.69 $Y2=0.48
r115 40 42 1.37196 $w=4.18e-07 $l=5e-08 $layer=LI1_cond $X=5.64 $Y=0.575
+ $X2=5.69 $Y2=0.575
r116 37 43 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=4.97 $Y=0.44
+ $X2=5.69 $Y2=0.44
r117 36 40 18.3842 $w=4.18e-07 $l=6.7e-07 $layer=LI1_cond $X=4.97 $Y=0.575
+ $X2=5.64 $Y2=0.575
r118 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.97 $Y=0.48
+ $X2=4.97 $Y2=0.48
r119 30 37 0.788926 $w=3.7e-07 $l=2.055e-06 $layer=MET1_cond $X=2.915 $Y=0.44
+ $X2=4.97 $Y2=0.44
r120 29 33 5.9245 $w=5.33e-07 $l=2.65e-07 $layer=LI1_cond $X=2.737 $Y=0.48
+ $X2=2.737 $Y2=0.745
r121 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.915 $Y=0.48
+ $X2=2.915 $Y2=0.48
r122 23 30 0.717903 $w=3.7e-07 $l=1.87e-06 $layer=MET1_cond $X=1.045 $Y=0.44
+ $X2=2.915 $Y2=0.44
r123 22 26 7.80492 $w=5.88e-07 $l=3.85e-07 $layer=LI1_cond $X=0.865 $Y=0.48
+ $X2=0.865 $Y2=0.865
r124 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.045 $Y=0.48
+ $X2=1.045 $Y2=0.48
r125 19 50 0.0748616 $w=3.7e-07 $l=1.95e-07 $layer=MET1_cond $X=7.44 $Y=0.44
+ $X2=7.635 $Y2=0.44
r126 19 47 0.20155 $w=3.7e-07 $l=5.25e-07 $layer=MET1_cond $X=7.44 $Y=0.44
+ $X2=6.915 $Y2=0.44
r127 6 72 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=13.55
+ $Y=1.015 $X2=13.805 $Y2=1.31
r128 6 70 182 $w=1.7e-07 $l=3.42491e-07 $layer=licon1_NDIFF $count=1 $X=13.55
+ $Y=1.015 $X2=13.805 $Y2=0.81
r129 5 61 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.365
+ $Y=1.015 $X2=11.505 $Y2=1.225
r130 4 54 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=7.35
+ $Y=1.015 $X2=7.585 $Y2=1.29
r131 4 52 182 $w=1.7e-07 $l=3.14166e-07 $layer=licon1_NDIFF $count=1 $X=7.35
+ $Y=1.015 $X2=7.585 $Y2=0.83
r132 3 40 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=5.5
+ $Y=0.535 $X2=5.64 $Y2=0.69
r133 2 33 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.535 $X2=2.57 $Y2=0.745
r134 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.935
+ $Y=0.655 $X2=1.075 $Y2=0.865
.ends

