* NGSPICE file created from sky130_fd_sc_hvl__fill_4.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__fill_4 VGND VNB VPB VPWR
.ends

