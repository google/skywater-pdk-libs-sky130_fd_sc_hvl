# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hvl__dfsbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  17.76000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.515000 2.875000 2.145000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.498750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.300000 0.495000 17.635000 1.325000 ;
        RECT 17.300000 2.355000 17.635000 3.435000 ;
        RECT 17.405000 1.325000 17.635000 2.355000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.015000 0.495000 15.375000 3.755000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  6.985000 1.155000 10.330000 1.325000 ;
        RECT 10.160000 1.325000 10.330000 1.605000 ;
        RECT 10.160000 1.605000 10.885000 1.775000 ;
        RECT 10.715000 1.775000 10.885000 1.975000 ;
        RECT 10.715000 1.975000 12.830000 2.145000 ;
        RECT 12.150000 1.555000 12.830000 1.975000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.550000 0.890000 2.520000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.365000 1.490000 1.020000 ;
    END
    PORT
      LAYER li1 ;
        RECT 12.200000 0.365000 13.150000 0.975000 ;
    END
    PORT
      LAYER li1 ;
        RECT 13.900000 0.365000 14.835000 1.025000 ;
    END
    PORT
      LAYER li1 ;
        RECT 16.155000 0.365000 17.105000 1.305000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.220000 0.365000 2.470000 0.985000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.650000 0.365000 5.600000 0.905000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.785000 0.365000 7.735000 0.975000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 17.760000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 17.760000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 17.760000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 17.760000 4.155000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 17.760000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.650000 2.700000 1.240000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 10.715000 2.675000 11.665000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 13.870000 2.255000 14.820000 3.755000 ;
    END
    PORT
      LAYER li1 ;
        RECT 16.135000 2.355000 17.085000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.470000 2.675000 2.675000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.680000 2.905000 6.245000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.855000 2.895000 8.805000 3.705000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 17.760000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.110000 0.540000  0.360000 1.200000 ;
      RECT  0.110000 1.200000  1.590000 1.370000 ;
      RECT  0.110000 1.370000  0.380000 3.450000 ;
      RECT  1.260000 1.370000  1.590000 1.870000 ;
      RECT  1.420000 1.870000  1.590000 3.630000 ;
      RECT  1.420000 3.630000  2.290000 3.800000 ;
      RECT  1.670000 0.540000  2.000000 1.000000 ;
      RECT  1.770000 1.000000  2.000000 1.165000 ;
      RECT  1.770000 1.165000  2.820000 1.335000 ;
      RECT  1.770000 1.335000  1.940000 3.450000 ;
      RECT  2.120000 2.325000  3.025000 2.495000 ;
      RECT  2.120000 2.495000  2.290000 3.630000 ;
      RECT  2.650000 0.265000  4.460000 0.435000 ;
      RECT  2.650000 0.435000  2.820000 1.165000 ;
      RECT  2.855000 2.495000  3.025000 3.355000 ;
      RECT  2.855000 3.355000  5.500000 3.525000 ;
      RECT  3.000000 0.615000  3.375000 1.005000 ;
      RECT  3.205000 1.005000  3.375000 2.675000 ;
      RECT  3.205000 2.675000  3.545000 3.175000 ;
      RECT  3.555000 1.105000  3.725000 2.225000 ;
      RECT  3.555000 2.225000  4.800000 2.395000 ;
      RECT  3.725000 2.395000  3.895000 3.355000 ;
      RECT  3.780000 0.615000  4.110000 0.925000 ;
      RECT  3.905000 0.925000  4.075000 1.855000 ;
      RECT  3.905000 1.855000  8.060000 2.025000 ;
      RECT  4.075000 2.675000  4.405000 3.005000 ;
      RECT  4.075000 3.005000  5.150000 3.175000 ;
      RECT  4.255000 1.105000  4.585000 1.505000 ;
      RECT  4.255000 1.505000  9.470000 1.675000 ;
      RECT  4.290000 0.435000  4.460000 1.105000 ;
      RECT  4.585000 2.395000  4.800000 2.555000 ;
      RECT  4.945000 1.085000  6.150000 1.325000 ;
      RECT  4.980000 2.025000  5.150000 3.005000 ;
      RECT  5.330000 2.205000  7.025000 2.375000 ;
      RECT  5.330000 2.555000  6.595000 2.725000 ;
      RECT  5.330000 2.725000  5.500000 3.355000 ;
      RECT  5.820000 0.515000  6.150000 1.085000 ;
      RECT  6.425000 2.725000  6.595000 3.355000 ;
      RECT  6.425000 3.355000  7.675000 3.525000 ;
      RECT  6.775000 2.375000  7.025000 3.175000 ;
      RECT  7.505000 2.545000  9.120000 2.715000 ;
      RECT  7.505000 2.715000  7.675000 3.355000 ;
      RECT  7.730000 2.025000  8.060000 2.365000 ;
      RECT  8.185000 0.375000 11.110000 0.545000 ;
      RECT  8.185000 0.545000  8.515000 0.975000 ;
      RECT  8.755000 0.725000 10.680000 0.975000 ;
      RECT  8.870000 1.885000  9.120000 2.545000 ;
      RECT  9.300000 1.675000  9.470000 2.305000 ;
      RECT  9.300000 2.305000 10.185000 2.475000 ;
      RECT  9.345000 2.675000  9.675000 3.585000 ;
      RECT  9.345000 3.585000 10.535000 3.755000 ;
      RECT  9.650000 1.505000  9.980000 1.955000 ;
      RECT  9.650000 1.955000 10.535000 2.125000 ;
      RECT  9.855000 2.475000 10.185000 2.555000 ;
      RECT 10.365000 2.125000 10.535000 2.325000 ;
      RECT 10.365000 2.325000 13.180000 2.495000 ;
      RECT 10.365000 2.495000 10.535000 3.585000 ;
      RECT 10.510000 0.975000 10.680000 1.255000 ;
      RECT 10.510000 1.255000 11.460000 1.425000 ;
      RECT 10.860000 0.545000 11.110000 1.075000 ;
      RECT 11.290000 0.515000 11.660000 0.975000 ;
      RECT 11.290000 0.975000 11.460000 1.255000 ;
      RECT 11.640000 1.155000 11.970000 1.205000 ;
      RECT 11.640000 1.205000 14.395000 1.375000 ;
      RECT 11.640000 1.375000 11.970000 1.795000 ;
      RECT 12.035000 2.495000 13.180000 3.175000 ;
      RECT 13.010000 1.555000 14.045000 1.725000 ;
      RECT 13.010000 1.725000 13.180000 2.325000 ;
      RECT 13.360000 1.905000 14.395000 2.075000 ;
      RECT 13.360000 2.075000 13.690000 2.675000 ;
      RECT 13.390000 0.825000 13.720000 1.205000 ;
      RECT 14.225000 1.375000 14.395000 1.905000 ;
      RECT 15.625000 0.825000 15.975000 1.505000 ;
      RECT 15.625000 1.505000 17.175000 1.675000 ;
      RECT 15.625000 1.675000 15.955000 3.185000 ;
      RECT 16.845000 1.675000 17.175000 2.175000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.570000  0.395000  0.740000 0.565000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.680000  3.505000  0.850000 3.675000 ;
      RECT  0.930000  0.395000  1.100000 0.565000 ;
      RECT  1.040000  3.505000  1.210000 3.675000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.290000  0.395000  1.460000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.250000  0.395000  2.420000 0.565000 ;
      RECT  2.490000  3.505000  2.660000 3.675000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.680000  0.395000  4.850000 0.565000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.040000  0.395000  5.210000 0.565000 ;
      RECT  5.400000  0.395000  5.570000 0.565000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.695000  3.505000  5.865000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.055000  3.505000  6.225000 3.675000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.815000  0.395000  6.985000 0.565000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.175000  0.395000  7.345000 0.565000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.535000  0.395000  7.705000 0.565000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  7.885000  3.505000  8.055000 3.675000 ;
      RECT  8.245000  3.505000  8.415000 3.675000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.605000  3.505000  8.775000 3.675000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.745000  3.505000 10.915000 3.675000 ;
      RECT 11.105000  3.505000 11.275000 3.675000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.465000  3.505000 11.635000 3.675000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.230000  0.395000 12.400000 0.565000 ;
      RECT 12.590000  0.395000 12.760000 0.565000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 12.950000  0.395000 13.120000 0.565000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.900000  3.505000 14.070000 3.675000 ;
      RECT 13.920000  0.395000 14.090000 0.565000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.260000  3.505000 14.430000 3.675000 ;
      RECT 14.280000  0.395000 14.450000 0.565000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.620000  3.505000 14.790000 3.675000 ;
      RECT 14.640000  0.395000 14.810000 0.565000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.165000  3.505000 16.335000 3.675000 ;
      RECT 16.185000  0.395000 16.355000 0.565000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.525000  3.505000 16.695000 3.675000 ;
      RECT 16.545000  0.395000 16.715000 0.565000 ;
      RECT 16.885000  3.505000 17.055000 3.675000 ;
      RECT 16.905000  0.395000 17.075000 0.565000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
  END
END sky130_fd_sc_hvl__dfsbp_1
END LIBRARY
