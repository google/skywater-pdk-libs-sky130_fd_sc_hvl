# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__nand3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__nand3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.455000 0.810000 2.725000 1.725000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 0.810000 2.275000 1.725000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.505000 0.995000 1.835000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.065000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.200000 1.905000 3.235000 2.075000 ;
        RECT 1.200000 2.075000 1.370000 3.755000 ;
        RECT 2.905000 0.495000 3.235000 1.325000 ;
        RECT 2.980000 1.325000 3.235000 1.905000 ;
        RECT 2.980000 2.075000 3.235000 3.755000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.360000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.360000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.985000 3.360000 4.155000 ;
      RECT 0.090000  0.365000 1.705000 1.325000 ;
      RECT 0.090000  2.175000 1.020000 3.755000 ;
      RECT 1.550000  2.255000 2.800000 3.755000 ;
    LAYER mcon ;
      RECT 0.095000  0.395000 0.265000 0.565000 ;
      RECT 0.110000  3.505000 0.280000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.455000  0.395000 0.625000 0.565000 ;
      RECT 0.470000  3.505000 0.640000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.815000  0.395000 0.985000 0.565000 ;
      RECT 0.830000  3.505000 1.000000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.175000  0.395000 1.345000 0.565000 ;
      RECT 1.535000  0.395000 1.705000 0.565000 ;
      RECT 1.550000  3.505000 1.720000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.910000  3.505000 2.080000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.270000  3.505000 2.440000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.630000  3.505000 2.800000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
  END
END sky130_fd_sc_hvl__nand3_1
END LIBRARY
