* File: sky130_fd_sc_hvl__conb_1.pxi.spice
* Created: Wed Sep  2 09:04:34 2020
* 
x_PM_SKY130_FD_SC_HVL__CONB_1%VNB N_VNB_X0_noxref_D0 VNB N_VNB_c_3_p VNB
+ PM_SKY130_FD_SC_HVL__CONB_1%VNB
x_PM_SKY130_FD_SC_HVL__CONB_1%VPB N_VPB_X0_noxref_D1 VPB N_VPB_c_22_p VPB
+ PM_SKY130_FD_SC_HVL__CONB_1%VPB
x_PM_SKY130_FD_SC_HVL__CONB_1%HI N_HI_R0_pos N_HI_c_49_p N_HI_c_41_n HI HI HI HI
+ N_HI_c_43_n PM_SKY130_FD_SC_HVL__CONB_1%HI
x_PM_SKY130_FD_SC_HVL__CONB_1%VPWR N_VPWR_R0_neg N_VPWR_c_77_n VPWR
+ N_VPWR_c_82_n N_VPWR_c_85_n PM_SKY130_FD_SC_HVL__CONB_1%VPWR
x_PM_SKY130_FD_SC_HVL__CONB_1%VGND N_VGND_R1_pos VGND N_VGND_c_103_n
+ N_VGND_c_105_n N_VGND_c_106_n N_VGND_c_108_n PM_SKY130_FD_SC_HVL__CONB_1%VGND
x_PM_SKY130_FD_SC_HVL__CONB_1%LO N_LO_R1_neg N_LO_c_127_n N_LO_c_132_n
+ N_LO_c_135_n LO LO LO LO LO PM_SKY130_FD_SC_HVL__CONB_1%LO
cc_1 N_VNB_X0_noxref_D0 N_HI_R0_pos 0.0883427f $X=-0.33 $Y=-0.265 $X2=0.84
+ $Y2=1.82
cc_2 N_VNB_X0_noxref_D0 N_HI_c_41_n 0.0293472f $X=-0.33 $Y=-0.265 $X2=0.455
+ $Y2=0.565
cc_3 N_VNB_c_3_p N_HI_c_41_n 0.00264305f $X=0.24 $Y=0 $X2=0.455 $Y2=0.565
cc_4 N_VNB_X0_noxref_D0 N_HI_c_43_n 0.14553f $X=-0.33 $Y=-0.265 $X2=0.84
+ $Y2=0.735
cc_5 N_VNB_c_3_p N_HI_c_43_n 0.00376473f $X=0.24 $Y=0 $X2=0.84 $Y2=0.735
cc_6 N_VNB_X0_noxref_D0 N_VPWR_c_77_n 0.00236338f $X=-0.33 $Y=-0.265 $X2=0.84
+ $Y2=1.82
cc_7 N_VNB_X0_noxref_D0 N_VGND_R1_pos 0.0883596f $X=-0.33 $Y=-0.265 $X2=0.84
+ $Y2=1.82
cc_8 N_VNB_X0_noxref_D0 N_VGND_c_103_n 0.123365f $X=-0.33 $Y=-0.265 $X2=1.115
+ $Y2=1.95
cc_9 N_VNB_c_3_p N_VGND_c_103_n 0.0010769f $X=0.24 $Y=0 $X2=1.115 $Y2=1.95
cc_10 N_VNB_X0_noxref_D0 N_VGND_c_105_n 0.0312779f $X=-0.33 $Y=-0.265 $X2=1.115
+ $Y2=2.32
cc_11 N_VNB_X0_noxref_D0 N_VGND_c_106_n 0.0473041f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_c_3_p N_VGND_c_106_n 0.00210617f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_13 N_VNB_X0_noxref_D0 N_VGND_c_108_n 0.0766646f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_c_3_p N_VGND_c_108_n 0.25664f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_15 N_VNB_X0_noxref_D0 N_LO_c_127_n 0.0023634f $X=-0.33 $Y=-0.265 $X2=0.84
+ $Y2=1.82
cc_16 N_VNB_X0_noxref_D0 LO 0.0106843f $X=-0.33 $Y=-0.265 $X2=0.577 $Y2=1.07
cc_17 N_VNB_c_3_p LO 0.00101616f $X=0.24 $Y=0 $X2=0.577 $Y2=1.07
cc_18 N_VNB_X0_noxref_D0 LO 0.00254362f $X=-0.33 $Y=-0.265 $X2=1.115 $Y2=2.69
cc_19 N_VPB_X0_noxref_D1 HI 0.00254166f $X=-0.33 $Y=1.885 $X2=1.115 $Y2=1.95
cc_20 N_VPB_X0_noxref_D1 HI 0.0021711f $X=-0.33 $Y=1.885 $X2=1.115 $Y2=2.32
cc_21 VPB HI 6.27922e-19 $X=0 $Y=3.955 $X2=1.115 $Y2=2.32
cc_22 N_VPB_c_22_p HI 0.00594087f $X=2.16 $Y=4.07 $X2=1.115 $Y2=2.32
cc_23 N_VPB_X0_noxref_D1 N_VPWR_c_77_n 0.151979f $X=-0.33 $Y=1.885 $X2=0.84
+ $Y2=1.82
cc_24 N_VPB_X0_noxref_D1 VPWR 0.0553552f $X=-0.33 $Y=1.885 $X2=0.74 $Y2=1.07
cc_25 VPB VPWR 0.251383f $X=0 $Y=3.955 $X2=0.74 $Y2=1.07
cc_26 N_VPB_c_22_p VPWR 0.0106344f $X=2.16 $Y=4.07 $X2=0.74 $Y2=1.07
cc_27 N_VPB_X0_noxref_D1 N_VPWR_c_82_n 0.0298923f $X=-0.33 $Y=1.885 $X2=0.455
+ $Y2=0.565
cc_28 VPB N_VPWR_c_82_n 0.00293269f $X=0 $Y=3.955 $X2=0.455 $Y2=0.565
cc_29 N_VPB_c_22_p N_VPWR_c_82_n 0.0371775f $X=2.16 $Y=4.07 $X2=0.455 $Y2=0.565
cc_30 N_VPB_X0_noxref_D1 N_VPWR_c_85_n 0.113624f $X=-0.33 $Y=1.885 $X2=0.577
+ $Y2=1.07
cc_31 VPB N_VPWR_c_85_n 0.0155031f $X=0 $Y=3.955 $X2=0.577 $Y2=1.07
cc_32 N_VPB_c_22_p N_VPWR_c_85_n 0.0243396f $X=2.16 $Y=4.07 $X2=0.577 $Y2=1.07
cc_33 N_VPB_X0_noxref_D1 N_LO_c_127_n 0.151962f $X=-0.33 $Y=1.885 $X2=0.84
+ $Y2=1.82
cc_34 N_VPB_X0_noxref_D1 N_LO_c_132_n 0.0118858f $X=-0.33 $Y=1.885 $X2=0.577
+ $Y2=0.565
cc_35 VPB N_LO_c_132_n 0.00277232f $X=0 $Y=3.955 $X2=0.577 $Y2=0.565
cc_36 N_VPB_c_22_p N_LO_c_132_n 0.0391267f $X=2.16 $Y=4.07 $X2=0.577 $Y2=0.565
cc_37 N_VPB_X0_noxref_D1 N_LO_c_135_n 0.122676f $X=-0.33 $Y=1.885 $X2=0.455
+ $Y2=0.565
cc_38 VPB N_LO_c_135_n 0.0155031f $X=0 $Y=3.955 $X2=0.455 $Y2=0.565
cc_39 N_VPB_c_22_p N_LO_c_135_n 0.0241291f $X=2.16 $Y=4.07 $X2=0.455 $Y2=0.565
cc_40 N_HI_c_49_p N_VPWR_c_77_n 0.00639527f $X=0.74 $Y=1.935 $X2=0 $Y2=0
cc_41 HI N_VPWR_c_77_n 0.0488317f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_42 HI N_VPWR_c_77_n 0.0539637f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_43 HI VPWR 0.0227576f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_44 HI N_VPWR_c_82_n 0.0135149f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_45 HI N_VPWR_c_85_n 0.0114027f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_46 N_HI_R0_pos N_VGND_R1_pos 0.0468073f $X=0.84 $Y=1.82 $X2=0 $Y2=0
cc_47 N_HI_c_49_p N_VGND_R1_pos 6.15994e-19 $X=0.74 $Y=1.935 $X2=0 $Y2=0
cc_48 N_HI_c_41_n N_VGND_c_103_n 5.39121e-19 $X=0.455 $Y=0.565 $X2=0.24 $Y2=0
cc_49 N_HI_c_43_n N_VGND_c_103_n 0.0468073f $X=0.84 $Y=0.735 $X2=0.24 $Y2=0
cc_50 N_HI_c_43_n N_VGND_c_105_n 2.23249e-19 $X=0.84 $Y=0.735 $X2=0.24 $Y2=0
cc_51 N_HI_c_41_n N_VGND_c_106_n 5.8995e-19 $X=0.455 $Y=0.565 $X2=2.16 $Y2=0
cc_52 N_HI_c_43_n N_VGND_c_106_n 5.78764e-19 $X=0.84 $Y=0.735 $X2=2.16 $Y2=0
cc_53 N_HI_c_41_n N_VGND_c_108_n 0.0574565f $X=0.455 $Y=0.565 $X2=2.16 $Y2=0
cc_54 N_HI_c_43_n N_VGND_c_108_n 0.0194647f $X=0.84 $Y=0.735 $X2=2.16 $Y2=0
cc_55 N_HI_c_49_p N_LO_c_127_n 2.01985e-19 $X=0.74 $Y=1.935 $X2=0 $Y2=0
cc_56 HI N_LO_c_127_n 0.0068883f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_57 HI N_LO_c_127_n 0.0260954f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_58 HI N_LO_c_135_n 0.00908035f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_59 N_HI_R0_pos LO 0.0126907f $X=0.84 $Y=1.82 $X2=0 $Y2=0
cc_60 N_HI_c_41_n LO 0.0745733f $X=0.455 $Y=0.565 $X2=0 $Y2=0
cc_61 N_HI_c_43_n LO 0.016085f $X=0.84 $Y=0.735 $X2=0 $Y2=0
cc_62 N_HI_R0_pos LO 0.00822143f $X=0.84 $Y=1.82 $X2=0 $Y2=0
cc_63 N_HI_c_49_p LO 0.0205809f $X=0.74 $Y=1.935 $X2=0 $Y2=0
cc_64 HI LO 0.0225842f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_65 N_HI_c_49_p LO 0.00429459f $X=0.74 $Y=1.935 $X2=0 $Y2=0
cc_66 HI LO 0.0168217f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_67 HI LO 0.083884f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_68 N_VPWR_c_77_n N_LO_c_127_n 0.0660389f $X=0.84 $Y=3.175 $X2=0 $Y2=0
cc_69 VPWR N_LO_c_132_n 0.0706387f $X=0 $Y=3.445 $X2=-0.33 $Y2=-0.265
cc_70 N_VPWR_c_82_n N_LO_c_132_n 0.00218825f $X=0.455 $Y=3.34 $X2=-0.33
+ $Y2=-0.265
cc_71 N_VPWR_c_85_n N_LO_c_132_n 0.00152479f $X=0.84 $Y=3.51 $X2=-0.33
+ $Y2=-0.265
cc_72 VPWR N_LO_c_135_n 0.0183133f $X=0 $Y=3.445 $X2=0 $Y2=0
cc_73 N_VPWR_c_82_n N_LO_c_135_n 0.00109474f $X=0.455 $Y=3.34 $X2=0 $Y2=0
cc_74 N_VPWR_c_85_n N_LO_c_135_n 0.0660389f $X=0.84 $Y=3.51 $X2=0 $Y2=0
cc_75 N_VPWR_c_77_n LO 8.00354e-19 $X=0.84 $Y=3.175 $X2=0 $Y2=0
cc_76 N_VGND_R1_pos LO 0.0257746f $X=1.56 $Y=1.82 $X2=0 $Y2=0
cc_77 N_VGND_c_103_n LO 0.0200561f $X=1.945 $Y=0.565 $X2=0 $Y2=0
cc_78 N_VGND_c_105_n LO 0.0165104f $X=1.945 $Y=0.565 $X2=0 $Y2=0
cc_79 N_VGND_c_106_n LO 0.00816771f $X=2.04 $Y=0.48 $X2=0 $Y2=0
cc_80 N_VGND_c_108_n LO 0.0307914f $X=2.04 $Y=0.48 $X2=0 $Y2=0
cc_81 N_VGND_R1_pos LO 0.0491992f $X=1.56 $Y=1.82 $X2=0 $Y2=0
cc_82 N_VGND_c_105_n LO 5.00804e-19 $X=1.945 $Y=0.565 $X2=0 $Y2=0
cc_83 N_VGND_R1_pos LO 0.00529894f $X=1.56 $Y=1.82 $X2=0 $Y2=0
