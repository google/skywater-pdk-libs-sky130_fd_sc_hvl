* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbufhv2lv_simple_1 A LVPWR VGND VNB VPB VPWR X
M1000 a_762_107# a_662_81# X VNB nhv w=750000u l=500000u
+  ad=3.0405e+11p pd=2.5e+06u as=1.9875e+11p ps=2.03e+06u
M1001 LVPWR a_662_81# X LVPWR phv w=1.5e+06u l=500000u
+  ad=5.1e+11p pd=3.79e+06u as=4.275e+11p ps=3.57e+06u
M1002 a_662_81# A a_762_107# VNB nhv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1003 a_662_81# A LVPWR LVPWR phv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
.ends
