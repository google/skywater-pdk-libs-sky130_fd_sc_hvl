* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 VPWR SCE a_116_451# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 VGND SCE a_116_451# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_1510_100# a_1212_471# a_2360_115# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_2574_543# a_2616_417# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 VGND RESET_B a_2904_181# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_1212_100# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VGND a_3417_443# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X7 a_294_126# SCE a_65_649# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR a_3417_443# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_1610_126# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_3417_443# a_2360_115# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 a_524_649# D a_65_649# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_2360_115# a_1212_100# a_2539_181# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 a_137_126# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 a_2539_181# a_2616_417# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 a_222_649# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X16 VPWR CLK a_1212_100# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X17 a_65_649# RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X18 a_1468_641# a_1510_100# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 VPWR RESET_B a_2616_417# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 a_3417_443# a_2360_115# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X21 a_65_649# a_116_451# a_592_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 a_1312_126# a_1212_100# a_1468_641# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X23 VPWR a_1312_126# a_1510_100# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X24 VGND a_1312_126# a_1510_100# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X25 a_1468_126# a_1510_100# a_1610_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X26 a_2904_181# a_2360_115# a_2616_417# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 VPWR SCE a_524_649# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X28 a_65_649# a_1212_471# a_1312_126# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X29 VPWR RESET_B a_1312_126# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X30 a_2360_115# a_1212_471# a_2574_543# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X31 a_1212_471# a_1212_100# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X32 a_1312_126# a_1212_471# a_1468_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X33 a_1212_471# a_1212_100# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X34 a_137_126# SCD a_294_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X35 a_65_649# a_116_451# a_222_649# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X36 a_2616_417# a_2360_115# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X37 a_65_649# a_1212_100# a_1312_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X38 a_592_126# D a_137_126# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X39 a_1510_100# a_1212_100# a_2360_115# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
.ends
