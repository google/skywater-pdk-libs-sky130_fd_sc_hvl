# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__diode_2
  CLASS CORE ANTENNACELL ;
  FOREIGN sky130_fd_sc_hvl__diode_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.960000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN DIODE
    ANTENNADIFFAREA  0.607200 ;
    ANTENNAGATEAREA  0.607200 ;
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.515000 0.855000 3.280000 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 0.960000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 0.960000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 0.960000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 0.960000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.960000 0.085000 ;
      RECT 0.000000  3.985000 0.960000 4.155000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
  END
END sky130_fd_sc_hvl__diode_2
END LIBRARY
