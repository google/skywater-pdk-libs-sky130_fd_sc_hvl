* File: sky130_fd_sc_hvl__inv_1.pxi.spice
* Created: Fri Aug 28 09:35:59 2020
* 
x_PM_SKY130_FD_SC_HVL__INV_1%VNB N_VNB_M1001_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__INV_1%VNB
x_PM_SKY130_FD_SC_HVL__INV_1%VPB N_VPB_M1000_b VPB N_VPB_c_13_p VPB
+ PM_SKY130_FD_SC_HVL__INV_1%VPB
x_PM_SKY130_FD_SC_HVL__INV_1%A N_A_M1000_g N_A_M1001_g A A N_A_c_30_n
+ PM_SKY130_FD_SC_HVL__INV_1%A
x_PM_SKY130_FD_SC_HVL__INV_1%VPWR N_VPWR_M1000_s VPWR N_VPWR_c_52_n
+ PM_SKY130_FD_SC_HVL__INV_1%VPWR
x_PM_SKY130_FD_SC_HVL__INV_1%Y N_Y_M1001_d N_Y_M1000_d Y Y Y Y Y Y Y N_Y_c_60_n
+ Y PM_SKY130_FD_SC_HVL__INV_1%Y
x_PM_SKY130_FD_SC_HVL__INV_1%VGND N_VGND_M1001_s VGND N_VGND_c_80_n
+ PM_SKY130_FD_SC_HVL__INV_1%VGND
cc_1 N_VNB_M1001_b N_A_M1001_g 0.0551724f $X=-0.33 $Y=-0.265 $X2=0.755 $Y2=0.91
cc_2 N_VNB_c_2_p N_A_M1001_g 0.0015174f $X=0.24 $Y=0 $X2=0.755 $Y2=0.91
cc_3 N_VNB_M1001_b A 0.019602f $X=-0.33 $Y=-0.265 $X2=0.635 $Y2=1.58
cc_4 N_VNB_M1001_b N_A_c_30_n 0.0545387f $X=-0.33 $Y=-0.265 $X2=0.67 $Y2=1.77
cc_5 N_VNB_M1001_b N_Y_c_60_n 0.0741071f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_c_2_p N_Y_c_60_n 7.68678e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_7 N_VNB_M1001_b VGND 0.0512888f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_8 N_VNB_c_2_p VGND 0.154031f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_9 N_VNB_M1001_b N_VGND_c_80_n 0.0710585f $X=-0.33 $Y=-0.265 $X2=0.755
+ $Y2=0.91
cc_10 N_VNB_c_2_p N_VGND_c_80_n 0.00166879f $X=0.24 $Y=0 $X2=0.755 $Y2=0.91
cc_11 N_VPB_M1000_b N_A_M1000_g 0.0451728f $X=-0.33 $Y=1.885 $X2=0.735 $Y2=2.965
cc_12 VPB N_A_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.735 $Y2=2.965
cc_13 N_VPB_c_13_p N_A_M1000_g 0.0170743f $X=1.2 $Y=4.07 $X2=0.735 $Y2=2.965
cc_14 N_VPB_M1000_b A 0.0061311f $X=-0.33 $Y=1.885 $X2=0.635 $Y2=1.58
cc_15 N_VPB_M1000_b N_A_c_30_n 0.0258169f $X=-0.33 $Y=1.885 $X2=0.67 $Y2=1.77
cc_16 N_VPB_M1000_b VPWR 0.0405637f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_17 VPB VPWR 0.153123f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_18 N_VPB_c_13_p VPWR 0.00690123f $X=1.2 $Y=4.07 $X2=0 $Y2=0
cc_19 N_VPB_M1000_b N_VPWR_c_52_n 0.0684885f $X=-0.33 $Y=1.885 $X2=0.755
+ $Y2=0.91
cc_20 VPB N_VPWR_c_52_n 0.00213862f $X=0 $Y=3.955 $X2=0.755 $Y2=0.91
cc_21 N_VPB_c_13_p N_VPWR_c_52_n 0.0303036f $X=1.2 $Y=4.07 $X2=0.755 $Y2=0.91
cc_22 N_VPB_M1000_b Y 0.00859775f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_23 N_VPB_M1000_b N_Y_c_60_n 0.0159301f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_24 N_VPB_M1000_b Y 0.0504529f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_25 VPB Y 0.0012155f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_26 N_VPB_c_13_p Y 0.0201437f $X=1.2 $Y=4.07 $X2=0 $Y2=0
cc_27 N_A_M1000_g VPWR 0.0168776f $X=0.735 $Y=2.965 $X2=0 $Y2=0
cc_28 N_A_M1000_g N_VPWR_c_52_n 0.0641117f $X=0.735 $Y=2.965 $X2=0 $Y2=0
cc_29 A N_VPWR_c_52_n 0.0371565f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_30 N_A_M1000_g Y 0.00604919f $X=0.735 $Y=2.965 $X2=0.24 $Y2=0
cc_31 N_A_c_30_n Y 0.0010557f $X=0.67 $Y=1.77 $X2=0.24 $Y2=0
cc_32 N_A_M1000_g N_Y_c_60_n 0.0044012f $X=0.735 $Y=2.965 $X2=0.72 $Y2=0.058
cc_33 N_A_M1001_g N_Y_c_60_n 0.0362734f $X=0.755 $Y=0.91 $X2=0.72 $Y2=0.058
cc_34 A N_Y_c_60_n 0.030872f $X=0.635 $Y=1.58 $X2=0.72 $Y2=0.058
cc_35 N_A_M1000_g Y 0.0293331f $X=0.735 $Y=2.965 $X2=0 $Y2=0
cc_36 N_A_M1001_g VGND 0.0211718f $X=0.755 $Y=0.91 $X2=0 $Y2=0
cc_37 N_A_M1001_g N_VGND_c_80_n 0.0418762f $X=0.755 $Y=0.91 $X2=0 $Y2=0
cc_38 A N_VGND_c_80_n 0.0390377f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_39 N_A_c_30_n N_VGND_c_80_n 6.20505e-19 $X=0.67 $Y=1.77 $X2=0 $Y2=0
cc_40 N_VPWR_c_52_n Y 0.07917f $X=0.345 $Y=2.34 $X2=0 $Y2=0
cc_41 VPWR Y 0.0492493f $X=0 $Y=3.445 $X2=0 $Y2=0
cc_42 N_Y_M1001_d VGND 3.33633e-19 $X=1.005 $Y=0.535 $X2=0 $Y2=0
cc_43 N_Y_c_60_n VGND 0.034001f $X=1.145 $Y=0.66 $X2=0 $Y2=0
cc_44 N_Y_c_60_n N_VGND_c_80_n 0.021149f $X=1.145 $Y=0.66 $X2=0 $Y2=0
