* File: sky130_fd_sc_hvl__einvp_1.spice
* Created: Wed Sep  2 09:06:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__einvp_1.pex.spice"
.subckt sky130_fd_sc_hvl__einvp_1  VNB VPB TE A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE	TE
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_TE_M1005_g N_A_30_189#_M1005_s N_VNB_M1005_b NHV L=0.5
+ W=0.42 AD=0.128746 AS=0.1197 PD=0.990769 PS=1.41 NRD=68.2746 NRS=0 M=1 R=0.84
+ SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1001 A_413_123# N_TE_M1001_g N_VGND_M1005_d N_VNB_M1005_b NHV L=0.5 W=0.75
+ AD=0.135 AS=0.229904 PD=1.11 PS=1.76923 NRD=18.9924 NRS=0 M=1 R=1.5 SA=250001
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1003 N_Z_M1003_d N_A_M1003_g A_413_123# N_VNB_M1005_b NHV L=0.5 W=0.75
+ AD=0.21375 AS=0.135 PD=2.07 PS=1.11 NRD=0 NRS=18.9924 M=1 R=1.5 SA=250002
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1002 N_VPWR_M1002_d N_TE_M1002_g N_A_30_189#_M1002_s N_VPB_M1002_b PHV L=0.5
+ W=0.75 AD=0.16625 AS=0.21375 PD=1.25333 PS=2.07 NRD=25.4603 NRS=0 M=1 R=1.5
+ SA=250000 SB=250002 A=0.375 P=2.5 MULT=1
MM1004 A_413_443# N_A_30_189#_M1004_g N_VPWR_M1002_d N_VPB_M1002_b PHV L=0.5
+ W=1.5 AD=0.27 AS=0.3325 PD=1.86 PS=2.50667 NRD=15.9103 NRS=0 M=1 R=3 SA=250000
+ SB=250001 A=0.75 P=4 MULT=1
MM1000 N_Z_M1000_d N_A_M1000_g A_413_443# N_VPB_M1002_b PHV L=0.5 W=1.5
+ AD=0.4275 AS=0.27 PD=3.57 PS=1.86 NRD=0 NRS=15.9103 M=1 R=3 SA=250001
+ SB=250000 A=0.75 P=4 MULT=1
DX6_noxref N_VNB_M1005_b N_VPB_M1002_b NWDIODE A=10.452 P=13.24
*
.include "sky130_fd_sc_hvl__einvp_1.pxi.spice"
*
.ends
*
*
