* File: sky130_fd_sc_hvl__nor2_1.spice
* Created: Fri Aug 28 09:38:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__nor2_1.pex.spice"
.subckt sky130_fd_sc_hvl__nor2_1  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1002_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.21375 PD=1.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5 SA=250000 SB=250001
+ A=0.375 P=2.5 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g N_Y_M1002_d N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.21375 AS=0.105 PD=2.07 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250001 SB=250000
+ A=0.375 P=2.5 MULT=1
MM1000 A_251_443# N_A_M1000_g N_VPWR_M1000_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.1575 AS=0.4275 PD=1.71 PS=3.57 NRD=6.3603 NRS=0 M=1 R=3 SA=250000
+ SB=250001 A=0.75 P=4 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g A_251_443# N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.4275 AS=0.1575 PD=3.57 PS=1.71 NRD=0 NRS=6.3603 M=1 R=3 SA=250001
+ SB=250000 A=0.75 P=4 MULT=1
DX4_noxref N_VNB_M1002_b N_VPB_M1000_b NWDIODE A=7.956 P=11.32
*
.include "sky130_fd_sc_hvl__nor2_1.pxi.spice"
*
.ends
*
*
