* File: sky130_fd_sc_hvl__mux2_1.spice
* Created: Wed Sep  2 09:08:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__mux2_1.pex.spice"
.subckt sky130_fd_sc_hvl__mux2_1  VNB VPB S A0 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A0	A0
* S	S
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_94_81#_M1009_g N_X_M1009_s N_VNB_M1009_b NHV L=0.5
+ W=0.75 AD=0.166635 AS=0.21375 PD=1.46795 PS=2.07 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250002 A=0.375 P=2.5 MULT=1
MM1001 A_373_107# N_S_M1001_g N_VGND_M1009_d N_VNB_M1009_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0933154 PD=0.63 PS=0.822051 NRD=13.566 NRS=31.2132 M=1 R=0.84
+ SA=250001 SB=250003 A=0.21 P=1.84 MULT=1
MM1006 N_A_94_81#_M1006_d N_A1_M1006_g A_373_107# N_VNB_M1009_b NHV L=0.5 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250002
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1011 A_671_107# N_A0_M1011_g N_A_94_81#_M1006_d N_VNB_M1009_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84 SA=250002
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1003 N_VGND_M1003_d N_A_713_81#_M1003_g A_671_107# N_VNB_M1009_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250003 SB=250001 A=0.21 P=1.84 MULT=1
MM1008 N_A_713_81#_M1008_d N_S_M1008_g N_VGND_M1003_d N_VNB_M1009_b NHV L=0.5
+ W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250004
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1002 N_VPWR_M1002_d N_A_94_81#_M1002_g N_X_M1002_s N_VPB_M1002_b PHV L=0.5
+ W=1.5 AD=0.370078 AS=0.4275 PD=2.96094 PS=3.57 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250001 A=0.75 P=4 MULT=1
MM1004 A_373_491# N_S_M1004_g N_VPWR_M1002_d N_VPB_M1002_b PHV L=0.5 W=0.42
+ AD=0.0441 AS=0.103622 PD=0.63 PS=0.829062 NRD=22.729 NRS=52.2958 M=1 R=0.84
+ SA=250001 SB=250003 A=0.21 P=1.84 MULT=1
MM1007 N_A_94_81#_M1007_d N_A0_M1007_g A_373_491# N_VPB_M1002_b PHV L=0.5 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84 SA=250002
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1000 A_671_491# N_A1_M1000_g N_A_94_81#_M1007_d N_VPB_M1002_b PHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84 SA=250002
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1005 N_VPWR_M1005_d N_A_713_81#_M1005_g A_671_491# N_VPB_M1002_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250003 SB=250001 A=0.21 P=1.84 MULT=1
MM1010 N_A_713_81#_M1010_d N_S_M1010_g N_VPWR_M1005_d N_VPB_M1002_b PHV L=0.5
+ W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250004
+ SB=250000 A=0.21 P=1.84 MULT=1
DX12_noxref N_VNB_M1009_b N_VPB_M1002_b NWDIODE A=15.444 P=17.08
*
.include "sky130_fd_sc_hvl__mux2_1.pxi.spice"
*
.ends
*
*
