* File: sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1.pex.spice
* Created: Wed Sep  2 09:07:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%VNB 9 11 12 23 35 42 49
r108 29 49 4.1576 $w=2.3e-07 $l=6.48e-06 $layer=MET1_cond $X=0.24 $Y=8.14
+ $X2=6.72 $Y2=8.14
r109 17 42 4.1576 $w=2.3e-07 $l=6.48e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=6.72
+ $Y2=0
r110 12 35 4.31158 $w=2.3e-07 $l=6.72e-06 $layer=MET1_cond $X=6.96 $Y=8.14
+ $X2=13.68 $Y2=8.14
r111 12 49 0.153985 $w=2.3e-07 $l=2.4e-07 $layer=MET1_cond $X=6.96 $Y=8.14
+ $X2=6.72 $Y2=8.14
r112 11 23 4.31158 $w=2.3e-07 $l=6.72e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=13.68 $Y2=0
r113 11 42 0.153985 $w=2.3e-07 $l=2.4e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.72
+ $Y2=0
r114 9 35 0.641379 $w=1.7e-07 $l=2.465e-06 $layer=mcon $count=14 $X=13.68
+ $Y=8.14 $X2=13.68 $Y2=8.14
r115 9 29 0.641379 $w=1.7e-07 $l=2.465e-06 $layer=mcon $count=14 $X=0.24 $Y=8.14
+ $X2=0.24 $Y2=8.14
r116 9 23 0.641379 $w=1.7e-07 $l=2.465e-06 $layer=mcon $count=14 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r117 9 17 0.641379 $w=1.7e-07 $l=2.465e-06 $layer=mcon $count=14 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%VPB 4 8 10 12 20 27
c78 10 0 2.72384e-19 $X=0 $Y=3.955
r79 21 27 3.92662 $w=2.3e-07 $l=6.12e-06 $layer=MET1_cond $X=0.6 $Y=4.07
+ $X2=6.72 $Y2=4.07
r80 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.6 $Y=4.07 $X2=0.6
+ $Y2=4.07
r81 18 20 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.445 $Y=4.07
+ $X2=0.6 $Y2=4.07
r82 15 21 0.230978 $w=2.3e-07 $l=3.6e-07 $layer=MET1_cond $X=0.24 $Y=4.07
+ $X2=0.6 $Y2=4.07
r83 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r84 12 18 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.36 $Y=4.07
+ $X2=0.445 $Y2=4.07
r85 12 14 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.36 $Y=4.07
+ $X2=0.24 $Y2=4.07
r86 10 27 0.153985 $w=2.3e-07 $l=2.4e-07 $layer=MET1_cond $X=6.96 $Y=4.07
+ $X2=6.72 $Y2=4.07
r87 6 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.445 $Y=4.155
+ $X2=0.445 $Y2=4.07
r88 6 8 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.445 $Y=4.155
+ $X2=0.445 $Y2=4.935
r89 4 14 182 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=1 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
r90 4 8 182 $w=1.7e-07 $l=1.1512e-06 $layer=licon1_NTAP_notbjt $count=1 $X=0
+ $Y=3.985 $X2=0.445 $Y2=4.935
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%LVPWR 1 2 10 16 19 22 27
+ 28 34 35 38
c63 34 0 1.02552e-19 $X=9.78 $Y=3.165
r64 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.78 $Y=3.165
+ $X2=9.78 $Y2=3.165
r65 28 35 1.4055 $w=2.85e-07 $l=2.82e-06 $layer=MET1_cond $X=6.96 $Y=3.162
+ $X2=9.78 $Y2=3.162
r66 28 38 0.119617 $w=2.85e-07 $l=2.4e-07 $layer=MET1_cond $X=6.96 $Y=3.162
+ $X2=6.72 $Y2=3.162
r67 22 24 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=9.87 $Y=4.94 $X2=9.87
+ $Y2=5.64
r68 20 27 5.16603 $w=3.3e-07 $l=1.96914e-07 $layer=LI1_cond $X=9.87 $Y=4.235
+ $X2=9.8 $Y2=4.07
r69 20 22 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=9.87 $Y=4.235
+ $X2=9.87 $Y2=4.94
r70 19 27 5.16603 $w=3.3e-07 $l=1.96914e-07 $layer=LI1_cond $X=9.73 $Y=3.905
+ $X2=9.8 $Y2=4.07
r71 18 19 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=9.73 $Y=3.365
+ $X2=9.73 $Y2=3.905
r72 14 34 1.67021 $w=3.43e-07 $l=5e-08 $layer=LI1_cond $X=9.73 $Y=3.192 $X2=9.78
+ $Y2=3.192
r73 14 18 0.986088 $w=3.3e-07 $l=1.73e-07 $layer=LI1_cond $X=9.73 $Y=3.192
+ $X2=9.73 $Y2=3.365
r74 14 16 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=9.73 $Y=3.02
+ $X2=9.73 $Y2=2.5
r75 10 27 91 $w=1.7e-07 $l=6.36082e-07 $layer=licon1_NTAP_notbjt $count=2 $X=9.1
+ $Y=3.985 $X2=9.695 $Y2=4.07
r76 2 24 400 $w=1.7e-07 $l=9.39694e-07 $layer=licon1_PDIFF $count=1 $X=9.67
+ $Y=4.795 $X2=9.87 $Y2=5.64
r77 2 22 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=9.67
+ $Y=4.795 $X2=9.87 $Y2=4.94
r78 1 14 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=9.585
+ $Y=2.225 $X2=9.73 $Y2=3.2
r79 1 16 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=9.585
+ $Y=2.225 $X2=9.73 $Y2=2.5
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_229_967# 1 2 9 12 13 15
+ 18 22 26 30 33 35 36 37
r71 37 38 29.436 $w=8.9e-07 $l=3.4e-07 $layer=POLY_cond $X=1.59 $Y=5.175
+ $X2=1.59 $Y2=4.835
r72 34 37 31.4858 $w=8.9e-07 $l=5.45e-07 $layer=POLY_cond $X=1.59 $Y=5.72
+ $X2=1.59 $Y2=5.175
r73 33 35 7.04571 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.87 $Y=5.72
+ $X2=2.035 $Y2=5.72
r74 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.87
+ $Y=5.72 $X2=1.87 $Y2=5.72
r75 28 30 29.073 $w=2.18e-07 $l=5.55e-07 $layer=LI1_cond $X=5.565 $Y=5.665
+ $X2=5.565 $Y2=5.11
r76 27 36 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=3.515 $Y=5.775
+ $X2=3.405 $Y2=5.775
r77 26 28 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=5.455 $Y=5.775
+ $X2=5.565 $Y2=5.665
r78 26 27 101.625 $w=2.18e-07 $l=1.94e-06 $layer=LI1_cond $X=5.455 $Y=5.775
+ $X2=3.515 $Y2=5.775
r79 22 24 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=3.405 $Y=6.61
+ $X2=3.405 $Y2=7.29
r80 20 36 1.34256 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=3.405 $Y=5.885
+ $X2=3.405 $Y2=5.775
r81 20 22 37.9782 $w=2.18e-07 $l=7.25e-07 $layer=LI1_cond $X=3.405 $Y=5.885
+ $X2=3.405 $Y2=6.61
r82 18 36 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=3.295 $Y=5.775
+ $X2=3.405 $Y2=5.775
r83 18 35 66.0036 $w=2.18e-07 $l=1.26e-06 $layer=LI1_cond $X=3.295 $Y=5.775
+ $X2=2.035 $Y2=5.775
r84 13 37 9.1487 $w=6.8e-07 $l=4.45e-07 $layer=POLY_cond $X=2.035 $Y=5.175
+ $X2=1.59 $Y2=5.175
r85 13 15 7.79706 $w=6.8e-07 $l=1.1e-07 $layer=POLY_cond $X=2.035 $Y=5.175
+ $X2=2.145 $Y2=5.175
r86 12 38 217.757 $w=5e-07 $l=2.035e-06 $layer=POLY_cond $X=1.455 $Y=2.8
+ $X2=1.455 $Y2=4.835
r87 9 12 161.579 $w=5e-07 $l=1.51e-06 $layer=POLY_cond $X=1.455 $Y=1.29
+ $X2=1.455 $Y2=2.8
r88 2 30 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.425
+ $Y=4.965 $X2=5.565 $Y2=5.11
r89 1 24 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1 $X=3.265
+ $Y=6.465 $X2=3.405 $Y2=7.29
r90 1 22 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.265
+ $Y=6.465 $X2=3.405 $Y2=6.61
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_507_107# 1 2 9 13 17 22
+ 24 25 27
c37 17 0 1.87386e-19 $X=4.315 $Y=2.57
r38 23 27 53.3453 $w=8e-07 $l=8.3e-07 $layer=POLY_cond $X=2.935 $Y=1.995
+ $X2=2.935 $Y2=1.165
r39 22 24 7.04571 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=1.995
+ $X2=3.32 $Y2=1.995
r40 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.155
+ $Y=1.995 $X2=3.155 $Y2=1.995
r41 17 19 53.4314 $w=2.18e-07 $l=1.02e-06 $layer=LI1_cond $X=4.315 $Y=2.57
+ $X2=4.315 $Y2=3.59
r42 15 25 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.315 $Y=2.16
+ $X2=4.315 $Y2=2.05
r43 15 17 21.4773 $w=2.18e-07 $l=4.1e-07 $layer=LI1_cond $X=4.315 $Y=2.16
+ $X2=4.315 $Y2=2.57
r44 11 25 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.315 $Y=1.94
+ $X2=4.315 $Y2=2.05
r45 11 13 59.1937 $w=2.18e-07 $l=1.13e-06 $layer=LI1_cond $X=4.315 $Y=1.94
+ $X2=4.315 $Y2=0.81
r46 9 25 1.34256 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.205 $Y=2.05
+ $X2=4.315 $Y2=2.05
r47 9 24 46.3596 $w=2.18e-07 $l=8.85e-07 $layer=LI1_cond $X=4.205 $Y=2.05
+ $X2=3.32 $Y2=2.05
r48 2 19 300 $w=1.7e-07 $l=1.23301e-06 $layer=licon1_PDIFF $count=2 $X=4.175
+ $Y=2.425 $X2=4.315 $Y2=3.59
r49 2 17 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.175
+ $Y=2.425 $X2=4.315 $Y2=2.57
r50 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.175
+ $Y=0.665 $X2=4.315 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_176_993# 1 2 3 12 13 18
+ 20 21 22 25 31 36 40 41 45
r87 38 41 1.31569 $w=4.98e-07 $l=5.5e-08 $layer=LI1_cond $X=2.615 $Y=4.545
+ $X2=2.67 $Y2=4.545
r88 38 40 15.8918 $w=4.98e-07 $l=5.05e-07 $layer=LI1_cond $X=2.615 $Y=4.545
+ $X2=2.11 $Y2=4.545
r89 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.615
+ $Y=4.46 $X2=2.615 $Y2=4.46
r90 36 41 5.5681 $w=2.2e-07 $l=2.5e-07 $layer=LI1_cond $X=2.67 $Y=4.295 $X2=2.67
+ $Y2=4.545
r91 35 45 0.853166 $w=2.2e-07 $l=1.13e-07 $layer=LI1_cond $X=2.67 $Y=3.085
+ $X2=2.67 $Y2=2.972
r92 35 36 63.3844 $w=2.18e-07 $l=1.21e-06 $layer=LI1_cond $X=2.67 $Y=3.085
+ $X2=2.67 $Y2=4.295
r93 31 34 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=2.37 $Y=0.81 $X2=2.37
+ $Y2=1.49
r94 29 45 15.3659 $w=2.23e-07 $l=3e-07 $layer=LI1_cond $X=2.37 $Y=2.972 $X2=2.67
+ $Y2=2.972
r95 29 34 71.7658 $w=2.18e-07 $l=1.37e-06 $layer=LI1_cond $X=2.37 $Y=2.86
+ $X2=2.37 $Y2=1.49
r96 25 27 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=1.845 $Y=6.61
+ $X2=1.845 $Y2=7.29
r97 23 25 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=1.845 $Y=6.275
+ $X2=1.845 $Y2=6.61
r98 21 23 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=1.735 $Y=6.165
+ $X2=1.845 $Y2=6.275
r99 21 22 32.4779 $w=2.18e-07 $l=6.2e-07 $layer=LI1_cond $X=1.735 $Y=6.165
+ $X2=1.115 $Y2=6.165
r100 20 40 52.1219 $w=2.18e-07 $l=9.95e-07 $layer=LI1_cond $X=1.115 $Y=4.685
+ $X2=2.11 $Y2=4.685
r101 16 22 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=1.005 $Y=6.055
+ $X2=1.115 $Y2=6.165
r102 16 18 49.5027 $w=2.18e-07 $l=9.45e-07 $layer=LI1_cond $X=1.005 $Y=6.055
+ $X2=1.005 $Y2=5.11
r103 15 20 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=1.005 $Y=4.795
+ $X2=1.115 $Y2=4.685
r104 15 18 16.5009 $w=2.18e-07 $l=3.15e-07 $layer=LI1_cond $X=1.005 $Y=4.795
+ $X2=1.005 $Y2=5.11
r105 13 39 141.638 $w=3.3e-07 $l=8.1e-07 $layer=POLY_cond $X=3.425 $Y=4.46
+ $X2=2.615 $Y2=4.46
r106 12 13 73.1039 $w=1.22e-06 $l=1e-06 $layer=POLY_cond $X=4.425 $Y=4.905
+ $X2=3.425 $Y2=4.905
r107 3 18 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.88
+ $Y=4.965 $X2=1.005 $Y2=5.11
r108 2 34 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.665 $X2=2.395 $Y2=1.49
r109 2 31 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.665 $X2=2.395 $Y2=0.81
r110 1 27 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1
+ $X=1.705 $Y=6.465 $X2=1.845 $Y2=7.29
r111 1 25 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1
+ $X=1.705 $Y=6.465 $X2=1.845 $Y2=6.61
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%SLEEP_B 3 7 9 12 13 14 17
+ 19 21 23 27 31
r58 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.235
+ $Y=1.995 $X2=5.235 $Y2=1.995
r59 27 31 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.065 $Y=1.995
+ $X2=5.235 $Y2=1.995
r60 19 21 234.521 $w=6e-07 $l=2.63e-06 $layer=POLY_cond $X=7.895 $Y=1.195
+ $X2=7.895 $Y2=3.825
r61 15 19 153.878 $w=3.3e-07 $l=8.8e-07 $layer=POLY_cond $X=7.015 $Y=1.03
+ $X2=7.895 $Y2=1.03
r62 15 17 234.521 $w=6e-07 $l=2.63e-06 $layer=POLY_cond $X=7.015 $Y=1.195
+ $X2=7.015 $Y2=3.825
r63 13 15 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=6.715 $Y=1.03
+ $X2=7.015 $Y2=1.03
r64 13 14 229.943 $w=3.3e-07 $l=1.315e-06 $layer=POLY_cond $X=6.715 $Y=1.03
+ $X2=5.4 $Y2=1.03
r65 12 30 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.235 $Y=1.83
+ $X2=5.235 $Y2=1.995
r66 11 14 26.9307 $w=3.3e-07 $l=2.33345e-07 $layer=POLY_cond $X=5.235 $Y=1.195
+ $X2=5.4 $Y2=1.03
r67 11 12 111.037 $w=3.3e-07 $l=6.35e-07 $layer=POLY_cond $X=5.235 $Y=1.195
+ $X2=5.235 $Y2=1.83
r68 10 23 11.3528 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=4.175 $Y=1.995
+ $X2=3.925 $Y2=1.995
r69 9 30 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.07 $Y=1.995
+ $X2=5.235 $Y2=1.995
r70 9 10 156.501 $w=3.3e-07 $l=8.95e-07 $layer=POLY_cond $X=5.07 $Y=1.995
+ $X2=4.175 $Y2=1.995
r71 5 23 14.2643 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.925 $Y=2.16
+ $X2=3.925 $Y2=1.995
r72 5 7 108.611 $w=5e-07 $l=1.015e-06 $layer=POLY_cond $X=3.925 $Y=2.16
+ $X2=3.925 $Y2=3.175
r73 1 23 14.2643 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.925 $Y=1.83
+ $X2=3.925 $Y2=1.995
r74 1 3 84.5347 $w=5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.925 $Y=1.83 $X2=3.925
+ $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_553_1225# 1 2 9 11 12 15
+ 17 20 22 23 24 25 26 29 33
r56 36 38 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=9.37 $Y=5.77
+ $X2=9.37 $Y2=6.79
r57 33 36 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=9.37 $Y=4.94
+ $X2=9.37 $Y2=5.77
r58 31 38 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=9.37 $Y=7.075
+ $X2=9.37 $Y2=6.79
r59 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.255
+ $Y=7.24 $X2=8.255 $Y2=7.24
r60 26 31 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=9.205 $Y=7.24
+ $X2=9.37 $Y2=7.075
r61 26 28 33.1764 $w=3.28e-07 $l=9.5e-07 $layer=LI1_cond $X=9.205 $Y=7.24
+ $X2=8.255 $Y2=7.24
r62 24 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.915 $Y=7.24
+ $X2=8.255 $Y2=7.24
r63 24 25 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.915 $Y=7.24
+ $X2=7.75 $Y2=7.24
r64 22 25 921.242 $w=1.8e-07 $l=2.37e-06 $layer=POLY_cond $X=5.38 $Y=7.315
+ $X2=7.75 $Y2=7.315
r65 20 22 26.9307 $w=1.8e-07 $l=1.27279e-07 $layer=POLY_cond $X=5.29 $Y=7.225
+ $X2=5.38 $Y2=7.315
r66 19 20 357.613 $w=1.8e-07 $l=9.2e-07 $layer=POLY_cond $X=5.29 $Y=6.305
+ $X2=5.29 $Y2=7.225
r67 18 23 43.0828 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=4.045 $Y=6.215
+ $X2=3.795 $Y2=6.215
r68 17 19 26.9307 $w=1.8e-07 $l=1.27279e-07 $layer=POLY_cond $X=5.2 $Y=6.215
+ $X2=5.29 $Y2=6.305
r69 17 18 448.96 $w=1.8e-07 $l=1.155e-06 $layer=POLY_cond $X=5.2 $Y=6.215
+ $X2=4.045 $Y2=6.215
r70 13 23 7.60666 $w=5e-07 $l=9e-08 $layer=POLY_cond $X=3.795 $Y=6.305 $X2=3.795
+ $Y2=6.215
r71 13 15 70.6239 $w=5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.795 $Y=6.305
+ $X2=3.795 $Y2=6.965
r72 11 23 43.0828 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=3.545 $Y=6.215
+ $X2=3.795 $Y2=6.215
r73 11 12 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=3.545 $Y=6.215
+ $X2=3.265 $Y2=6.215
r74 7 12 35.539 $w=1.8e-07 $l=2.91548e-07 $layer=POLY_cond $X=3.015 $Y=6.305
+ $X2=3.265 $Y2=6.215
r75 7 9 70.6239 $w=5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.015 $Y=6.305 $X2=3.015
+ $Y2=6.965
r76 2 36 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=9.225
+ $Y=4.795 $X2=9.37 $Y2=5.77
r77 2 33 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=9.225
+ $Y=4.795 $X2=9.37 $Y2=4.94
r78 1 38 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=9.225
+ $Y=6.645 $X2=9.37 $Y2=6.79
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_241_1225# 1 2 9 11 12 15
+ 18 19 20 22 23 24 26 27 28 31 33 35 36 38 45 50 52 56 57
r111 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.21
+ $Y=6.29 $X2=10.21 $Y2=6.29
r112 52 54 5.27442 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.3 $Y=3.2
+ $X2=10.3 $Y2=3.365
r113 52 53 5.27442 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.3 $Y=3.2
+ $X2=10.3 $Y2=3.035
r114 50 56 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.37 $Y=6.125
+ $X2=10.37 $Y2=6.29
r115 50 54 96.3861 $w=3.28e-07 $l=2.76e-06 $layer=LI1_cond $X=10.37 $Y=6.125
+ $X2=10.37 $Y2=3.365
r116 48 53 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=10.23 $Y=2.37
+ $X2=10.23 $Y2=3.035
r117 45 48 51.3361 $w=3.28e-07 $l=1.47e-06 $layer=LI1_cond $X=10.23 $Y=0.9
+ $X2=10.23 $Y2=2.37
r118 39 40 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.595 $Y=6.365
+ $X2=9.595 $Y2=6.455
r119 38 57 91.8022 $w=3.3e-07 $l=5.25e-07 $layer=POLY_cond $X=9.685 $Y=6.29
+ $X2=10.21 $Y2=6.29
r120 38 39 29.1532 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.595 $Y=6.29
+ $X2=9.595 $Y2=6.365
r121 33 38 118.763 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=9.595 $Y=5.99
+ $X2=9.595 $Y2=6.29
r122 33 35 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.595 $Y=5.99
+ $X2=9.595 $Y2=5.355
r123 31 40 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.585 $Y=7.015
+ $X2=9.585 $Y2=6.455
r124 27 39 2.83073 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.505 $Y=6.365
+ $X2=9.595 $Y2=6.365
r125 27 28 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.505 $Y=6.365
+ $X2=8.93 $Y2=6.365
r126 25 28 26.9307 $w=1.8e-07 $l=1.27279e-07 $layer=POLY_cond $X=8.84 $Y=6.455
+ $X2=8.93 $Y2=6.365
r127 25 26 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=8.84 $Y=6.455
+ $X2=8.84 $Y2=6.665
r128 23 26 26.9307 $w=1.8e-07 $l=1.27279e-07 $layer=POLY_cond $X=8.75 $Y=6.755
+ $X2=8.84 $Y2=6.665
r129 23 24 1158.35 $w=1.8e-07 $l=2.98e-06 $layer=POLY_cond $X=8.75 $Y=6.755
+ $X2=5.77 $Y2=6.755
r130 22 24 26.9307 $w=1.8e-07 $l=1.27279e-07 $layer=POLY_cond $X=5.68 $Y=6.665
+ $X2=5.77 $Y2=6.755
r131 21 22 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=5.68 $Y=5.915
+ $X2=5.68 $Y2=6.665
r132 19 21 26.9307 $w=1.8e-07 $l=1.27279e-07 $layer=POLY_cond $X=5.59 $Y=5.825
+ $X2=5.68 $Y2=5.915
r133 19 20 1206.94 $w=1.8e-07 $l=3.105e-06 $layer=POLY_cond $X=5.59 $Y=5.825
+ $X2=2.485 $Y2=5.825
r134 18 36 11.696 $w=3.4e-07 $l=2e-07 $layer=POLY_cond $X=2.395 $Y=6.125
+ $X2=2.235 $Y2=6.215
r135 17 20 26.9307 $w=1.8e-07 $l=1.27279e-07 $layer=POLY_cond $X=2.395 $Y=5.915
+ $X2=2.485 $Y2=5.825
r136 17 18 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=2.395 $Y=5.915
+ $X2=2.395 $Y2=6.125
r137 13 36 11.696 $w=3.4e-07 $l=9e-08 $layer=POLY_cond $X=2.235 $Y=6.305
+ $X2=2.235 $Y2=6.215
r138 13 15 70.6239 $w=5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.235 $Y=6.305
+ $X2=2.235 $Y2=6.965
r139 11 36 14.6411 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=1.985 $Y=6.215
+ $X2=2.235 $Y2=6.215
r140 11 12 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=1.985 $Y=6.215
+ $X2=1.705 $Y2=6.215
r141 7 12 35.539 $w=1.8e-07 $l=2.91548e-07 $layer=POLY_cond $X=1.455 $Y=6.305
+ $X2=1.705 $Y2=6.215
r142 7 9 70.6239 $w=5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.455 $Y=6.305
+ $X2=1.455 $Y2=6.965
r143 2 52 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.08
+ $Y=2.225 $X2=10.23 $Y2=3.2
r144 2 48 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.08
+ $Y=2.225 $X2=10.23 $Y2=2.37
r145 1 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.09
+ $Y=0.755 $X2=10.23 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A 1 3 6 8 9 10 14
c24 1 0 1.69832e-19 $X=10.005 $Y=2.15
r25 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.73
+ $Y=1.85 $X2=9.73 $Y2=1.85
r26 10 14 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=9.56 $Y=1.85
+ $X2=9.73 $Y2=1.85
r27 8 13 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=9.915 $Y=1.85
+ $X2=9.73 $Y2=1.85
r28 8 9 5.03009 $w=3.3e-07 $l=1.1887e-07 $layer=POLY_cond $X=9.915 $Y=1.85
+ $X2=10.005 $Y2=1.917
r29 4 9 37.0704 $w=1.5e-07 $l=2.36947e-07 $layer=POLY_cond $X=10.015 $Y=1.685
+ $X2=10.005 $Y2=1.917
r30 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.015 $Y=1.685
+ $X2=10.015 $Y2=1.125
r31 1 9 37.0704 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=10.005 $Y=2.15
+ $X2=10.005 $Y2=1.917
r32 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.005 $Y=2.15
+ $X2=10.005 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%X 1 2 9 13 19 25 27
r16 22 27 21.4773 $w=2.18e-07 $l=4.1e-07 $layer=LI1_cond $X=0.865 $Y=2.405
+ $X2=0.865 $Y2=1.995
r17 21 25 7.94788 $w=2.88e-07 $l=2e-07 $layer=LI1_cond $X=0.865 $Y=2.55
+ $X2=1.065 $Y2=2.55
r18 21 22 2.35727 $w=2.2e-07 $l=1.45e-07 $layer=LI1_cond $X=0.865 $Y=2.55
+ $X2=0.865 $Y2=2.405
r19 16 27 20.4297 $w=2.18e-07 $l=3.9e-07 $layer=LI1_cond $X=0.865 $Y=1.605
+ $X2=0.865 $Y2=1.995
r20 15 19 7.94788 $w=2.88e-07 $l=2e-07 $layer=LI1_cond $X=0.865 $Y=1.46
+ $X2=1.065 $Y2=1.46
r21 15 16 2.35727 $w=2.2e-07 $l=1.45e-07 $layer=LI1_cond $X=0.865 $Y=1.46
+ $X2=0.865 $Y2=1.605
r22 11 25 2.35727 $w=2.2e-07 $l=1.45e-07 $layer=LI1_cond $X=1.065 $Y=2.695
+ $X2=1.065 $Y2=2.55
r23 11 13 11.2625 $w=2.18e-07 $l=2.15e-07 $layer=LI1_cond $X=1.065 $Y=2.695
+ $X2=1.065 $Y2=2.91
r24 7 19 2.35727 $w=2.2e-07 $l=1.45e-07 $layer=LI1_cond $X=1.065 $Y=1.315
+ $X2=1.065 $Y2=1.46
r25 7 9 13.3579 $w=2.18e-07 $l=2.55e-07 $layer=LI1_cond $X=1.065 $Y=1.315
+ $X2=1.065 $Y2=1.06
r26 2 25 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.94
+ $Y=2.425 $X2=1.065 $Y2=2.57
r27 2 13 600 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=1 $X=0.94
+ $Y=2.425 $X2=1.065 $Y2=2.91
r28 1 19 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=0.915 $X2=1.065 $Y2=1.4
r29 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=0.915 $X2=1.065 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%VPWR 1 2 3 12 16 20 25 26
+ 29 31 32 36 39 45 53 57
c109 25 0 1.87386e-19 $X=3.535 $Y=4.41
r110 46 53 1.22274 $w=3.7e-07 $l=3.185e-06 $layer=MET1_cond $X=3.535 $Y=3.63
+ $X2=6.72 $Y2=3.63
r111 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.535 $Y=3.59
+ $X2=3.535 $Y2=3.59
r112 42 46 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=3.175 $Y=3.63
+ $X2=3.535 $Y2=3.63
r113 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.175 $Y=3.59
+ $X2=3.175 $Y2=3.59
r114 39 45 0.369424 $w=2.9e-07 $l=1.1e-07 $layer=LI1_cond $X=3.425 $Y=3.59
+ $X2=3.535 $Y2=3.59
r115 39 41 9.93485 $w=2.88e-07 $l=2.5e-07 $layer=LI1_cond $X=3.425 $Y=3.59
+ $X2=3.175 $Y2=3.59
r116 37 42 0.360871 $w=3.7e-07 $l=9.4e-07 $layer=MET1_cond $X=2.235 $Y=3.63
+ $X2=3.175 $Y2=3.63
r117 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.235 $Y=3.59
+ $X2=2.235 $Y2=3.59
r118 32 57 0.0921373 $w=3.7e-07 $l=2.4e-07 $layer=MET1_cond $X=6.96 $Y=4.51
+ $X2=6.72 $Y2=4.51
r119 31 53 0.0921373 $w=3.7e-07 $l=2.4e-07 $layer=MET1_cond $X=6.96 $Y=3.63
+ $X2=6.72 $Y2=3.63
r120 27 29 13.0959 $w=2.18e-07 $l=2.5e-07 $layer=LI1_cond $X=3.285 $Y=4.52
+ $X2=3.535 $Y2=4.52
r121 26 36 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=1.93 $Y=3.59
+ $X2=2.235 $Y2=3.59
r122 25 29 0.716491 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=3.535 $Y=4.41
+ $X2=3.535 $Y2=4.52
r123 24 45 6.45878 $w=2.2e-07 $l=1.45e-07 $layer=LI1_cond $X=3.535 $Y=3.735
+ $X2=3.535 $Y2=3.59
r124 24 25 35.359 $w=2.18e-07 $l=6.75e-07 $layer=LI1_cond $X=3.535 $Y=3.735
+ $X2=3.535 $Y2=4.41
r125 20 23 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=3.535 $Y=2.57
+ $X2=3.535 $Y2=3.25
r126 18 45 6.45878 $w=2.2e-07 $l=1.45e-07 $layer=LI1_cond $X=3.535 $Y=3.445
+ $X2=3.535 $Y2=3.59
r127 18 23 10.2148 $w=2.18e-07 $l=1.95e-07 $layer=LI1_cond $X=3.535 $Y=3.445
+ $X2=3.535 $Y2=3.25
r128 14 27 0.716491 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=3.285 $Y=4.63
+ $X2=3.285 $Y2=4.52
r129 14 16 25.1442 $w=2.18e-07 $l=4.8e-07 $layer=LI1_cond $X=3.285 $Y=4.63
+ $X2=3.285 $Y2=5.11
r130 10 26 7.43784 $w=2.9e-07 $l=1.8262e-07 $layer=LI1_cond $X=1.845 $Y=3.445
+ $X2=1.93 $Y2=3.59
r131 10 12 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.845 $Y=3.445
+ $X2=1.845 $Y2=2.57
r132 3 45 600 $w=1.7e-07 $l=1.22591e-06 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.425 $X2=3.535 $Y2=3.59
r133 3 23 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.425 $X2=3.535 $Y2=3.25
r134 3 20 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.425 $X2=3.535 $Y2=2.57
r135 2 16 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.145
+ $Y=4.965 $X2=3.285 $Y2=5.11
r136 1 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.705
+ $Y=2.425 $X2=1.845 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_188_1293# 1 2 3 4 5 18
+ 22 23 26 30 34 38 41 42 43 46 50 54 58 59 60
r96 54 57 231.536 $w=2.18e-07 $l=4.42e-06 $layer=LI1_cond $X=8.335 $Y=1.47
+ $X2=8.335 $Y2=5.89
r97 52 57 21.2154 $w=2.18e-07 $l=4.05e-07 $layer=LI1_cond $X=8.335 $Y=6.295
+ $X2=8.335 $Y2=5.89
r98 51 60 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=6.685 $Y=6.405
+ $X2=6.575 $Y2=6.405
r99 50 52 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=8.225 $Y=6.405
+ $X2=8.335 $Y2=6.295
r100 50 51 80.671 $w=2.18e-07 $l=1.54e-06 $layer=LI1_cond $X=8.225 $Y=6.405
+ $X2=6.685 $Y2=6.405
r101 46 49 231.536 $w=2.18e-07 $l=4.42e-06 $layer=LI1_cond $X=6.575 $Y=1.47
+ $X2=6.575 $Y2=5.89
r102 44 60 1.34256 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=6.575 $Y=6.295
+ $X2=6.575 $Y2=6.405
r103 44 49 21.2154 $w=2.18e-07 $l=4.05e-07 $layer=LI1_cond $X=6.575 $Y=6.295
+ $X2=6.575 $Y2=5.89
r104 42 60 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=6.465 $Y=6.405
+ $X2=6.575 $Y2=6.405
r105 42 43 81.9806 $w=2.18e-07 $l=1.565e-06 $layer=LI1_cond $X=6.465 $Y=6.405
+ $X2=4.9 $Y2=6.405
r106 40 43 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=4.79 $Y=6.515
+ $X2=4.9 $Y2=6.405
r107 40 41 58.146 $w=2.18e-07 $l=1.11e-06 $layer=LI1_cond $X=4.79 $Y=6.515
+ $X2=4.79 $Y2=7.625
r108 39 59 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.295 $Y=7.735
+ $X2=4.185 $Y2=7.735
r109 38 41 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=4.68 $Y=7.735
+ $X2=4.79 $Y2=7.625
r110 38 39 20.1678 $w=2.18e-07 $l=3.85e-07 $layer=LI1_cond $X=4.68 $Y=7.735
+ $X2=4.295 $Y2=7.735
r111 34 37 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=4.185 $Y=6.61
+ $X2=4.185 $Y2=7.29
r112 32 59 1.34256 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.185 $Y=7.625
+ $X2=4.185 $Y2=7.735
r113 32 37 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=4.185 $Y=7.625
+ $X2=4.185 $Y2=7.29
r114 31 58 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=2.735 $Y=7.735
+ $X2=2.625 $Y2=7.735
r115 30 59 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.075 $Y=7.735
+ $X2=4.185 $Y2=7.735
r116 30 31 70.1943 $w=2.18e-07 $l=1.34e-06 $layer=LI1_cond $X=4.075 $Y=7.735
+ $X2=2.735 $Y2=7.735
r117 26 29 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=2.625 $Y=6.61
+ $X2=2.625 $Y2=7.29
r118 24 58 1.34256 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=2.625 $Y=7.625
+ $X2=2.625 $Y2=7.735
r119 24 29 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=2.625 $Y=7.625
+ $X2=2.625 $Y2=7.29
r120 22 58 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=2.515 $Y=7.735
+ $X2=2.625 $Y2=7.735
r121 22 23 70.1943 $w=2.18e-07 $l=1.34e-06 $layer=LI1_cond $X=2.515 $Y=7.735
+ $X2=1.175 $Y2=7.735
r122 18 21 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=1.065 $Y=6.61
+ $X2=1.065 $Y2=7.29
r123 16 23 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=1.065 $Y=7.625
+ $X2=1.175 $Y2=7.735
r124 16 21 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=1.065 $Y=7.625
+ $X2=1.065 $Y2=7.29
r125 5 57 26 $w=1.7e-07 $l=4.63447e-06 $layer=licon1_NDIFF $count=7 $X=8.195
+ $Y=1.325 $X2=8.335 $Y2=5.89
r126 5 54 26 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=7 $X=8.195
+ $Y=1.325 $X2=8.335 $Y2=1.47
r127 4 49 26 $w=1.7e-07 $l=4.62708e-06 $layer=licon1_NDIFF $count=7 $X=6.45
+ $Y=1.325 $X2=6.575 $Y2=5.89
r128 4 46 26 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=7 $X=6.45
+ $Y=1.325 $X2=6.575 $Y2=1.47
r129 3 37 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1
+ $X=4.045 $Y=6.465 $X2=4.185 $Y2=7.29
r130 3 34 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1
+ $X=4.045 $Y=6.465 $X2=4.185 $Y2=6.61
r131 2 29 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1
+ $X=2.485 $Y=6.465 $X2=2.625 $Y2=7.29
r132 2 26 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1
+ $X=2.485 $Y=6.465 $X2=2.625 $Y2=6.61
r133 1 21 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=6.465 $X2=1.065 $Y2=7.29
r134 1 18 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=6.465 $X2=1.065 $Y2=6.61
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%VGND 1 2 3 4 5 18 20 24 30
+ 36 40 42 43 47 52 58 64 65 70 71 77 83
r86 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.18 $Y=7.635
+ $X2=10.18 $Y2=7.635
r87 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.78 $Y=0.51
+ $X2=9.78 $Y2=0.51
r88 59 65 0.825397 $w=3.7e-07 $l=2.15e-06 $layer=MET1_cond $X=7.63 $Y=0.44
+ $X2=9.78 $Y2=0.44
r89 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.63 $Y=0.51
+ $X2=7.63 $Y2=0.51
r90 55 58 8.76859 $w=2.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.455 $Y=0.51
+ $X2=7.63 $Y2=0.51
r91 53 77 1.17859 $w=3.7e-07 $l=3.07e-06 $layer=MET1_cond $X=3.65 $Y=0.44
+ $X2=6.72 $Y2=0.44
r92 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.65 $Y=0.51
+ $X2=3.65 $Y2=0.51
r93 49 52 8.76859 $w=2.28e-07 $l=1.75e-07 $layer=LI1_cond $X=3.475 $Y=0.51
+ $X2=3.65 $Y2=0.51
r94 48 53 0.681432 $w=3.7e-07 $l=1.775e-06 $layer=MET1_cond $X=1.875 $Y=0.44
+ $X2=3.65 $Y2=0.44
r95 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.875 $Y=0.51
+ $X2=1.875 $Y2=0.51
r96 43 71 1.23618 $w=3.7e-07 $l=3.22e-06 $layer=MET1_cond $X=6.96 $Y=7.7
+ $X2=10.18 $Y2=7.7
r97 43 83 0.0921373 $w=3.7e-07 $l=2.4e-07 $layer=MET1_cond $X=6.96 $Y=7.7
+ $X2=6.72 $Y2=7.7
r98 42 59 0.257217 $w=3.7e-07 $l=6.7e-07 $layer=MET1_cond $X=6.96 $Y=0.44
+ $X2=7.63 $Y2=0.44
r99 42 77 0.0921373 $w=3.7e-07 $l=2.4e-07 $layer=MET1_cond $X=6.96 $Y=0.44
+ $X2=6.72 $Y2=0.44
r100 38 70 15.5329 $w=2.28e-07 $l=3.1e-07 $layer=LI1_cond $X=9.87 $Y=7.635
+ $X2=10.18 $Y2=7.635
r101 38 40 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=9.87 $Y=7.52
+ $X2=9.87 $Y2=6.79
r102 34 64 2.50531 $w=2.28e-07 $l=5e-08 $layer=LI1_cond $X=9.73 $Y=0.51 $X2=9.78
+ $Y2=0.51
r103 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.73 $Y=0.625
+ $X2=9.73 $Y2=0.9
r104 30 32 221.469 $w=2.28e-07 $l=4.42e-06 $layer=LI1_cond $X=7.455 $Y=1.47
+ $X2=7.455 $Y2=5.89
r105 28 55 0.716491 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=7.455 $Y=0.625
+ $X2=7.455 $Y2=0.51
r106 28 30 42.3398 $w=2.28e-07 $l=8.45e-07 $layer=LI1_cond $X=7.455 $Y=0.625
+ $X2=7.455 $Y2=1.47
r107 24 26 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.475 $Y=0.81
+ $X2=3.475 $Y2=1.49
r108 22 49 0.716491 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=3.475 $Y=0.625
+ $X2=3.475 $Y2=0.51
r109 22 24 9.26965 $w=2.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.475 $Y=0.625
+ $X2=3.475 $Y2=0.81
r110 18 47 3.40825 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=1.875 $Y=0.625
+ $X2=1.875 $Y2=0.51
r111 18 20 21.7962 $w=2.28e-07 $l=4.35e-07 $layer=LI1_cond $X=1.875 $Y=0.625
+ $X2=1.875 $Y2=1.06
r112 5 40 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=9.66
+ $Y=6.645 $X2=9.87 $Y2=6.79
r113 4 36 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=9.585
+ $Y=0.755 $X2=9.73 $Y2=0.9
r114 3 32 26 $w=1.7e-07 $l=4.63447e-06 $layer=licon1_NDIFF $count=7 $X=7.315
+ $Y=1.325 $X2=7.455 $Y2=5.89
r115 3 30 26 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=7 $X=7.315
+ $Y=1.325 $X2=7.455 $Y2=1.47
r116 2 26 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1
+ $X=3.335 $Y=0.665 $X2=3.475 $Y2=1.49
r117 2 24 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1
+ $X=3.335 $Y=0.665 $X2=3.475 $Y2=0.81
r118 1 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.705
+ $Y=0.915 $X2=1.845 $Y2=1.06
.ends

