* File: sky130_fd_sc_hvl__nor2_1.pex.spice
* Created: Fri Aug 28 09:38:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__NOR2_1%VNB 5 7 11 25
r18 7 25 5.20833e-05 $w=2.4e-06 $l=1e-09 $layer=MET1_cond $X=1.2 $Y=0.057
+ $X2=1.2 $Y2=0.058
r19 7 11 0.00296875 $w=2.4e-06 $l=5.7e-08 $layer=MET1_cond $X=1.2 $Y=0.057
+ $X2=1.2 $Y2=0
r20 5 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r21 5 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR2_1%VPB 4 6 14 21
r17 10 21 0.00296875 $w=2.4e-06 $l=5.7e-08 $layer=MET1_cond $X=1.2 $Y=4.07
+ $X2=1.2 $Y2=4.013
r18 10 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=4.07
+ $X2=2.16 $Y2=4.07
r19 9 14 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=2.16 $Y2=4.07
r20 9 10 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r21 6 21 5.20833e-05 $w=2.4e-06 $l=1e-09 $layer=MET1_cond $X=1.2 $Y=4.012
+ $X2=1.2 $Y2=4.013
r22 4 14 72.8 $w=1.7e-07 $l=2.20209e-06 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=2.16 $Y2=4.07
r23 4 9 72.8 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR2_1%A 3 7 9 10 11 16
r26 16 19 19.2482 $w=5.7e-07 $l=1.95e-07 $layer=POLY_cond $X=0.97 $Y=1.89
+ $X2=0.97 $Y2=2.085
r27 16 18 45.5303 $w=5.7e-07 $l=4.75e-07 $layer=POLY_cond $X=0.97 $Y=1.89
+ $X2=0.97 $Y2=1.415
r28 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.91
+ $Y=1.89 $X2=0.91 $Y2=1.89
r29 11 17 9.6872 $w=3.43e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=1.947 $X2=0.91
+ $Y2=1.947
r30 10 17 6.34679 $w=3.43e-07 $l=1.9e-07 $layer=LI1_cond $X=0.72 $Y=1.947
+ $X2=0.91 $Y2=1.947
r31 9 10 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.947 $X2=0.72
+ $Y2=1.947
r32 7 19 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.005 $Y=2.965
+ $X2=1.005 $Y2=2.085
r33 3 18 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.935 $Y=0.91 $X2=0.935
+ $Y2=1.415
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR2_1%B 1 4 8 10
r23 7 10 115.031 $w=5e-07 $l=1.075e-06 $layer=POLY_cond $X=1.715 $Y=1.89
+ $X2=1.715 $Y2=2.965
r24 7 8 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.66 $Y=1.89
+ $X2=1.66 $Y2=1.89
r25 4 7 104.866 $w=5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.715 $Y=0.91 $X2=1.715
+ $Y2=1.89
r26 1 8 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.66 $Y=2.035
+ $X2=1.66 $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR2_1%VPWR 1 4 7 14
r17 10 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.645 $Y=3.59
+ $X2=1.645 $Y2=3.59
r18 10 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.205 $Y=3.59
+ $X2=0.205 $Y2=3.59
r19 7 10 8.80299 $w=1.668e-06 $l=1.205e-06 $layer=LI1_cond $X=0.925 $Y=2.385
+ $X2=0.925 $Y2=3.59
r20 4 14 0.170838 $w=3.7e-07 $l=4.45e-07 $layer=MET1_cond $X=1.2 $Y=3.63
+ $X2=1.645 $Y2=3.63
r21 4 11 0.381986 $w=3.7e-07 $l=9.95e-07 $layer=MET1_cond $X=1.2 $Y=3.63
+ $X2=0.205 $Y2=3.63
r22 1 10 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.47
+ $Y=2.215 $X2=0.615 $Y2=3.59
r23 1 7 300 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=2 $X=0.47
+ $Y=2.215 $X2=0.615 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR2_1%Y 1 2 9 11 12 13 14 15 16 17 24 26
r29 24 26 3.16357 $w=2.53e-07 $l=7e-08 $layer=LI1_cond $X=2.147 $Y=1.595
+ $X2=2.147 $Y2=1.665
r30 17 38 20.1113 $w=2.53e-07 $l=4.45e-07 $layer=LI1_cond $X=2.147 $Y=3.145
+ $X2=2.147 $Y2=3.59
r31 16 17 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.147 $Y=2.775
+ $X2=2.147 $Y2=3.145
r32 15 16 19.6593 $w=2.53e-07 $l=4.35e-07 $layer=LI1_cond $X=2.147 $Y=2.34
+ $X2=2.147 $Y2=2.775
r33 14 15 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=2.147 $Y=2.035
+ $X2=2.147 $Y2=2.34
r34 13 24 2.87766 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.147 $Y=1.51
+ $X2=2.147 $Y2=1.595
r35 13 14 16.4054 $w=2.53e-07 $l=3.63e-07 $layer=LI1_cond $X=2.147 $Y=1.672
+ $X2=2.147 $Y2=2.035
r36 13 26 0.316357 $w=2.53e-07 $l=7e-09 $layer=LI1_cond $X=2.147 $Y=1.672
+ $X2=2.147 $Y2=1.665
r37 11 13 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.02 $Y=1.51
+ $X2=2.147 $Y2=1.51
r38 11 12 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.02 $Y=1.51
+ $X2=1.53 $Y2=1.51
r39 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.365 $Y=1.425
+ $X2=1.53 $Y2=1.51
r40 7 9 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=1.365 $Y=1.425
+ $X2=1.365 $Y2=0.66
r41 2 38 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.965
+ $Y=2.215 $X2=2.105 $Y2=3.59
r42 2 15 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.965
+ $Y=2.215 $X2=2.105 $Y2=2.34
r43 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.185
+ $Y=0.535 $X2=1.325 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR2_1%VGND 1 2 7 10 19 20
r19 19 23 3.64905 $w=5.88e-07 $l=1.8e-07 $layer=LI1_cond $X=2.015 $Y=0.48
+ $X2=2.015 $Y2=0.66
r20 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.195 $Y=0.48
+ $X2=2.195 $Y2=0.48
r21 11 14 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.195 $Y=0.44
+ $X2=0.915 $Y2=0.44
r22 10 16 2.36129 $w=9.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.555 $Y=0.48
+ $X2=0.555 $Y2=0.66
r23 10 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.915 $Y=0.48
+ $X2=0.915 $Y2=0.48
r24 10 11 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.195 $Y=0.48
+ $X2=0.195 $Y2=0.48
r25 7 20 0.381986 $w=3.7e-07 $l=9.95e-07 $layer=MET1_cond $X=1.2 $Y=0.44
+ $X2=2.195 $Y2=0.44
r26 7 14 0.109413 $w=3.7e-07 $l=2.85e-07 $layer=MET1_cond $X=1.2 $Y=0.44
+ $X2=0.915 $Y2=0.44
r27 2 23 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.965
+ $Y=0.535 $X2=2.105 $Y2=0.66
r28 1 16 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.4
+ $Y=0.535 $X2=0.545 $Y2=0.66
.ends

