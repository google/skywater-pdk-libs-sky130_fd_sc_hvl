# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__einvn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__einvn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275000 1.725000 2.780000 2.540000 ;
        RECT 2.505000 1.160000 2.780000 1.725000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.335000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.825000 1.795000 2.025000 ;
        RECT 0.635000 2.025000 1.795000 2.120000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.950000 0.495000 3.235000 3.755000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.360000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.360000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.985000 3.360000 4.155000 ;
      RECT 0.090000  0.910000 0.440000 1.425000 ;
      RECT 0.090000  1.425000 2.065000 1.645000 ;
      RECT 0.090000  1.645000 0.345000 2.195000 ;
      RECT 0.090000  2.195000 0.455000 2.300000 ;
      RECT 0.090000  2.300000 0.535000 3.025000 ;
      RECT 0.440000  0.365000 2.770000 0.740000 ;
      RECT 0.610000  0.740000 2.770000 0.900000 ;
      RECT 0.610000  0.900000 2.335000 1.245000 ;
      RECT 0.740000  2.300000 2.105000 2.710000 ;
      RECT 0.740000  2.710000 2.770000 3.755000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.440000  0.395000 0.610000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.770000  3.505000 0.940000 3.675000 ;
      RECT 0.800000  0.395000 0.970000 0.565000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.130000  3.505000 1.300000 3.675000 ;
      RECT 1.160000  0.395000 1.330000 0.565000 ;
      RECT 1.490000  3.505000 1.660000 3.675000 ;
      RECT 1.520000  0.395000 1.690000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.850000  3.505000 2.020000 3.675000 ;
      RECT 1.880000  0.395000 2.050000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.210000  3.505000 2.380000 3.675000 ;
      RECT 2.240000  0.395000 2.410000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.570000  3.505000 2.740000 3.675000 ;
      RECT 2.600000  0.395000 2.770000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
  END
END sky130_fd_sc_hvl__einvn_1
END LIBRARY
