* File: sky130_fd_sc_hvl__einvp_1.pex.spice
* Created: Wed Sep  2 09:06:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__EINVP_1%VNB 5 7 11 25
r23 7 25 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0.058
r24 7 11 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0
r25 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r26 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVP_1%VPB 4 6 14 21
r27 10 21 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=4.07
+ $X2=1.68 $Y2=4.013
r28 10 14 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=4.07
+ $X2=3.12 $Y2=4.07
r29 9 14 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=3.12 $Y2=4.07
r30 9 10 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r31 6 21 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=4.012
+ $X2=1.68 $Y2=4.013
r32 4 14 52 $w=1.7e-07 $l=3.16221e-06 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=3.12 $Y2=4.07
r33 4 9 52 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVP_1%TE 4 7 9 10 11 13 14 15 19
r38 19 22 34.8628 $w=7.5e-07 $l=4.25e-07 $layer=POLY_cond $X=0.81 $Y=1.66
+ $X2=0.81 $Y2=2.085
r39 19 21 17.0382 $w=7.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.81 $Y=1.66
+ $X2=0.81 $Y2=1.495
r40 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.02
+ $Y=1.66 $X2=1.02 $Y2=1.66
r41 15 20 8.46693 $w=2.43e-07 $l=1.8e-07 $layer=LI1_cond $X=1.2 $Y=1.627
+ $X2=1.02 $Y2=1.627
r42 14 20 14.1115 $w=2.43e-07 $l=3e-07 $layer=LI1_cond $X=0.72 $Y=1.627 $X2=1.02
+ $Y2=1.627
r43 11 13 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.815 $Y=0.505
+ $X2=1.815 $Y2=0.99
r44 9 11 27.7928 $w=3.65e-07 $l=3.29014e-07 $layer=POLY_cond $X=1.565 $Y=0.322
+ $X2=1.815 $Y2=0.505
r45 9 10 99.5991 $w=3.65e-07 $l=6.3e-07 $layer=POLY_cond $X=1.565 $Y=0.322
+ $X2=0.935 $Y2=0.322
r46 7 22 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.935 $Y=2.59 $X2=0.935
+ $Y2=2.085
r47 4 21 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.685 $Y=1.155 $X2=0.685
+ $Y2=1.495
r48 1 10 27.7928 $w=3.65e-07 $l=3.29014e-07 $layer=POLY_cond $X=0.685 $Y=0.505
+ $X2=0.935 $Y2=0.322
r49 1 4 69.5538 $w=5e-07 $l=6.5e-07 $layer=POLY_cond $X=0.685 $Y=0.505 $X2=0.685
+ $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVP_1%A_30_189# 1 2 9 10 14 17 21 23 27 30 31 34
r49 30 34 20.7297 $w=6.7e-07 $l=2.15e-07 $layer=POLY_cond $X=1.73 $Y=1.89
+ $X2=1.73 $Y2=2.105
r50 29 31 6.09592 $w=3.73e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=1.912
+ $X2=1.475 $Y2=1.912
r51 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.56
+ $Y=1.89 $X2=1.56 $Y2=1.89
r52 23 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.9
+ $Y=1.89 $X2=1.9 $Y2=1.89
r53 21 29 3.13464 $w=3.73e-07 $l=1.02e-07 $layer=LI1_cond $X=1.662 $Y=1.912
+ $X2=1.56 $Y2=1.912
r54 21 23 7.31417 $w=3.73e-07 $l=2.38e-07 $layer=LI1_cond $X=1.662 $Y=1.912
+ $X2=1.9 $Y2=1.912
r55 20 27 3.72223 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.65 $Y=2.015
+ $X2=0.412 $Y2=2.015
r56 20 31 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.65 $Y=2.015
+ $X2=1.475 $Y2=2.015
r57 15 27 2.94878 $w=3.22e-07 $l=8.5e-08 $layer=LI1_cond $X=0.412 $Y=2.1
+ $X2=0.412 $Y2=2.015
r58 15 17 6.04334 $w=4.73e-07 $l=2.4e-07 $layer=LI1_cond $X=0.412 $Y=2.1
+ $X2=0.412 $Y2=2.34
r59 14 27 2.94878 $w=3.22e-07 $l=1.898e-07 $layer=LI1_cond $X=0.26 $Y=1.93
+ $X2=0.412 $Y2=2.015
r60 14 26 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=0.26 $Y=1.93
+ $X2=0.26 $Y2=1.335
r61 10 26 5.87448 $w=2.03e-07 $l=1.02e-07 $layer=LI1_cond $X=0.277 $Y=1.233
+ $X2=0.277 $Y2=1.335
r62 10 12 4.64195 $w=2.05e-07 $l=7.8e-08 $layer=LI1_cond $X=0.277 $Y=1.233
+ $X2=0.277 $Y2=1.155
r63 9 34 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.815 $Y=2.965 $X2=1.815
+ $Y2=2.105
r64 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.4
+ $Y=2.215 $X2=0.545 $Y2=2.34
r65 1 12 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.945 $X2=0.295 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVP_1%A 3 7 9 10 12 20 21 31
r39 29 36 0.110517 $w=3.65e-07 $l=1.65e-07 $layer=LI1_cond $X=2.627 $Y=1.955
+ $X2=2.627 $Y2=1.79
r40 29 31 2.5259 $w=3.63e-07 $l=8e-08 $layer=LI1_cond $X=2.627 $Y=1.955
+ $X2=2.627 $Y2=2.035
r41 24 36 0.110517 $w=3.65e-07 $l=1.65e-07 $layer=LI1_cond $X=2.627 $Y=1.625
+ $X2=2.627 $Y2=1.79
r42 20 23 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.61 $Y=1.79
+ $X2=2.61 $Y2=1.955
r43 20 22 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.61 $Y=1.79
+ $X2=2.61 $Y2=1.625
r44 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.78
+ $Y=1.79 $X2=2.78 $Y2=1.79
r45 10 21 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.64 $Y=1.79
+ $X2=2.78 $Y2=1.79
r46 10 36 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=2.64 $Y=1.79
+ $X2=2.627 $Y2=1.79
r47 10 12 11.6192 $w=3.63e-07 $l=3.68e-07 $layer=LI1_cond $X=2.627 $Y=2.037
+ $X2=2.627 $Y2=2.405
r48 10 31 0.0631476 $w=3.63e-07 $l=2e-09 $layer=LI1_cond $X=2.627 $Y=2.037
+ $X2=2.627 $Y2=2.035
r49 10 24 0.726197 $w=3.63e-07 $l=2.3e-08 $layer=LI1_cond $X=2.627 $Y=1.602
+ $X2=2.627 $Y2=1.625
r50 9 10 9.69315 $w=3.63e-07 $l=3.07e-07 $layer=LI1_cond $X=2.627 $Y=1.295
+ $X2=2.627 $Y2=1.602
r51 7 23 108.076 $w=5e-07 $l=1.01e-06 $layer=POLY_cond $X=2.675 $Y=2.965
+ $X2=2.675 $Y2=1.955
r52 3 22 67.9487 $w=5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.675 $Y=0.99
+ $X2=2.675 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVP_1%VPWR 1 4 11 14
r21 11 14 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.715 $Y=3.59
+ $X2=2.715 $Y2=3.59
r22 11 12 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.915 $Y=3.59
+ $X2=0.915 $Y2=3.59
r23 9 11 2.72081 $w=1.816e-06 $l=4.05e-07 $layer=LI1_cond $X=1.815 $Y=3.185
+ $X2=1.815 $Y2=3.59
r24 7 9 5.50881 $w=1.816e-06 $l=8.2e-07 $layer=LI1_cond $X=1.815 $Y=2.365
+ $X2=1.815 $Y2=3.185
r25 4 14 0.397342 $w=3.7e-07 $l=1.035e-06 $layer=MET1_cond $X=1.68 $Y=3.63
+ $X2=2.715 $Y2=3.63
r26 4 12 0.293688 $w=3.7e-07 $l=7.65e-07 $layer=MET1_cond $X=1.68 $Y=3.63
+ $X2=0.915 $Y2=3.63
r27 1 9 300 $w=1.7e-07 $l=1.08337e-06 $layer=licon1_PDIFF $count=2 $X=1.185
+ $Y=2.215 $X2=1.425 $Y2=3.185
r28 1 7 300 $w=1.7e-07 $l=3.05941e-07 $layer=licon1_PDIFF $count=2 $X=1.185
+ $Y=2.215 $X2=1.425 $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVP_1%Z 1 2 8 10 11 12 13 14 15 16 27 33
r25 25 33 1.4914 $w=2.53e-07 $l=3.3e-08 $layer=LI1_cond $X=3.107 $Y=1.328
+ $X2=3.107 $Y2=1.295
r26 16 47 20.1113 $w=2.53e-07 $l=4.45e-07 $layer=LI1_cond $X=3.107 $Y=3.145
+ $X2=3.107 $Y2=3.59
r27 15 16 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.107 $Y=2.775
+ $X2=3.107 $Y2=3.145
r28 14 15 19.6593 $w=2.53e-07 $l=4.35e-07 $layer=LI1_cond $X=3.107 $Y=2.34
+ $X2=3.107 $Y2=2.775
r29 12 13 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.135 $Y=1.665
+ $X2=3.135 $Y2=2.035
r30 12 50 11.6455 $w=1.98e-07 $l=2.1e-07 $layer=LI1_cond $X=3.135 $Y=1.665
+ $X2=3.135 $Y2=1.455
r31 11 50 5.13232 $w=2.53e-07 $l=1.01e-07 $layer=LI1_cond $X=3.107 $Y=1.354
+ $X2=3.107 $Y2=1.455
r32 11 25 1.17504 $w=2.53e-07 $l=2.6e-08 $layer=LI1_cond $X=3.107 $Y=1.354
+ $X2=3.107 $Y2=1.328
r33 11 33 1.17504 $w=2.53e-07 $l=2.6e-08 $layer=LI1_cond $X=3.107 $Y=1.269
+ $X2=3.107 $Y2=1.295
r34 10 11 15.5467 $w=2.53e-07 $l=3.44e-07 $layer=LI1_cond $X=3.107 $Y=0.925
+ $X2=3.107 $Y2=1.269
r35 10 27 8.36086 $w=2.53e-07 $l=1.85e-07 $layer=LI1_cond $X=3.107 $Y=0.925
+ $X2=3.107 $Y2=0.74
r36 9 13 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=3.135 $Y=2.125
+ $X2=3.135 $Y2=2.035
r37 8 14 3.97706 $w=2.53e-07 $l=8.8e-08 $layer=LI1_cond $X=3.107 $Y=2.252
+ $X2=3.107 $Y2=2.34
r38 8 9 6.30736 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=3.107 $Y=2.252
+ $X2=3.107 $Y2=2.125
r39 2 47 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.925
+ $Y=2.215 $X2=3.065 $Y2=3.59
r40 2 14 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.925
+ $Y=2.215 $X2=3.065 $Y2=2.34
r41 1 27 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.925
+ $Y=0.615 $X2=3.065 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HVL__EINVP_1%VGND 1 4 10 12
r28 12 14 2.41902 $w=2.093e-06 $l=4.15e-07 $layer=LI1_cond $X=1.635 $Y=0.74
+ $X2=1.635 $Y2=1.155
r29 7 12 1.51553 $w=2.093e-06 $l=2.6e-07 $layer=LI1_cond $X=1.635 $Y=0.48
+ $X2=1.635 $Y2=0.74
r30 7 10 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.715 $Y=0.48
+ $X2=2.715 $Y2=0.48
r31 7 8 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.555 $Y=0.48
+ $X2=0.555 $Y2=0.48
r32 4 10 0.397342 $w=3.7e-07 $l=1.035e-06 $layer=MET1_cond $X=1.68 $Y=0.44
+ $X2=2.715 $Y2=0.44
r33 4 8 0.431894 $w=3.7e-07 $l=1.125e-06 $layer=MET1_cond $X=1.68 $Y=0.44
+ $X2=0.555 $Y2=0.44
r34 1 14 91 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=2 $X=0.935
+ $Y=0.945 $X2=1.075 $Y2=1.155
r35 1 12 182 $w=1.7e-07 $l=5.83567e-07 $layer=licon1_NDIFF $count=1 $X=0.935
+ $Y=0.945 $X2=1.425 $Y2=0.74
.ends

