* NGSPICE file created from sky130_fd_sc_hvl__dfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__dfxtp_1 CLK D VGND VNB VPB VPWR Q
M1000 a_982_543# a_30_127# a_780_574# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=2.5915e+11p ps=2.17e+06u
M1001 a_339_559# a_30_127# VPWR VPB phv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=1.3412e+12p ps=1.246e+07u
M1002 a_1687_113# a_30_127# a_1455_543# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1003 a_1024_371# a_780_574# VPWR VPB phv w=1e+06u l=500000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1004 a_339_559# a_30_127# VGND VNB nhv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=1.09365e+12p ps=9.95e+06u
M1005 a_1015_113# a_339_559# a_780_574# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.995e+11p ps=1.79e+06u
M1006 VPWR a_1024_371# a_982_543# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_1024_371# a_1015_113# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_1729_87# a_1687_113# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Q a_1729_87# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=3.975e+11p pd=3.53e+06u as=0p ps=0u
M1010 a_1455_543# a_339_559# a_1024_371# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=2.5995e+11p ps=2.29e+06u
M1011 VPWR CLK a_30_127# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u
M1012 a_780_574# a_339_559# a_605_563# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=1.652e+11p ps=1.7e+06u
M1013 a_780_574# a_30_127# a_605_563# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.68e+11p ps=1.64e+06u
M1014 a_1731_543# a_339_559# a_1455_543# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=8.162e+11p ps=3.76e+06u
M1015 VPWR a_1729_87# a_1731_543# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_605_563# D VGND VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_605_563# D VPWR VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1729_87# a_1455_543# VPWR VPB phv w=1e+06u l=500000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1019 a_1729_87# a_1455_543# VGND VNB nhv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
M1020 a_1455_543# a_30_127# a_1024_371# VPB phv w=1e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1024_371# a_780_574# VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND CLK a_30_127# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1023 Q a_1729_87# VGND VNB nhv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
.ends

