* File: sky130_fd_sc_hvl__dfrbp_1.pex.spice
* Created: Wed Sep  2 09:04:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%VNB 5 7 11
r114 7 11 0.000424107 $w=1.68e-05 $l=5.7e-08 $layer=MET1_cond $X=8.4 $Y=0.057
+ $X2=8.4 $Y2=0
r115 5 11 0.531429 $w=1.7e-07 $l=2.975e-06 $layer=mcon $count=17 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r116 5 11 0.531429 $w=1.7e-07 $l=2.975e-06 $layer=mcon $count=17 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%VPB 4 6 14
c149 4 0 2.95049e-19 $X=-0.33 $Y=1.885
r150 10 14 0.531429 $w=1.7e-07 $l=2.975e-06 $layer=mcon $count=17 $X=16.56
+ $Y=4.07 $X2=16.56 $Y2=4.07
r151 9 14 1064.73 $w=1.68e-07 $l=1.632e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=16.56 $Y2=4.07
r152 9 10 0.531429 $w=1.7e-07 $l=2.975e-06 $layer=mcon $count=17 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r153 6 10 0.000424107 $w=1.68e-05 $l=5.7e-08 $layer=MET1_cond $X=8.4 $Y=4.013
+ $X2=8.4 $Y2=4.07
r154 4 14 10.4 $w=1.7e-07 $l=1.66024e-05 $layer=licon1_NTAP_notbjt $count=17
+ $X=0 $Y=3.985 $X2=16.56 $Y2=4.07
r155 4 9 10.4 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=17 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%CLK 1 4 10
r23 7 10 188.33 $w=5e-07 $l=1.76e-06 $layer=POLY_cond $X=0.72 $Y=1.28 $X2=0.72
+ $Y2=3.04
r24 4 7 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=0.72 $Y=0.745 $X2=0.72
+ $Y2=1.28
r25 1 7 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.76 $Y=1.28
+ $X2=0.76 $Y2=1.28
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%A_37_107# 1 2 9 13 17 22 23 24 27 30 33 35
+ 39 40 43 44 45 47 48 49 51 52 53 56 57 60 61 64 65 66 68 69 70 74 75 76 77 78
+ 79 80 81 83 90 95 98
c265 98 0 3.83042e-19 $X=10.32 $Y=0.745
c266 81 0 2.55801e-20 $X=5.522 $Y=2.96
c267 77 0 2.32009e-19 $X=9.375 $Y=1.315
c268 75 0 1.95406e-19 $X=9.29 $Y=1.985
c269 60 0 1.47443e-19 $X=5.48 $Y=3.6
c270 57 0 3.16608e-19 $X=5.485 $Y=2.715
c271 51 0 3.11168e-19 $X=3.82 $Y=3.6
c272 48 0 1.52052e-19 $X=3.735 $Y=2.735
r273 84 98 52.4329 $w=5e-07 $l=4.9e-07 $layer=POLY_cond $X=10.32 $Y=1.235
+ $X2=10.32 $Y2=0.745
r274 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.255
+ $Y=1.235 $X2=10.255 $Y2=1.235
r275 76 83 3.23493 $w=2.83e-07 $l=8e-08 $layer=LI1_cond $X=10.232 $Y=1.315
+ $X2=10.232 $Y2=1.235
r276 76 77 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=10.09 $Y=1.315
+ $X2=9.375 $Y2=1.315
r277 75 95 88.2799 $w=5e-07 $l=8.25e-07 $layer=POLY_cond $X=9.25 $Y=1.985
+ $X2=9.25 $Y2=2.81
r278 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.29
+ $Y=1.985 $X2=9.29 $Y2=1.985
r279 72 74 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=9.29 $Y=2.7
+ $X2=9.29 $Y2=1.985
r280 71 77 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.29 $Y=1.4
+ $X2=9.375 $Y2=1.315
r281 71 74 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=9.29 $Y=1.4
+ $X2=9.29 $Y2=1.985
r282 69 72 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.205 $Y=2.785
+ $X2=9.29 $Y2=2.7
r283 69 70 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=9.205 $Y=2.785
+ $X2=7.735 $Y2=2.785
r284 67 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.65 $Y=2.87
+ $X2=7.735 $Y2=2.785
r285 67 68 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=7.65 $Y=2.87
+ $X2=7.65 $Y2=3.635
r286 65 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.565 $Y=3.72
+ $X2=7.65 $Y2=3.635
r287 65 66 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.565 $Y=3.72
+ $X2=7.035 $Y2=3.72
r288 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.95 $Y=3.635
+ $X2=7.035 $Y2=3.72
r289 63 64 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.95 $Y=3.045
+ $X2=6.95 $Y2=3.635
r290 62 81 2.15711 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=5.65 $Y=2.96
+ $X2=5.522 $Y2=2.96
r291 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.865 $Y=2.96
+ $X2=6.95 $Y2=3.045
r292 61 62 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=6.865 $Y=2.96
+ $X2=5.65 $Y2=2.96
r293 59 81 4.27425 $w=2.12e-07 $l=1.03899e-07 $layer=LI1_cond $X=5.48 $Y=3.045
+ $X2=5.522 $Y2=2.96
r294 59 60 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.48 $Y=3.045
+ $X2=5.48 $Y2=3.6
r295 57 90 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=5.42 $Y=2.715
+ $X2=5.42 $Y2=3.25
r296 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.485
+ $Y=2.715 $X2=5.485 $Y2=2.715
r297 54 81 4.27425 $w=2.12e-07 $l=8.5e-08 $layer=LI1_cond $X=5.522 $Y=2.875
+ $X2=5.522 $Y2=2.96
r298 54 56 7.23101 $w=2.53e-07 $l=1.6e-07 $layer=LI1_cond $X=5.522 $Y=2.875
+ $X2=5.522 $Y2=2.715
r299 52 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.395 $Y=3.685
+ $X2=5.48 $Y2=3.6
r300 52 53 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=5.395 $Y=3.685
+ $X2=3.905 $Y2=3.685
r301 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.82 $Y=3.6
+ $X2=3.905 $Y2=3.685
r302 50 51 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.82 $Y=2.82
+ $X2=3.82 $Y2=3.6
r303 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.735 $Y=2.735
+ $X2=3.82 $Y2=2.82
r304 48 49 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.735 $Y=2.735
+ $X2=3.205 $Y2=2.735
r305 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.12 $Y=2.82
+ $X2=3.205 $Y2=2.735
r306 46 47 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.12 $Y=2.82
+ $X2=3.12 $Y2=3.635
r307 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.035 $Y=3.72
+ $X2=3.12 $Y2=3.635
r308 44 45 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=3.035 $Y=3.72
+ $X2=1.835 $Y2=3.72
r309 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.75 $Y=3.635
+ $X2=1.835 $Y2=3.72
r310 42 80 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.75 $Y=2.445
+ $X2=1.67 $Y2=2.36
r311 42 43 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=1.75 $Y=2.445
+ $X2=1.75 $Y2=3.635
r312 40 104 43.3056 $w=7.1e-07 $l=5.35e-07 $layer=POLY_cond $X=1.605 $Y=2
+ $X2=1.605 $Y2=2.535
r313 40 103 17.9591 $w=7.1e-07 $l=1.85e-07 $layer=POLY_cond $X=1.605 $Y=2
+ $X2=1.605 $Y2=1.815
r314 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.67 $Y=2
+ $X2=1.67 $Y2=2
r315 37 80 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.275
+ $X2=1.67 $Y2=2.36
r316 37 39 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.67 $Y=2.275
+ $X2=1.67 $Y2=2
r317 36 79 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.415 $Y=2.36
+ $X2=0.29 $Y2=2.36
r318 35 80 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=2.36
+ $X2=1.67 $Y2=2.36
r319 35 36 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=1.505 $Y=2.36
+ $X2=0.415 $Y2=2.36
r320 31 79 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.29 $Y=2.445
+ $X2=0.29 $Y2=2.36
r321 31 33 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=0.29 $Y=2.445
+ $X2=0.29 $Y2=2.79
r322 30 79 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.29 $Y=2.275
+ $X2=0.29 $Y2=2.36
r323 30 78 59.0051 $w=2.48e-07 $l=1.28e-06 $layer=LI1_cond $X=0.29 $Y=2.275
+ $X2=0.29 $Y2=0.995
r324 25 78 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.33 $Y=0.83
+ $X2=0.33 $Y2=0.995
r325 25 27 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.33 $Y=0.83
+ $X2=0.33 $Y2=0.745
r326 23 57 5.88532 $w=5e-07 $l=5.5e-08 $layer=POLY_cond $X=5.42 $Y=2.66 $X2=5.42
+ $Y2=2.715
r327 23 24 47.4204 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.42 $Y=2.66 $X2=5.42
+ $Y2=2.41
r328 22 24 168.339 $w=1.95e-07 $l=4.95e-07 $layer=POLY_cond $X=5.267 $Y=1.915
+ $X2=5.267 $Y2=2.41
r329 21 22 74.1719 $w=5e-07 $l=5e-07 $layer=POLY_cond $X=4.997 $Y=1.415
+ $X2=4.997 $Y2=1.915
r330 17 21 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.88 $Y=1.075 $X2=4.88
+ $Y2=1.415
r331 13 104 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.71 $Y=3.04
+ $X2=1.71 $Y2=2.535
r332 9 103 114.496 $w=5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.5 $Y=0.745 $X2=1.5
+ $Y2=1.815
r333 2 33 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.185
+ $Y=2.665 $X2=0.33 $Y2=2.79
r334 1 27 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.535 $X2=0.33 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%RESET_B 3 5 7 8 10 13 17 21 24 25 26 28 29
+ 30 31 37 39 40 41 43 44 45 46 47 51 53 56 64 67
c194 51 0 9.84974e-20 $X=11.675 $Y=1.25
c195 46 0 4.39293e-20 $X=8.43 $Y=1.21
c196 45 0 1.30913e-19 $X=11.075 $Y=1.045
c197 39 0 1.92054e-19 $X=8.43 $Y=1.825
c198 31 0 1.01253e-19 $X=8.345 $Y=1.91
c199 21 0 1.0678e-19 $X=7.265 $Y=2.645
c200 3 0 1.67177e-19 $X=3.08 $Y=3.25
r201 62 64 26.2164 $w=5e-07 $l=2.45e-07 $layer=POLY_cond $X=3.145 $Y=1.645
+ $X2=3.39 $Y2=1.645
r202 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.145
+ $Y=1.64 $X2=3.145 $Y2=1.64
r203 59 62 6.95538 $w=5e-07 $l=6.5e-08 $layer=POLY_cond $X=3.08 $Y=1.645
+ $X2=3.145 $Y2=1.645
r204 53 63 0.486211 $w=6.13e-07 $l=2.5e-08 $layer=LI1_cond $X=3.12 $Y=1.812
+ $X2=3.145 $Y2=1.812
r205 51 68 26.7574 $w=5.7e-07 $l=2.75e-07 $layer=POLY_cond $X=11.775 $Y=1.25
+ $X2=11.775 $Y2=1.525
r206 51 67 18.3095 $w=5.7e-07 $l=1.85e-07 $layer=POLY_cond $X=11.775 $Y=1.25
+ $X2=11.775 $Y2=1.065
r207 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.675
+ $Y=1.25 $X2=11.675 $Y2=1.25
r208 47 50 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=11.675 $Y=1.045
+ $X2=11.675 $Y2=1.25
r209 44 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.51 $Y=1.045
+ $X2=11.675 $Y2=1.045
r210 44 45 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=11.51 $Y=1.045
+ $X2=11.075 $Y2=1.045
r211 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.99 $Y=0.96
+ $X2=11.075 $Y2=1.045
r212 42 43 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=10.99 $Y=0.435
+ $X2=10.99 $Y2=0.96
r213 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.905 $Y=0.35
+ $X2=10.99 $Y2=0.435
r214 40 41 155.925 $w=1.68e-07 $l=2.39e-06 $layer=LI1_cond $X=10.905 $Y=0.35
+ $X2=8.515 $Y2=0.35
r215 38 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.43 $Y=1.295
+ $X2=8.43 $Y2=1.21
r216 38 39 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.43 $Y=1.295
+ $X2=8.43 $Y2=1.825
r217 37 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.43 $Y=1.125
+ $X2=8.43 $Y2=1.21
r218 36 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.43 $Y=0.435
+ $X2=8.515 $Y2=0.35
r219 36 37 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.43 $Y=0.435
+ $X2=8.43 $Y2=1.125
r220 34 56 89.3499 $w=5e-07 $l=8.35e-07 $layer=POLY_cond $X=7.265 $Y=1.91
+ $X2=7.265 $Y2=1.075
r221 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.33
+ $Y=1.91 $X2=7.33 $Y2=1.91
r222 31 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.345 $Y=1.91
+ $X2=8.43 $Y2=1.825
r223 31 33 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=8.345 $Y=1.91
+ $X2=7.33 $Y2=1.91
r224 29 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.345 $Y=1.21
+ $X2=8.43 $Y2=1.21
r225 29 30 112.214 $w=1.68e-07 $l=1.72e-06 $layer=LI1_cond $X=8.345 $Y=1.21
+ $X2=6.625 $Y2=1.21
r226 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.54 $Y=1.125
+ $X2=6.625 $Y2=1.21
r227 27 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=6.54 $Y=0.63
+ $X2=6.54 $Y2=1.125
r228 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.455 $Y=0.545
+ $X2=6.54 $Y2=0.63
r229 25 26 182.021 $w=1.68e-07 $l=2.79e-06 $layer=LI1_cond $X=6.455 $Y=0.545
+ $X2=3.665 $Y2=0.545
r230 24 63 8.46007 $w=6.13e-07 $l=4.35e-07 $layer=LI1_cond $X=3.58 $Y=1.812
+ $X2=3.145 $Y2=1.812
r231 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.58 $Y=0.63
+ $X2=3.665 $Y2=0.545
r232 23 24 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=3.58 $Y=0.63
+ $X2=3.58 $Y2=1.505
r233 21 34 78.6493 $w=5e-07 $l=7.35e-07 $layer=POLY_cond $X=7.265 $Y=2.645
+ $X2=7.265 $Y2=1.91
r234 17 67 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.81 $Y=0.745
+ $X2=11.81 $Y2=1.065
r235 13 68 106.471 $w=5e-07 $l=9.95e-07 $layer=POLY_cond $X=11.74 $Y=2.52
+ $X2=11.74 $Y2=1.525
r236 8 21 74.7205 $w=2.85e-07 $l=3.55e-07 $layer=POLY_cond $X=6.91 $Y=2.787
+ $X2=7.265 $Y2=2.787
r237 8 10 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.91 $Y=2.93 $X2=6.91
+ $Y2=3.25
r238 5 64 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.39 $Y=1.395 $X2=3.39
+ $Y2=1.645
r239 5 7 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.39 $Y=1.395 $X2=3.39
+ $Y2=1.075
r240 1 59 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.08 $Y=1.895 $X2=3.08
+ $Y2=1.645
r241 1 3 144.993 $w=5e-07 $l=1.355e-06 $layer=POLY_cond $X=3.08 $Y=1.895
+ $X2=3.08 $Y2=3.25
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%D 3 7 8 10 11 12 16
c50 11 0 1.67177e-19 $X=4.08 $Y=0.925
c51 10 0 1.18418e-19 $X=4.1 $Y=1.915
c52 8 0 1.62027e-19 $X=3.895 $Y=2.635
r53 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.015
+ $Y=1.6 $X2=4.015 $Y2=1.6
r54 16 19 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.1 $Y=1.075 $X2=4.1
+ $Y2=1.6
r55 12 20 11.1586 $w=3.13e-07 $l=3.05e-07 $layer=LI1_cond $X=4.007 $Y=1.295
+ $X2=4.007 $Y2=1.6
r56 11 12 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=4.007 $Y=0.925
+ $X2=4.007 $Y2=1.295
r57 9 19 6.95538 $w=5e-07 $l=6.5e-08 $layer=POLY_cond $X=4.1 $Y=1.665 $X2=4.1
+ $Y2=1.6
r58 9 10 32.941 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.1 $Y=1.665 $X2=4.1
+ $Y2=1.915
r59 7 8 59.6925 $w=5e-07 $l=5e-07 $layer=POLY_cond $X=3.895 $Y=2.135 $X2=3.895
+ $Y2=2.635
r60 7 10 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=4.015 $Y=2.135
+ $X2=4.015 $Y2=1.915
r61 3 8 65.8086 $w=5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.86 $Y=3.25 $X2=3.86
+ $Y2=2.635
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%A_350_107# 1 2 9 11 13 14 15 20 25 29 30 35
+ 37 39 43 45 46 47 48 51 57 58 61 69 71 72 79
c187 47 0 1.98216e-19 $X=9.695 $Y=1.665
c188 39 0 3.64387e-20 $X=5.76 $Y=1.595
c189 30 0 3.15614e-19 $X=4.78 $Y=2.315
c190 29 0 2.80445e-19 $X=4.78 $Y=2.315
c191 15 0 1.50919e-19 $X=9.5 $Y=1.492
c192 11 0 2.2109e-19 $X=9.25 $Y=1.395
c193 9 0 2.55801e-20 $X=4.64 $Y=3.25
r194 69 72 25.4802 $w=6.85e-07 $l=2.75e-07 $layer=POLY_cond $X=10.052 $Y=1.925
+ $X2=10.052 $Y2=2.2
r195 69 71 53.5705 $w=6.85e-07 $l=1.85e-07 $layer=POLY_cond $X=10.052 $Y=1.925
+ $X2=10.052 $Y2=1.74
r196 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.895
+ $Y=1.925 $X2=9.895 $Y2=1.925
r197 58 70 8.94433 $w=3.33e-07 $l=2.6e-07 $layer=LI1_cond $X=9.892 $Y=1.665
+ $X2=9.892 $Y2=1.925
r198 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=1.665
+ $X2=9.84 $Y2=1.665
r199 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.665
+ $X2=5.04 $Y2=1.665
r200 51 79 6.47738 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=2.145 $Y=1.665
+ $X2=2.145 $Y2=1.55
r201 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=1.665
r202 48 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.665
+ $X2=5.04 $Y2=1.665
r203 47 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=9.84 $Y2=1.665
r204 47 48 5.58167 $w=1.4e-07 $l=4.51e-06 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=5.185 $Y2=1.665
r205 46 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=1.665
+ $X2=2.16 $Y2=1.665
r206 45 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=5.04 $Y2=1.665
r207 45 46 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=2.305 $Y2=1.665
r208 43 55 23.2584 $w=2.73e-07 $l=5.55e-07 $layer=LI1_cond $X=5.595 $Y=1.642
+ $X2=5.04 $Y2=1.642
r209 42 43 1.82517 $w=2.75e-07 $l=1.65e-07 $layer=LI1_cond $X=5.76 $Y=1.642
+ $X2=5.595 $Y2=1.642
r210 40 61 55.6431 $w=5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.825 $Y=1.595
+ $X2=5.825 $Y2=1.075
r211 39 42 1.64136 $w=3.28e-07 $l=4.7e-08 $layer=LI1_cond $X=5.76 $Y=1.595
+ $X2=5.76 $Y2=1.642
r212 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.76
+ $Y=1.595 $X2=5.76 $Y2=1.595
r213 37 55 7.33373 $w=2.73e-07 $l=1.75e-07 $layer=LI1_cond $X=4.865 $Y=1.642
+ $X2=5.04 $Y2=1.642
r214 33 35 5.02353 $w=4.98e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=0.745
+ $X2=2.1 $Y2=0.745
r215 30 67 56.7941 $w=5.7e-07 $l=5.95e-07 $layer=POLY_cond $X=4.675 $Y=2.315
+ $X2=4.675 $Y2=2.91
r216 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.78
+ $Y=2.315 $X2=4.78 $Y2=2.315
r217 27 37 7.32204 $w=2.75e-07 $l=1.75425e-07 $layer=LI1_cond $X=4.78 $Y=1.78
+ $X2=4.865 $Y2=1.642
r218 27 29 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=4.78 $Y=1.78
+ $X2=4.78 $Y2=2.315
r219 23 51 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=2.145 $Y=1.68
+ $X2=2.145 $Y2=1.665
r220 23 25 49.2005 $w=2.58e-07 $l=1.11e-06 $layer=LI1_cond $X=2.145 $Y=1.68
+ $X2=2.145 $Y2=2.79
r221 21 35 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=2.1 $Y=0.995 $X2=2.1
+ $Y2=0.745
r222 21 79 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.1 $Y=0.995
+ $X2=2.1 $Y2=1.55
r223 20 72 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.145 $Y=2.52
+ $X2=10.145 $Y2=2.2
r224 16 71 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=9.785 $Y=1.59
+ $X2=9.785 $Y2=1.74
r225 14 16 27.531 $w=1.95e-07 $l=1.30208e-07 $layer=POLY_cond $X=9.71 $Y=1.492
+ $X2=9.785 $Y2=1.59
r226 14 15 71.4166 $w=1.95e-07 $l=2.1e-07 $layer=POLY_cond $X=9.71 $Y=1.492
+ $X2=9.5 $Y2=1.492
r227 11 15 34.3048 $w=1.95e-07 $l=2.94534e-07 $layer=POLY_cond $X=9.25 $Y=1.395
+ $X2=9.5 $Y2=1.492
r228 11 13 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.25 $Y=1.395
+ $X2=9.25 $Y2=0.91
r229 9 67 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.64 $Y=3.25 $X2=4.64
+ $Y2=2.91
r230 2 25 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=2.665 $X2=2.1 $Y2=2.79
r231 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.535 $X2=1.89 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%A_1176_466# 1 2 7 9 13 18 22 23 25 26 29 31
c90 26 0 1.0678e-19 $X=6.785 $Y=2.26
c91 25 0 7.92603e-20 $X=8.695 $Y=2.26
c92 9 0 5.91168e-20 $X=6.13 $Y=3.25
c93 7 0 2.28267e-19 $X=6.13 $Y=2.91
r94 31 33 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=8.86 $Y=2.26
+ $X2=8.86 $Y2=2.435
r95 27 31 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.86 $Y=2.175
+ $X2=8.86 $Y2=2.26
r96 27 29 51.5107 $w=3.28e-07 $l=1.475e-06 $layer=LI1_cond $X=8.86 $Y=2.175
+ $X2=8.86 $Y2=0.7
r97 25 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=2.26
+ $X2=8.86 $Y2=2.26
r98 25 26 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=8.695 $Y=2.26
+ $X2=6.785 $Y2=2.26
r99 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.62
+ $Y=1.91 $X2=6.62 $Y2=1.91
r100 20 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.62 $Y=2.175
+ $X2=6.785 $Y2=2.26
r101 20 22 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=6.62 $Y=2.175
+ $X2=6.62 $Y2=1.91
r102 18 23 24.1792 $w=5.2e-07 $l=2.35e-07 $layer=POLY_cond $X=6.545 $Y=1.675
+ $X2=6.545 $Y2=1.91
r103 18 19 26.7515 $w=5.2e-07 $l=2.6e-07 $layer=POLY_cond $X=6.545 $Y=1.675
+ $X2=6.545 $Y2=1.415
r104 17 23 43.2139 $w=5.2e-07 $l=4.2e-07 $layer=POLY_cond $X=6.545 $Y=2.33
+ $X2=6.545 $Y2=1.91
r105 13 19 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.535 $Y=1.075
+ $X2=6.535 $Y2=1.415
r106 7 17 50.3854 $w=3.97e-07 $l=5.40902e-07 $layer=POLY_cond $X=6.13 $Y=2.62
+ $X2=6.545 $Y2=2.33
r107 7 9 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.13 $Y=2.91 $X2=6.13
+ $Y2=3.25
r108 2 33 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=8.72
+ $Y=2.31 $X2=8.86 $Y2=2.435
r109 1 29 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=8.72
+ $Y=0.535 $X2=8.86 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%A_978_608# 1 2 3 10 12 15 19 20 21 24 26 28
+ 31 34 35 38 41 42 45 49 50 53
c144 41 0 5.91168e-20 $X=5.03 $Y=3.25
c145 31 0 1.91828e-19 $X=8 $Y=1.56
c146 20 0 1.98216e-19 $X=5.215 $Y=2.285
c147 10 0 8.109e-20 $X=8.47 $Y=1.395
r148 45 47 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=1.075
+ $X2=5.435 $Y2=1.24
r149 41 42 11.2873 $w=3.48e-07 $l=2.5e-07 $layer=LI1_cond $X=5.04 $Y=3.25
+ $X2=5.04 $Y2=3
r150 36 38 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.3 $Y=2.695
+ $X2=7.3 $Y2=3.225
r151 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.215 $Y=2.61
+ $X2=7.3 $Y2=2.695
r152 34 35 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=7.215 $Y=2.61
+ $X2=6.275 $Y2=2.61
r153 32 53 50.2928 $w=5e-07 $l=4.7e-07 $layer=POLY_cond $X=8 $Y=1.645 $X2=8.47
+ $Y2=1.645
r154 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8 $Y=1.56
+ $X2=8 $Y2=1.56
r155 29 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.275 $Y=1.56
+ $X2=6.19 $Y2=1.56
r156 29 31 112.54 $w=1.68e-07 $l=1.725e-06 $layer=LI1_cond $X=6.275 $Y=1.56
+ $X2=8 $Y2=1.56
r157 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.19 $Y=2.525
+ $X2=6.275 $Y2=2.61
r158 27 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.19 $Y=2.37
+ $X2=6.19 $Y2=2.285
r159 27 28 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.19 $Y=2.37
+ $X2=6.19 $Y2=2.525
r160 26 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.19 $Y=2.2 $X2=6.19
+ $Y2=2.285
r161 25 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.19 $Y=1.645
+ $X2=6.19 $Y2=1.56
r162 25 26 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=6.19 $Y=1.645
+ $X2=6.19 $Y2=2.2
r163 24 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.19 $Y=1.475
+ $X2=6.19 $Y2=1.56
r164 23 24 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.19 $Y=1.325
+ $X2=6.19 $Y2=1.475
r165 22 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.6 $Y=1.24
+ $X2=5.435 $Y2=1.24
r166 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.105 $Y=1.24
+ $X2=6.19 $Y2=1.325
r167 21 22 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=6.105 $Y=1.24
+ $X2=5.6 $Y2=1.24
r168 19 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.105 $Y=2.285
+ $X2=6.19 $Y2=2.285
r169 19 20 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=6.105 $Y=2.285
+ $X2=5.215 $Y2=2.285
r170 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.13 $Y=2.37
+ $X2=5.215 $Y2=2.285
r171 17 42 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.13 $Y=2.37
+ $X2=5.13 $Y2=3
r172 13 53 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.47 $Y=1.895
+ $X2=8.47 $Y2=1.645
r173 13 15 97.9104 $w=5e-07 $l=9.15e-07 $layer=POLY_cond $X=8.47 $Y=1.895
+ $X2=8.47 $Y2=2.81
r174 10 53 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.47 $Y=1.395
+ $X2=8.47 $Y2=1.645
r175 10 12 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=8.47 $Y=1.395
+ $X2=8.47 $Y2=0.91
r176 3 38 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=7.16
+ $Y=3.04 $X2=7.3 $Y2=3.225
r177 2 41 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=3.04 $X2=5.03 $Y2=3.25
r178 1 45 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=5.13
+ $Y=0.865 $X2=5.435 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%A_2122_348# 1 2 9 12 13 15 18 20 22 27 33
+ 36 38
c76 22 0 1.68113e-19 $X=11.095 $Y=1.395
r77 33 35 10.5766 $w=3.63e-07 $l=2.3e-07 $layer=LI1_cond $X=12.892 $Y=0.745
+ $X2=12.892 $Y2=0.975
r78 27 30 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=12.13 $Y=2.435
+ $X2=12.13 $Y2=2.52
r79 23 38 69.5538 $w=5e-07 $l=6.5e-07 $layer=POLY_cond $X=11.03 $Y=1.395
+ $X2=11.03 $Y2=0.745
r80 22 25 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=11.095 $Y=1.395
+ $X2=11.095 $Y2=1.615
r81 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.095
+ $Y=1.395 $X2=11.095 $Y2=1.395
r82 19 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.795 $Y=1.7
+ $X2=12.795 $Y2=1.615
r83 19 20 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=12.795 $Y=1.7
+ $X2=12.795 $Y2=2.35
r84 18 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.795 $Y=1.53
+ $X2=12.795 $Y2=1.615
r85 18 35 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=12.795 $Y=1.53
+ $X2=12.795 $Y2=0.975
r86 16 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.295 $Y=2.435
+ $X2=12.13 $Y2=2.435
r87 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.71 $Y=2.435
+ $X2=12.795 $Y2=2.35
r88 15 16 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=12.71 $Y=2.435
+ $X2=12.295 $Y2=2.435
r89 14 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.26 $Y=1.615
+ $X2=11.095 $Y2=1.615
r90 13 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.71 $Y=1.615
+ $X2=12.795 $Y2=1.615
r91 13 14 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=12.71 $Y=1.615
+ $X2=11.26 $Y2=1.615
r92 11 23 36.917 $w=5e-07 $l=3.45e-07 $layer=POLY_cond $X=11.03 $Y=1.74
+ $X2=11.03 $Y2=1.395
r93 11 12 36.7334 $w=6.7e-07 $l=4.6e-07 $layer=POLY_cond $X=10.945 $Y=1.74
+ $X2=10.945 $Y2=2.2
r94 9 12 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.86 $Y=2.52 $X2=10.86
+ $Y2=2.2
r95 2 30 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.99
+ $Y=2.31 $X2=12.13 $Y2=2.52
r96 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.77
+ $Y=0.535 $X2=12.91 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%A_1900_107# 1 2 9 11 13 14 18 22 24 28 32
+ 34 35 36 38 40 42 45 46 47 53 56 57
r151 56 59 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=12.365 $Y=1.985
+ $X2=12.365 $Y2=2.085
r152 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.365
+ $Y=1.985 $X2=12.365 $Y2=1.985
r153 51 53 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=9.745 $Y=0.805
+ $X2=9.91 $Y2=0.805
r154 47 54 5.47079 $w=2.64e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.725 $Y=2.085
+ $X2=10.64 $Y2=2.17
r155 46 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.2 $Y=2.085
+ $X2=12.365 $Y2=2.085
r156 46 47 96.2299 $w=1.68e-07 $l=1.475e-06 $layer=LI1_cond $X=12.2 $Y=2.085
+ $X2=10.725 $Y2=2.085
r157 45 54 3.3128 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=10.64 $Y=2 $X2=10.64
+ $Y2=2.17
r158 44 45 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=10.64 $Y=0.785
+ $X2=10.64 $Y2=2
r159 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.555 $Y=0.7
+ $X2=10.64 $Y2=0.785
r160 42 53 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=10.555 $Y=0.7
+ $X2=9.91 $Y2=0.7
r161 41 49 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.805 $Y=2.355
+ $X2=9.68 $Y2=2.355
r162 40 54 20.0276 $w=2.64e-07 $l=4.83735e-07 $layer=LI1_cond $X=10.24 $Y=2.355
+ $X2=10.64 $Y2=2.17
r163 40 41 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=10.24 $Y=2.355
+ $X2=9.805 $Y2=2.355
r164 36 49 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.68 $Y=2.44
+ $X2=9.68 $Y2=2.355
r165 36 38 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=9.68 $Y=2.44
+ $X2=9.68 $Y2=2.81
r166 30 35 20.4101 $w=5e-07 $l=3.39963e-07 $layer=POLY_cond $X=15.24 $Y=1.415
+ $X2=15.23 $Y2=1.75
r167 30 32 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=15.24 $Y=1.415
+ $X2=15.24 $Y2=1.075
r168 26 35 20.4101 $w=5e-07 $l=3.39963e-07 $layer=POLY_cond $X=15.22 $Y=2.085
+ $X2=15.23 $Y2=1.75
r169 26 28 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=15.22 $Y=2.085
+ $X2=15.22 $Y2=2.59
r170 25 34 12.05 $w=5e-07 $l=2.73e-07 $layer=POLY_cond $X=14.12 $Y=1.835
+ $X2=13.847 $Y2=1.835
r171 24 35 5.30422 $w=5e-07 $l=2.995e-07 $layer=POLY_cond $X=14.97 $Y=1.835
+ $X2=15.23 $Y2=1.75
r172 24 25 90.955 $w=5e-07 $l=8.5e-07 $layer=POLY_cond $X=14.97 $Y=1.835
+ $X2=14.12 $Y2=1.835
r173 20 34 12.05 $w=5e-07 $l=2.61247e-07 $layer=POLY_cond $X=13.87 $Y=1.585
+ $X2=13.847 $Y2=1.835
r174 20 22 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=13.87 $Y=1.585
+ $X2=13.87 $Y2=1.08
r175 16 34 12.05 $w=5e-07 $l=2.60768e-07 $layer=POLY_cond $X=13.825 $Y=2.085
+ $X2=13.847 $Y2=1.835
r176 16 18 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=13.825 $Y=2.085
+ $X2=13.825 $Y2=2.965
r177 15 57 5.30422 $w=5e-07 $l=6.17981e-07 $layer=POLY_cond $X=12.77 $Y=1.835
+ $X2=12.2 $Y2=1.735
r178 14 34 12.05 $w=5e-07 $l=2.72e-07 $layer=POLY_cond $X=13.575 $Y=1.835
+ $X2=13.847 $Y2=1.835
r179 14 15 86.1397 $w=5e-07 $l=8.05e-07 $layer=POLY_cond $X=13.575 $Y=1.835
+ $X2=12.77 $Y2=1.835
r180 11 57 20.4101 $w=5e-07 $l=6.04173e-07 $layer=POLY_cond $X=12.52 $Y=2.2
+ $X2=12.2 $Y2=1.735
r181 11 13 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=12.52 $Y=2.2 $X2=12.52
+ $Y2=2.52
r182 7 57 20.4101 $w=5e-07 $l=3.87814e-07 $layer=POLY_cond $X=12.52 $Y=1.585
+ $X2=12.2 $Y2=1.735
r183 7 9 89.8849 $w=5e-07 $l=8.4e-07 $layer=POLY_cond $X=12.52 $Y=1.585
+ $X2=12.52 $Y2=0.745
r184 2 49 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=9.5
+ $Y=2.31 $X2=9.64 $Y2=2.435
r185 2 38 300 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_PDIFF $count=2 $X=9.5
+ $Y=2.31 $X2=9.64 $Y2=2.81
r186 1 51 182 $w=1.7e-07 $l=3.41138e-07 $layer=licon1_NDIFF $count=1 $X=9.5
+ $Y=0.535 $X2=9.745 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%A_2937_443# 1 2 9 13 17 21 25 26 28
r46 26 31 23.8503 $w=5.75e-07 $l=2.45e-07 $layer=POLY_cond $X=16.097 $Y=1.67
+ $X2=16.097 $Y2=1.915
r47 26 30 24.7808 $w=5.75e-07 $l=2.55e-07 $layer=POLY_cond $X=16.097 $Y=1.67
+ $X2=16.097 $Y2=1.415
r48 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.995
+ $Y=1.67 $X2=15.995 $Y2=1.67
r49 23 28 1.45028 $w=3.3e-07 $l=1.75e-07 $layer=LI1_cond $X=15.015 $Y=1.67
+ $X2=14.84 $Y2=1.67
r50 23 25 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=15.015 $Y=1.67
+ $X2=15.995 $Y2=1.67
r51 19 28 5.0389 $w=3.4e-07 $l=1.69926e-07 $layer=LI1_cond $X=14.83 $Y=1.835
+ $X2=14.84 $Y2=1.67
r52 19 21 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=14.83 $Y=1.835
+ $X2=14.83 $Y2=2.34
r53 15 28 5.0389 $w=3.4e-07 $l=1.65e-07 $layer=LI1_cond $X=14.84 $Y=1.505
+ $X2=14.84 $Y2=1.67
r54 15 17 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=14.84 $Y=1.505
+ $X2=14.84 $Y2=1.075
r55 13 30 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=16.135 $Y=0.91
+ $X2=16.135 $Y2=1.415
r56 9 31 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=16.115 $Y=2.965
+ $X2=16.115 $Y2=1.915
r57 2 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=14.685
+ $Y=2.215 $X2=14.83 $Y2=2.34
r58 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=14.705
+ $Y=0.865 $X2=14.85 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%VPWR 1 2 3 4 5 6 7 22 25 34 47 51 60 69 81
+ 89
r126 87 89 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=15.29 $Y=3.63
+ $X2=16.01 $Y2=3.63
r127 86 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.01 $Y=3.59
+ $X2=16.01 $Y2=3.59
r128 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.29 $Y=3.59
+ $X2=15.29 $Y2=3.59
r129 84 86 5.32947 $w=9.48e-07 $l=4.15e-07 $layer=LI1_cond $X=15.65 $Y=3.175
+ $X2=15.65 $Y2=3.59
r130 81 84 10.7232 $w=9.48e-07 $l=8.35e-07 $layer=LI1_cond $X=15.65 $Y=2.34
+ $X2=15.65 $Y2=3.175
r131 78 87 0.547065 $w=3.7e-07 $l=1.425e-06 $layer=MET1_cond $X=13.865 $Y=3.63
+ $X2=15.29 $Y2=3.63
r132 75 78 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=13.145 $Y=3.63
+ $X2=13.865 $Y2=3.63
r133 74 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.865 $Y=3.59
+ $X2=13.865 $Y2=3.59
r134 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.145 $Y=3.59
+ $X2=13.145 $Y2=3.59
r135 72 74 11.4461 $w=8.88e-07 $l=8.35e-07 $layer=LI1_cond $X=13.505 $Y=2.755
+ $X2=13.505 $Y2=3.59
r136 69 72 5.68876 $w=8.88e-07 $l=4.15e-07 $layer=LI1_cond $X=13.505 $Y=2.34
+ $X2=13.505 $Y2=2.755
r137 66 75 0.660317 $w=3.7e-07 $l=1.72e-06 $layer=MET1_cond $X=11.425 $Y=3.63
+ $X2=13.145 $Y2=3.63
r138 64 66 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.705 $Y=3.63
+ $X2=11.425 $Y2=3.63
r139 63 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.425 $Y=3.59
+ $X2=11.425 $Y2=3.59
r140 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.705 $Y=3.59
+ $X2=10.705 $Y2=3.59
r141 60 63 13.7411 $w=9.48e-07 $l=1.07e-06 $layer=LI1_cond $X=11.065 $Y=2.52
+ $X2=11.065 $Y2=3.59
r142 57 64 0.750535 $w=3.7e-07 $l=1.955e-06 $layer=MET1_cond $X=8.75 $Y=3.63
+ $X2=10.705 $Y2=3.63
r143 54 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.75 $Y=3.59
+ $X2=8.75 $Y2=3.59
r144 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.03 $Y=3.59
+ $X2=8.03 $Y2=3.59
r145 51 54 5.52211 $w=9.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.39 $Y=3.16
+ $X2=8.39 $Y2=3.59
r146 48 55 0.558582 $w=3.7e-07 $l=1.455e-06 $layer=MET1_cond $X=6.575 $Y=3.63
+ $X2=8.03 $Y2=3.63
r147 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.575 $Y=3.59
+ $X2=6.575 $Y2=3.59
r148 45 47 1.37051 $w=4.78e-07 $l=5.5e-08 $layer=LI1_cond $X=6.52 $Y=3.465
+ $X2=6.575 $Y2=3.465
r149 42 48 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.855 $Y=3.63
+ $X2=6.575 $Y2=3.63
r150 41 45 16.5707 $w=4.78e-07 $l=6.65e-07 $layer=LI1_cond $X=5.855 $Y=3.465
+ $X2=6.52 $Y2=3.465
r151 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.855 $Y=3.59
+ $X2=5.855 $Y2=3.59
r152 38 42 0.915614 $w=3.7e-07 $l=2.385e-06 $layer=MET1_cond $X=3.47 $Y=3.63
+ $X2=5.855 $Y2=3.63
r153 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.47 $Y=3.59
+ $X2=3.47 $Y2=3.59
r154 34 37 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.47 $Y=3.25
+ $X2=3.47 $Y2=3.59
r155 31 38 0.794684 $w=3.7e-07 $l=2.07e-06 $layer=MET1_cond $X=1.4 $Y=3.63
+ $X2=3.47 $Y2=3.63
r156 29 31 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.68 $Y=3.63
+ $X2=1.4 $Y2=3.63
r157 28 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.4 $Y=3.59
+ $X2=1.4 $Y2=3.59
r158 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.68 $Y=3.59
+ $X2=0.68 $Y2=3.59
r159 25 28 10.9663 $w=8.88e-07 $l=8e-07 $layer=LI1_cond $X=1.04 $Y=2.79 $X2=1.04
+ $Y2=3.59
r160 22 57 0.134367 $w=3.7e-07 $l=3.5e-07 $layer=MET1_cond $X=8.4 $Y=3.63
+ $X2=8.75 $Y2=3.63
r161 22 55 0.142045 $w=3.7e-07 $l=3.7e-07 $layer=MET1_cond $X=8.4 $Y=3.63
+ $X2=8.03 $Y2=3.63
r162 7 84 300 $w=1.7e-07 $l=1.08e-06 $layer=licon1_PDIFF $count=2 $X=15.47
+ $Y=2.215 $X2=15.725 $Y2=3.175
r163 7 81 300 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=2 $X=15.47
+ $Y=2.215 $X2=15.725 $Y2=2.34
r164 6 74 400 $w=1.7e-07 $l=1.57785e-06 $layer=licon1_PDIFF $count=1 $X=12.77
+ $Y=2.31 $X2=13.435 $Y2=3.59
r165 6 72 400 $w=1.7e-07 $l=8.59157e-07 $layer=licon1_PDIFF $count=1 $X=12.77
+ $Y=2.31 $X2=13.435 $Y2=2.755
r166 6 69 600 $w=1.7e-07 $l=6.79835e-07 $layer=licon1_PDIFF $count=1 $X=12.77
+ $Y=2.31 $X2=13.435 $Y2=2.34
r167 5 60 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.11
+ $Y=2.31 $X2=11.25 $Y2=2.52
r168 4 51 600 $w=1.7e-07 $l=9.19647e-07 $layer=licon1_PDIFF $count=1 $X=7.935
+ $Y=2.31 $X2=8.08 $Y2=3.16
r169 3 45 600 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=3.04 $X2=6.52 $Y2=3.32
r170 2 34 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.33
+ $Y=3.04 $X2=3.47 $Y2=3.25
r171 1 25 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.97
+ $Y=2.665 $X2=1.11 $Y2=2.79
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%A_509_608# 1 2 3 12 14 15 18 21 23 27 29 30
c64 27 0 1.38804e-19 $X=4.43 $Y=3.21
c65 23 0 1.77803e-19 $X=4.43 $Y=3
r66 25 27 4.93904 $w=4.18e-07 $l=1.8e-07 $layer=LI1_cond $X=4.25 $Y=3.21
+ $X2=4.43 $Y2=3.21
r67 23 27 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=4.43 $Y=3 $X2=4.43
+ $Y2=3.21
r68 22 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.43 $Y=2.47 $X2=4.43
+ $Y2=2.385
r69 22 23 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.43 $Y=2.47
+ $X2=4.43 $Y2=3
r70 21 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.43 $Y=2.3 $X2=4.43
+ $Y2=2.385
r71 21 29 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=4.43 $Y=2.3
+ $X2=4.43 $Y2=1.325
r72 16 29 8.09553 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=4.5 $Y=1.17 $X2=4.5
+ $Y2=1.325
r73 16 18 3.53168 $w=3.08e-07 $l=9.5e-08 $layer=LI1_cond $X=4.5 $Y=1.17 $X2=4.5
+ $Y2=1.075
r74 14 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.345 $Y=2.385
+ $X2=4.43 $Y2=2.385
r75 14 15 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=4.345 $Y=2.385
+ $X2=2.855 $Y2=2.385
r76 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.69 $Y=2.47
+ $X2=2.855 $Y2=2.385
r77 10 12 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=2.69 $Y=2.47
+ $X2=2.69 $Y2=3.25
r78 3 25 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.11
+ $Y=3.04 $X2=4.25 $Y2=3.25
r79 2 12 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=2.545
+ $Y=3.04 $X2=2.69 $Y2=3.25
r80 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.35
+ $Y=0.865 $X2=4.49 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%Q_N 1 2 7 9 13 14 15 22 28
r26 20 28 0.303274 $w=3.78e-07 $l=1e-08 $layer=LI1_cond $X=14.235 $Y=1.305
+ $X2=14.235 $Y2=1.295
r27 14 15 11.1632 $w=3.53e-07 $l=3.23e-07 $layer=LI1_cond $X=14.235 $Y=1.342
+ $X2=14.235 $Y2=1.665
r28 14 20 1.26811 $w=3.8e-07 $l=3.7e-08 $layer=LI1_cond $X=14.235 $Y=1.342
+ $X2=14.235 $Y2=1.305
r29 14 28 1.15244 $w=3.78e-07 $l=3.8e-08 $layer=LI1_cond $X=14.235 $Y=1.257
+ $X2=14.235 $Y2=1.295
r30 13 14 10.0687 $w=3.78e-07 $l=3.32e-07 $layer=LI1_cond $X=14.235 $Y=0.925
+ $X2=14.235 $Y2=1.257
r31 13 22 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=14.235 $Y=0.925
+ $X2=14.235 $Y2=0.83
r32 9 11 57.6222 $w=2.48e-07 $l=1.25e-06 $layer=LI1_cond $X=14.255 $Y=2.34
+ $X2=14.255 $Y2=3.59
r33 7 15 5.02948 $w=3.53e-07 $l=1.24599e-07 $layer=LI1_cond $X=14.255 $Y=1.78
+ $X2=14.235 $Y2=1.665
r34 7 9 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=14.255 $Y=1.78
+ $X2=14.255 $Y2=2.34
r35 2 11 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=14.075
+ $Y=2.215 $X2=14.215 $Y2=3.59
r36 2 9 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=14.075
+ $Y=2.215 $X2=14.215 $Y2=2.34
r37 1 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=14.12
+ $Y=0.705 $X2=14.26 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%Q 1 2 7 8 9 10 11 12 13 22
r13 13 40 14.6525 $w=3.48e-07 $l=4.45e-07 $layer=LI1_cond $X=16.515 $Y=3.145
+ $X2=16.515 $Y2=3.59
r14 12 13 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=16.515 $Y=2.775
+ $X2=16.515 $Y2=3.145
r15 11 12 14.3232 $w=3.48e-07 $l=4.35e-07 $layer=LI1_cond $X=16.515 $Y=2.34
+ $X2=16.515 $Y2=2.775
r16 10 11 10.0427 $w=3.48e-07 $l=3.05e-07 $layer=LI1_cond $X=16.515 $Y=2.035
+ $X2=16.515 $Y2=2.34
r17 9 10 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=16.515 $Y=1.665
+ $X2=16.515 $Y2=2.035
r18 8 9 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=16.515 $Y=1.295
+ $X2=16.515 $Y2=1.665
r19 7 8 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=16.515 $Y=0.925
+ $X2=16.515 $Y2=1.295
r20 7 22 8.0671 $w=3.48e-07 $l=2.45e-07 $layer=LI1_cond $X=16.515 $Y=0.925
+ $X2=16.515 $Y2=0.68
r21 2 40 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=16.365
+ $Y=2.215 $X2=16.505 $Y2=3.59
r22 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=16.365
+ $Y=2.215 $X2=16.505 $Y2=2.34
r23 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=16.385
+ $Y=0.535 $X2=16.525 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRBP_1%VGND 1 2 3 4 5 6 19 22 31 46 56 60 67 71
c103 56 0 1.82514e-19 $X=12.09 $Y=0.48
r104 73 75 6.42105 $w=9.48e-07 $l=5e-07 $layer=LI1_cond $X=15.67 $Y=0.66
+ $X2=15.67 $Y2=1.16
r105 68 71 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=15.31 $Y=0.44
+ $X2=16.03 $Y2=0.44
r106 67 73 2.31158 $w=9.48e-07 $l=1.8e-07 $layer=LI1_cond $X=15.67 $Y=0.48
+ $X2=15.67 $Y2=0.66
r107 67 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.03 $Y=0.48
+ $X2=16.03 $Y2=0.48
r108 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.31 $Y=0.48
+ $X2=15.31 $Y2=0.48
r109 61 68 0.606571 $w=3.7e-07 $l=1.58e-06 $layer=MET1_cond $X=13.73 $Y=0.44
+ $X2=15.31 $Y2=0.44
r110 60 64 7.09538 $w=5.88e-07 $l=3.5e-07 $layer=LI1_cond $X=13.55 $Y=0.48
+ $X2=13.55 $Y2=0.83
r111 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.73 $Y=0.48
+ $X2=13.73 $Y2=0.48
r112 57 61 0.629605 $w=3.7e-07 $l=1.64e-06 $layer=MET1_cond $X=12.09 $Y=0.44
+ $X2=13.73 $Y2=0.44
r113 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.09 $Y=0.48
+ $X2=12.09 $Y2=0.48
r114 54 56 18.6057 $w=4.13e-07 $l=6.7e-07 $layer=LI1_cond $X=11.42 $Y=0.572
+ $X2=12.09 $Y2=0.572
r115 51 57 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=11.37 $Y=0.44
+ $X2=12.09 $Y2=0.44
r116 50 54 1.38849 $w=4.13e-07 $l=5e-08 $layer=LI1_cond $X=11.37 $Y=0.572
+ $X2=11.42 $Y2=0.572
r117 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.37 $Y=0.48
+ $X2=11.37 $Y2=0.48
r118 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=0.48
+ $X2=8.05 $Y2=0.48
r119 44 46 1.0311 $w=5.78e-07 $l=5e-08 $layer=LI1_cond $X=8 $Y=0.655 $X2=8.05
+ $Y2=0.655
r120 41 47 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.33 $Y=0.44
+ $X2=8.05 $Y2=0.44
r121 40 44 13.8168 $w=5.78e-07 $l=6.7e-07 $layer=LI1_cond $X=7.33 $Y=0.655 $X2=8
+ $Y2=0.655
r122 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.33 $Y=0.48
+ $X2=7.33 $Y2=0.48
r123 35 41 1.58553 $w=3.7e-07 $l=4.13e-06 $layer=MET1_cond $X=3.2 $Y=0.44
+ $X2=7.33 $Y2=0.44
r124 32 35 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.48 $Y=0.44
+ $X2=3.2 $Y2=0.44
r125 31 37 7.64105 $w=9.48e-07 $l=5.95e-07 $layer=LI1_cond $X=2.84 $Y=0.48
+ $X2=2.84 $Y2=1.075
r126 31 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.2 $Y=0.48
+ $X2=3.2 $Y2=0.48
r127 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.48 $Y=0.48
+ $X2=2.48 $Y2=0.48
r128 26 32 0.372388 $w=3.7e-07 $l=9.7e-07 $layer=MET1_cond $X=1.51 $Y=0.44
+ $X2=2.48 $Y2=0.44
r129 23 26 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.79 $Y=0.44
+ $X2=1.51 $Y2=0.44
r130 22 28 3.40316 $w=9.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.15 $Y=0.48
+ $X2=1.15 $Y2=0.745
r131 22 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.51 $Y=0.48
+ $X2=1.51 $Y2=0.48
r132 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.79 $Y=0.48
+ $X2=0.79 $Y2=0.48
r133 19 51 1.1402 $w=3.7e-07 $l=2.97e-06 $layer=MET1_cond $X=8.4 $Y=0.44
+ $X2=11.37 $Y2=0.44
r134 19 47 0.134367 $w=3.7e-07 $l=3.5e-07 $layer=MET1_cond $X=8.4 $Y=0.44
+ $X2=8.05 $Y2=0.44
r135 6 75 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=15.49
+ $Y=0.865 $X2=15.745 $Y2=1.16
r136 6 73 182 $w=1.7e-07 $l=3.42491e-07 $layer=licon1_NDIFF $count=1 $X=15.49
+ $Y=0.865 $X2=15.745 $Y2=0.66
r137 5 64 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=13.335
+ $Y=0.705 $X2=13.48 $Y2=0.83
r138 4 54 182 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=1 $X=11.28
+ $Y=0.535 $X2=11.42 $Y2=0.675
r139 3 44 182 $w=1.7e-07 $l=5.3493e-07 $layer=licon1_NDIFF $count=1 $X=7.515
+ $Y=0.865 $X2=8 $Y2=0.76
r140 2 37 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.855
+ $Y=0.865 $X2=3 $Y2=1.075
r141 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.97
+ $Y=0.535 $X2=1.11 $Y2=0.745
.ends

