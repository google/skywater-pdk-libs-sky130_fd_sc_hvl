* File: sky130_fd_sc_hvl__xor2_1.pxi.spice
* Created: Fri Aug 28 09:40:58 2020
* 
x_PM_SKY130_FD_SC_HVL__XOR2_1%VNB N_VNB_M1005_b VNB N_VNB_c_5_p VNB
+ PM_SKY130_FD_SC_HVL__XOR2_1%VNB
x_PM_SKY130_FD_SC_HVL__XOR2_1%VPB N_VPB_M1009_b VPB N_VPB_c_34_p VPB
+ PM_SKY130_FD_SC_HVL__XOR2_1%VPB
x_PM_SKY130_FD_SC_HVL__XOR2_1%B N_B_c_84_n N_B_M1001_g N_B_c_77_n N_B_c_78_n
+ N_B_c_103_p N_B_c_79_n N_B_c_105_p B N_B_M1005_g N_B_M1009_g N_B_M1004_g
+ PM_SKY130_FD_SC_HVL__XOR2_1%B
x_PM_SKY130_FD_SC_HVL__XOR2_1%A N_A_c_148_n N_A_M1007_g N_A_M1008_g N_A_c_151_n
+ N_A_M1006_g N_A_c_145_n N_A_M1003_g A A A N_A_c_147_n
+ PM_SKY130_FD_SC_HVL__XOR2_1%A
x_PM_SKY130_FD_SC_HVL__XOR2_1%A_30_443# N_A_30_443#_M1005_d N_A_30_443#_M1009_s
+ N_A_30_443#_M1002_g N_A_30_443#_c_199_n N_A_30_443#_M1000_g
+ N_A_30_443#_c_193_n N_A_30_443#_c_203_n N_A_30_443#_c_194_n
+ N_A_30_443#_c_195_n N_A_30_443#_c_217_n N_A_30_443#_c_196_n
+ N_A_30_443#_c_206_n N_A_30_443#_c_249_p N_A_30_443#_c_207_n
+ N_A_30_443#_c_223_n N_A_30_443#_c_255_p N_A_30_443#_c_198_n
+ PM_SKY130_FD_SC_HVL__XOR2_1%A_30_443#
x_PM_SKY130_FD_SC_HVL__XOR2_1%VPWR N_VPWR_M1007_d N_VPWR_M1001_d VPWR
+ N_VPWR_c_271_n N_VPWR_c_274_n N_VPWR_c_277_n PM_SKY130_FD_SC_HVL__XOR2_1%VPWR
x_PM_SKY130_FD_SC_HVL__XOR2_1%A_531_443# N_A_531_443#_M1006_d
+ N_A_531_443#_M1000_d N_A_531_443#_c_321_n N_A_531_443#_c_308_n
+ N_A_531_443#_c_311_n N_A_531_443#_c_312_n N_A_531_443#_c_313_n
+ N_A_531_443#_c_316_n PM_SKY130_FD_SC_HVL__XOR2_1%A_531_443#
x_PM_SKY130_FD_SC_HVL__XOR2_1%X N_X_M1004_d N_X_M1000_s X X X X N_X_c_341_n X
+ PM_SKY130_FD_SC_HVL__XOR2_1%X
x_PM_SKY130_FD_SC_HVL__XOR2_1%VGND N_VGND_M1005_s N_VGND_M1008_d N_VGND_M1002_d
+ VGND N_VGND_c_361_n N_VGND_c_363_n N_VGND_c_365_n N_VGND_c_367_n
+ PM_SKY130_FD_SC_HVL__XOR2_1%VGND
cc_1 N_VNB_M1005_b N_B_c_77_n 0.0111991f $X=-0.33 $Y=-0.265 $X2=3.545 $Y2=1.855
cc_2 N_VNB_M1005_b N_B_c_78_n 0.00413046f $X=-0.33 $Y=-0.265 $X2=1.34 $Y2=1.915
cc_3 N_VNB_M1005_b N_B_c_79_n 0.00354401f $X=-0.33 $Y=-0.265 $X2=3.415 $Y2=1.51
cc_4 N_VNB_M1005_b N_B_M1005_g 0.0950456f $X=-0.33 $Y=-0.265 $X2=0.685 $Y2=0.91
cc_5 N_VNB_c_5_p N_B_M1005_g 0.00119158f $X=0.24 $Y=0 $X2=0.685 $Y2=0.91
cc_6 N_VNB_M1005_b N_B_M1004_g 0.0823591f $X=-0.33 $Y=-0.265 $X2=3.545 $Y2=0.91
cc_7 N_VNB_c_5_p N_B_M1004_g 5.81826e-19 $X=0.24 $Y=0 $X2=3.545 $Y2=0.91
cc_8 N_VNB_M1005_b N_A_M1008_g 0.0477121f $X=-0.33 $Y=-0.265 $X2=3.545 $Y2=1.98
cc_9 N_VNB_c_5_p N_A_M1008_g 5.81826e-19 $X=0.24 $Y=0 $X2=3.545 $Y2=1.98
cc_10 N_VNB_M1005_b N_A_c_145_n 0.0420545f $X=-0.33 $Y=-0.265 $X2=0.725 $Y2=1.89
cc_11 N_VNB_M1005_b A 0.00461555f $X=-0.33 $Y=-0.265 $X2=3.415 $Y2=1.51
cc_12 N_VNB_M1005_b N_A_c_147_n 0.137285f $X=-0.33 $Y=-0.265 $X2=0.685 $Y2=2.965
cc_13 N_VNB_M1005_b N_A_30_443#_M1002_g 0.0750201f $X=-0.33 $Y=-0.265 $X2=1.34
+ $Y2=1.915
cc_14 N_VNB_c_5_p N_A_30_443#_M1002_g 0.00221559f $X=0.24 $Y=0 $X2=1.34
+ $Y2=1.915
cc_15 N_VNB_M1005_b N_A_30_443#_c_193_n 0.0146038f $X=-0.33 $Y=-0.265 $X2=1.51
+ $Y2=1.51
cc_16 N_VNB_M1005_b N_A_30_443#_c_194_n 0.00577343f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.965
cc_17 N_VNB_M1005_b N_A_30_443#_c_195_n 0.0100989f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.965
cc_18 N_VNB_M1005_b N_A_30_443#_c_196_n 0.0101821f $X=-0.33 $Y=-0.265 $X2=3.545
+ $Y2=1.67
cc_19 N_VNB_c_5_p N_A_30_443#_c_196_n 6.32535e-19 $X=0.24 $Y=0 $X2=3.545
+ $Y2=1.67
cc_20 N_VNB_M1005_b N_A_30_443#_c_198_n 0.0528038f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_21 N_VNB_M1005_b X 0.00962907f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_22 N_VNB_M1005_b N_X_c_341_n 0.015149f $X=-0.33 $Y=-0.265 $X2=3.515 $Y2=1.58
cc_23 N_VNB_c_5_p N_X_c_341_n 0.00184286f $X=0.24 $Y=0 $X2=3.515 $Y2=1.58
cc_24 N_VNB_M1005_b N_VGND_c_361_n 0.0614067f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_25 N_VNB_c_5_p N_VGND_c_361_n 0.00166879f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_26 N_VNB_M1005_b N_VGND_c_363_n 0.116714f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_27 N_VNB_c_5_p N_VGND_c_363_n 0.00660266f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_28 N_VNB_M1005_b N_VGND_c_365_n 0.0836368f $X=-0.33 $Y=-0.265 $X2=3.545
+ $Y2=1.67
cc_29 N_VNB_c_5_p N_VGND_c_365_n 0.00166879f $X=0.24 $Y=0 $X2=3.545 $Y2=1.67
cc_30 N_VNB_M1005_b N_VGND_c_367_n 0.0863165f $X=-0.33 $Y=-0.265 $X2=3.565
+ $Y2=1.67
cc_31 N_VNB_c_5_p N_VGND_c_367_n 0.564546f $X=0.24 $Y=0 $X2=3.565 $Y2=1.67
cc_32 N_VPB_M1009_b N_B_c_84_n 0.0376872f $X=-0.33 $Y=1.885 $X2=3.185 $Y2=2.105
cc_33 VPB N_B_c_84_n 0.00970178f $X=0 $Y=3.955 $X2=3.185 $Y2=2.105
cc_34 N_VPB_c_34_p N_B_c_84_n 0.015205f $X=5.04 $Y=4.07 $X2=3.185 $Y2=2.105
cc_35 N_VPB_M1009_b N_B_c_77_n 0.039288f $X=-0.33 $Y=1.885 $X2=3.545 $Y2=1.855
cc_36 N_VPB_M1009_b N_B_c_78_n 0.0026938f $X=-0.33 $Y=1.885 $X2=1.34 $Y2=1.915
cc_37 N_VPB_M1009_b N_B_M1005_g 0.0561778f $X=-0.33 $Y=1.885 $X2=0.685 $Y2=0.91
cc_38 VPB N_B_M1005_g 0.00970178f $X=0 $Y=3.955 $X2=0.685 $Y2=0.91
cc_39 N_VPB_c_34_p N_B_M1005_g 0.0152133f $X=5.04 $Y=4.07 $X2=0.685 $Y2=0.91
cc_40 N_VPB_M1009_b N_A_c_148_n 0.0345202f $X=-0.33 $Y=1.885 $X2=3.185 $Y2=2.105
cc_41 VPB N_A_c_148_n 0.00970178f $X=0 $Y=3.955 $X2=3.185 $Y2=2.105
cc_42 N_VPB_c_34_p N_A_c_148_n 0.0137101f $X=5.04 $Y=4.07 $X2=3.185 $Y2=2.105
cc_43 N_VPB_M1009_b N_A_c_151_n 0.0347709f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_44 VPB N_A_c_151_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_45 N_VPB_c_34_p N_A_c_151_n 0.0152133f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_46 N_VPB_M1009_b A 0.00503207f $X=-0.33 $Y=1.885 $X2=3.415 $Y2=1.51
cc_47 N_VPB_M1009_b N_A_c_147_n 0.0503613f $X=-0.33 $Y=1.885 $X2=0.685 $Y2=2.965
cc_48 N_VPB_M1009_b N_A_30_443#_c_199_n 0.0429698f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=1.89
cc_49 VPB N_A_30_443#_c_199_n 0.00970178f $X=0 $Y=3.955 $X2=0.725 $Y2=1.89
cc_50 N_VPB_c_34_p N_A_30_443#_c_199_n 0.015205f $X=5.04 $Y=4.07 $X2=0.725
+ $Y2=1.89
cc_51 N_VPB_M1009_b N_A_30_443#_c_193_n 0.0254803f $X=-0.33 $Y=1.885 $X2=1.51
+ $Y2=1.51
cc_52 N_VPB_M1009_b N_A_30_443#_c_203_n 0.0365978f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=0.91
cc_53 VPB N_A_30_443#_c_203_n 7.60114e-19 $X=0 $Y=3.955 $X2=0.685 $Y2=0.91
cc_54 N_VPB_c_34_p N_A_30_443#_c_203_n 0.0131049f $X=5.04 $Y=4.07 $X2=0.685
+ $Y2=0.91
cc_55 N_VPB_M1009_b N_A_30_443#_c_206_n 0.0130122f $X=-0.33 $Y=1.885 $X2=3.565
+ $Y2=1.67
cc_56 N_VPB_M1009_b N_A_30_443#_c_207_n 0.00704942f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_57 N_VPB_M1009_b N_A_30_443#_c_198_n 0.0449828f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_58 N_VPB_M1009_b N_VPWR_c_271_n 0.00343705f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=1.915
cc_59 VPB N_VPWR_c_271_n 0.00819601f $X=0 $Y=3.955 $X2=0.725 $Y2=1.915
cc_60 N_VPB_c_34_p N_VPWR_c_271_n 0.0990548f $X=5.04 $Y=4.07 $X2=0.725 $Y2=1.915
cc_61 N_VPB_M1009_b N_VPWR_c_274_n 0.0132463f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_274_n 0.0062727f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_63 N_VPB_c_34_p N_VPWR_c_274_n 0.0839896f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_64 N_VPB_M1009_b N_VPWR_c_277_n 0.0504527f $X=-0.33 $Y=1.885 $X2=3.545
+ $Y2=0.91
cc_65 VPB N_VPWR_c_277_n 0.56022f $X=0 $Y=3.955 $X2=3.545 $Y2=0.91
cc_66 N_VPB_c_34_p N_VPWR_c_277_n 0.0220721f $X=5.04 $Y=4.07 $X2=3.545 $Y2=0.91
cc_67 N_VPB_M1009_b N_A_531_443#_c_308_n 0.00127492f $X=-0.33 $Y=1.885 $X2=1.34
+ $Y2=1.915
cc_68 VPB N_A_531_443#_c_308_n 5.14916e-19 $X=0 $Y=3.955 $X2=1.34 $Y2=1.915
cc_69 N_VPB_c_34_p N_A_531_443#_c_308_n 0.00887752f $X=5.04 $Y=4.07 $X2=1.34
+ $Y2=1.915
cc_70 N_VPB_M1009_b N_A_531_443#_c_311_n 0.00806673f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=1.89
cc_71 N_VPB_M1009_b N_A_531_443#_c_312_n 0.0392785f $X=-0.33 $Y=1.885 $X2=1.425
+ $Y2=1.775
cc_72 N_VPB_M1009_b N_A_531_443#_c_313_n 0.0174969f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_73 VPB N_A_531_443#_c_313_n 7.60114e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_74 N_VPB_c_34_p N_A_531_443#_c_313_n 0.0131049f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_75 N_VPB_M1009_b N_A_531_443#_c_316_n 0.00704942f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=1.89
cc_76 N_VPB_M1009_b X 0.00842641f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_77 N_B_M1005_g N_A_M1008_g 0.0390642f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_78 N_B_c_84_n N_A_c_151_n 0.0321713f $X=3.185 $Y=2.105 $X2=0 $Y2=0
cc_79 N_B_M1004_g N_A_c_145_n 0.0839214f $X=3.545 $Y=0.91 $X2=0.24 $Y2=0
cc_80 N_B_c_84_n A 0.00930008f $X=3.185 $Y=2.105 $X2=5.04 $Y2=0
cc_81 N_B_c_77_n A 0.025289f $X=3.545 $Y=1.855 $X2=5.04 $Y2=0
cc_82 N_B_c_78_n A 0.00917551f $X=1.34 $Y=1.915 $X2=5.04 $Y2=0
cc_83 N_B_c_79_n A 0.0850219f $X=3.415 $Y=1.51 $X2=5.04 $Y2=0
cc_84 B A 0.00475644f $X=3.515 $Y=1.58 $X2=5.04 $Y2=0
cc_85 N_B_M1004_g A 0.00162635f $X=3.545 $Y=0.91 $X2=5.04 $Y2=0
cc_86 N_B_c_77_n N_A_c_147_n 0.0420942f $X=3.545 $Y=1.855 $X2=2.64 $Y2=0.058
cc_87 N_B_c_78_n N_A_c_147_n 0.0343944f $X=1.34 $Y=1.915 $X2=2.64 $Y2=0.058
cc_88 N_B_c_103_p N_A_c_147_n 0.0133413f $X=1.425 $Y=1.775 $X2=2.64 $Y2=0.058
cc_89 N_B_c_79_n N_A_c_147_n 0.0755539f $X=3.415 $Y=1.51 $X2=2.64 $Y2=0.058
cc_90 N_B_c_105_p N_A_c_147_n 0.00662797f $X=1.51 $Y=1.51 $X2=2.64 $Y2=0.058
cc_91 B N_A_c_147_n 2.95119e-19 $X=3.515 $Y=1.58 $X2=2.64 $Y2=0.058
cc_92 N_B_M1005_g N_A_c_147_n 0.138454f $X=0.685 $Y=0.91 $X2=2.64 $Y2=0.058
cc_93 N_B_M1004_g N_A_c_147_n 0.00474554f $X=3.545 $Y=0.91 $X2=2.64 $Y2=0.058
cc_94 B N_A_30_443#_M1002_g 3.79552e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_95 N_B_M1004_g N_A_30_443#_M1002_g 0.0241097f $X=3.545 $Y=0.91 $X2=0 $Y2=0
cc_96 N_B_c_78_n N_A_30_443#_c_193_n 0.0218761f $X=1.34 $Y=1.915 $X2=5.04 $Y2=0
cc_97 N_B_M1005_g N_A_30_443#_c_193_n 0.023819f $X=0.685 $Y=0.91 $X2=5.04 $Y2=0
cc_98 N_B_M1005_g N_A_30_443#_c_203_n 0.00260632f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_99 N_B_c_78_n N_A_30_443#_c_194_n 0.0443049f $X=1.34 $Y=1.915 $X2=2.64
+ $Y2=0.058
cc_100 N_B_c_105_p N_A_30_443#_c_194_n 0.0145092f $X=1.51 $Y=1.51 $X2=2.64
+ $Y2=0.058
cc_101 N_B_M1005_g N_A_30_443#_c_194_n 0.0372598f $X=0.685 $Y=0.91 $X2=2.64
+ $Y2=0.058
cc_102 N_B_c_84_n N_A_30_443#_c_217_n 0.00981169f $X=3.185 $Y=2.105 $X2=0 $Y2=0
cc_103 N_B_c_78_n N_A_30_443#_c_217_n 0.034563f $X=1.34 $Y=1.915 $X2=0 $Y2=0
cc_104 N_B_M1005_g N_A_30_443#_c_217_n 0.0341798f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_105 N_B_M1005_g N_A_30_443#_c_196_n 0.0240466f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_106 N_B_c_84_n N_A_30_443#_c_206_n 0.0202931f $X=3.185 $Y=2.105 $X2=0 $Y2=0
cc_107 N_B_c_77_n N_A_30_443#_c_206_n 0.00987234f $X=3.545 $Y=1.855 $X2=0 $Y2=0
cc_108 N_B_c_84_n N_A_30_443#_c_223_n 0.0212035f $X=3.185 $Y=2.105 $X2=0 $Y2=0
cc_109 N_B_c_77_n N_A_30_443#_c_198_n 0.0241097f $X=3.545 $Y=1.855 $X2=0 $Y2=0
cc_110 N_B_M1005_g N_VPWR_c_271_n 0.0575682f $X=0.685 $Y=0.91 $X2=0.24 $Y2=0
cc_111 N_B_c_84_n N_VPWR_c_274_n 0.0273029f $X=3.185 $Y=2.105 $X2=0 $Y2=0
cc_112 N_B_c_84_n N_VPWR_c_277_n 0.00428953f $X=3.185 $Y=2.105 $X2=0 $Y2=0
cc_113 N_B_M1005_g N_VPWR_c_277_n 0.00846141f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_114 N_B_c_84_n N_A_531_443#_c_308_n 0.00199892f $X=3.185 $Y=2.105 $X2=0 $Y2=0
cc_115 N_B_c_84_n N_A_531_443#_c_311_n 0.0273029f $X=3.185 $Y=2.105 $X2=0.24
+ $Y2=0
cc_116 N_B_c_84_n X 0.0095186f $X=3.185 $Y=2.105 $X2=0 $Y2=0
cc_117 B X 0.0239088f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_118 N_B_M1004_g X 0.0130211f $X=3.545 $Y=0.91 $X2=0 $Y2=0
cc_119 N_B_M1004_g N_X_c_341_n 0.00223015f $X=3.545 $Y=0.91 $X2=0 $Y2=0
cc_120 N_B_M1005_g N_VGND_c_361_n 0.0441237f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_121 N_B_c_79_n N_VGND_c_363_n 0.131884f $X=3.415 $Y=1.51 $X2=0 $Y2=0
cc_122 N_B_c_105_p N_VGND_c_363_n 0.0135978f $X=1.51 $Y=1.51 $X2=0 $Y2=0
cc_123 B N_VGND_c_363_n 0.0179963f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_124 N_B_M1005_g N_VGND_c_363_n 7.04443e-19 $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_125 N_B_M1004_g N_VGND_c_363_n 0.0560885f $X=3.545 $Y=0.91 $X2=0 $Y2=0
cc_126 N_B_M1005_g N_VGND_c_367_n 0.0140308f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_127 N_B_M1004_g N_VGND_c_367_n 0.00772948f $X=3.545 $Y=0.91 $X2=0 $Y2=0
cc_128 N_A_c_147_n N_A_30_443#_c_194_n 0.00180904f $X=2.405 $Y=1.75 $X2=2.64
+ $Y2=0.058
cc_129 N_A_c_148_n N_A_30_443#_c_217_n 0.0332631f $X=1.395 $Y=2.105 $X2=0 $Y2=0
cc_130 N_A_c_151_n N_A_30_443#_c_217_n 0.0328458f $X=2.405 $Y=2.105 $X2=0 $Y2=0
cc_131 A N_A_30_443#_c_217_n 0.0468433f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_132 N_A_c_147_n N_A_30_443#_c_217_n 0.0109032f $X=2.405 $Y=1.75 $X2=0 $Y2=0
cc_133 N_A_M1008_g N_A_30_443#_c_196_n 0.00473603f $X=1.465 $Y=0.91 $X2=0 $Y2=0
cc_134 N_A_c_151_n N_A_30_443#_c_223_n 9.75909e-19 $X=2.405 $Y=2.105 $X2=0 $Y2=0
cc_135 A N_A_30_443#_c_223_n 0.00847132f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_136 N_A_c_148_n N_VPWR_c_271_n 0.0648537f $X=1.395 $Y=2.105 $X2=0.24 $Y2=0
cc_137 N_A_c_151_n N_VPWR_c_271_n 0.0660048f $X=2.405 $Y=2.105 $X2=0.24 $Y2=0
cc_138 N_A_c_148_n N_VPWR_c_277_n 0.00207887f $X=1.395 $Y=2.105 $X2=0 $Y2=0
cc_139 N_A_c_151_n N_VPWR_c_277_n 0.00803362f $X=2.405 $Y=2.105 $X2=0 $Y2=0
cc_140 N_A_c_151_n N_A_531_443#_c_308_n 0.00198688f $X=2.405 $Y=2.105 $X2=0
+ $Y2=0
cc_141 N_A_M1008_g N_VGND_c_361_n 5.11463e-19 $X=1.465 $Y=0.91 $X2=0 $Y2=0
cc_142 N_A_M1008_g N_VGND_c_363_n 0.0534373f $X=1.465 $Y=0.91 $X2=0 $Y2=0
cc_143 N_A_c_145_n N_VGND_c_363_n 0.0828313f $X=2.835 $Y=1.395 $X2=0 $Y2=0
cc_144 N_A_c_147_n N_VGND_c_363_n 0.0236609f $X=2.405 $Y=1.75 $X2=0 $Y2=0
cc_145 N_A_M1008_g N_VGND_c_367_n 0.00772948f $X=1.465 $Y=0.91 $X2=0 $Y2=0
cc_146 N_A_30_443#_c_217_n A_187_443# 0.00254458f $X=3.06 $Y=2.52 $X2=0 $Y2=0
cc_147 N_A_30_443#_c_217_n N_VPWR_M1007_d 0.011726f $X=3.06 $Y=2.52 $X2=0 $Y2=0
cc_148 N_A_30_443#_c_206_n N_VPWR_M1001_d 0.00697699f $X=4.55 $Y=2.69 $X2=0
+ $Y2=0
cc_149 N_A_30_443#_c_203_n N_VPWR_c_271_n 0.041864f $X=0.295 $Y=2.755 $X2=0.24
+ $Y2=0
cc_150 N_A_30_443#_c_217_n N_VPWR_c_271_n 0.129096f $X=3.06 $Y=2.52 $X2=0.24
+ $Y2=0
cc_151 N_A_30_443#_c_199_n N_VPWR_c_274_n 0.0368618f $X=4.595 $Y=2.105 $X2=0
+ $Y2=0
cc_152 N_A_30_443#_M1009_s N_VPWR_c_277_n 0.00221032f $X=0.15 $Y=2.215 $X2=0
+ $Y2=0
cc_153 N_A_30_443#_c_199_n N_VPWR_c_277_n 0.00500332f $X=4.595 $Y=2.105 $X2=0
+ $Y2=0
cc_154 N_A_30_443#_c_203_n N_VPWR_c_277_n 0.0354327f $X=0.295 $Y=2.755 $X2=0
+ $Y2=0
cc_155 N_A_30_443#_c_217_n N_A_531_443#_M1006_d 0.00404642f $X=3.06 $Y=2.52
+ $X2=0 $Y2=0
cc_156 N_A_30_443#_c_217_n N_A_531_443#_c_321_n 0.0129403f $X=3.06 $Y=2.52 $X2=0
+ $Y2=0
cc_157 N_A_30_443#_c_199_n N_A_531_443#_c_311_n 0.0307871f $X=4.595 $Y=2.105
+ $X2=0.24 $Y2=0
cc_158 N_A_30_443#_c_217_n N_A_531_443#_c_311_n 0.00472848f $X=3.06 $Y=2.52
+ $X2=0.24 $Y2=0
cc_159 N_A_30_443#_c_206_n N_A_531_443#_c_311_n 0.0951326f $X=4.55 $Y=2.69
+ $X2=0.24 $Y2=0
cc_160 N_A_30_443#_c_223_n N_A_531_443#_c_311_n 0.0115442f $X=3.145 $Y=2.52
+ $X2=0.24 $Y2=0
cc_161 N_A_30_443#_c_199_n N_A_531_443#_c_312_n 0.00188943f $X=4.595 $Y=2.105
+ $X2=0 $Y2=0
cc_162 N_A_30_443#_c_249_p N_A_531_443#_c_312_n 0.0153818f $X=4.635 $Y=2.605
+ $X2=0 $Y2=0
cc_163 N_A_30_443#_c_199_n N_A_531_443#_c_313_n 0.00186266f $X=4.595 $Y=2.105
+ $X2=0 $Y2=0
cc_164 N_A_30_443#_c_206_n N_X_M1000_s 0.00568641f $X=4.55 $Y=2.69 $X2=0 $Y2=0
cc_165 N_A_30_443#_M1002_g X 0.0328435f $X=4.325 $Y=0.91 $X2=0 $Y2=0
cc_166 N_A_30_443#_c_199_n X 0.00800827f $X=4.595 $Y=2.105 $X2=0 $Y2=0
cc_167 N_A_30_443#_c_206_n X 0.0271029f $X=4.55 $Y=2.69 $X2=0 $Y2=0
cc_168 N_A_30_443#_c_255_p X 0.0537523f $X=4.715 $Y=1.83 $X2=0 $Y2=0
cc_169 N_A_30_443#_c_198_n X 0.0317518f $X=4.715 $Y=1.83 $X2=0 $Y2=0
cc_170 N_A_30_443#_M1002_g N_X_c_341_n 0.0268989f $X=4.325 $Y=0.91 $X2=0 $Y2=0
cc_171 N_A_30_443#_c_194_n N_VGND_c_361_n 0.0196695f $X=0.91 $Y=1.51 $X2=0 $Y2=0
cc_172 N_A_30_443#_c_195_n N_VGND_c_361_n 0.0219893f $X=0.38 $Y=1.51 $X2=0 $Y2=0
cc_173 N_A_30_443#_c_196_n N_VGND_c_361_n 0.0435428f $X=1.075 $Y=0.66 $X2=0
+ $Y2=0
cc_174 N_A_30_443#_M1002_g N_VGND_c_363_n 0.00110154f $X=4.325 $Y=0.91 $X2=0
+ $Y2=0
cc_175 N_A_30_443#_c_196_n N_VGND_c_363_n 0.0317942f $X=1.075 $Y=0.66 $X2=0
+ $Y2=0
cc_176 N_A_30_443#_M1002_g N_VGND_c_365_n 0.0227925f $X=4.325 $Y=0.91 $X2=0
+ $Y2=0
cc_177 N_A_30_443#_c_255_p N_VGND_c_365_n 0.0168751f $X=4.715 $Y=1.83 $X2=0
+ $Y2=0
cc_178 N_A_30_443#_c_198_n N_VGND_c_365_n 0.00874988f $X=4.715 $Y=1.83 $X2=0
+ $Y2=0
cc_179 N_A_30_443#_M1005_d N_VGND_c_367_n 0.00221032f $X=0.935 $Y=0.535 $X2=0
+ $Y2=0
cc_180 N_A_30_443#_M1002_g N_VGND_c_367_n 0.0137947f $X=4.325 $Y=0.91 $X2=0
+ $Y2=0
cc_181 N_A_30_443#_c_196_n N_VGND_c_367_n 0.0246119f $X=1.075 $Y=0.66 $X2=0
+ $Y2=0
cc_182 A_187_443# N_VPWR_c_271_n 0.00109099f $X=0.935 $Y=2.215 $X2=0 $Y2=0
cc_183 N_VPWR_c_277_n N_A_531_443#_M1006_d 0.00275991f $X=4.61 $Y=3.59 $X2=0
+ $Y2=3.985
cc_184 N_VPWR_c_277_n N_A_531_443#_M1000_d 5.49589e-19 $X=4.61 $Y=3.59 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_271_n N_A_531_443#_c_308_n 0.028177f $X=1.785 $Y=2.87 $X2=0.24
+ $Y2=4.07
cc_186 N_VPWR_c_274_n N_A_531_443#_c_308_n 0.0209803f $X=4.61 $Y=3.59 $X2=0.24
+ $Y2=4.07
cc_187 N_VPWR_c_277_n N_A_531_443#_c_308_n 0.0229098f $X=4.61 $Y=3.59 $X2=0.24
+ $Y2=4.07
cc_188 N_VPWR_M1001_d N_A_531_443#_c_311_n 0.00581692f $X=3.435 $Y=2.215 $X2=0
+ $Y2=0
cc_189 N_VPWR_c_274_n N_A_531_443#_c_311_n 0.105573f $X=4.61 $Y=3.59 $X2=0 $Y2=0
cc_190 N_VPWR_c_277_n N_A_531_443#_c_311_n 0.0219322f $X=4.61 $Y=3.59 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_274_n N_A_531_443#_c_313_n 0.0210514f $X=4.61 $Y=3.59 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_277_n N_A_531_443#_c_313_n 0.0354073f $X=4.61 $Y=3.59 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_274_n N_X_M1000_s 0.00494129f $X=4.61 $Y=3.59 $X2=0 $Y2=0
cc_194 N_A_531_443#_c_311_n N_X_M1000_s 0.00581692f $X=4.9 $Y=3.04 $X2=0 $Y2=0
cc_195 N_X_c_341_n N_VGND_c_363_n 0.0318609f $X=3.935 $Y=0.66 $X2=0 $Y2=0
cc_196 N_X_c_341_n N_VGND_c_365_n 0.062271f $X=3.935 $Y=0.66 $X2=0 $Y2=0
cc_197 N_X_M1004_d N_VGND_c_367_n 0.00221032f $X=3.795 $Y=0.535 $X2=0 $Y2=0
cc_198 N_X_c_341_n N_VGND_c_367_n 0.047798f $X=3.935 $Y=0.66 $X2=0 $Y2=0
cc_199 N_VGND_c_363_n A_617_107# 9.69903e-19 $X=3.585 $Y=0.48 $X2=0 $Y2=0
