* File: sky130_fd_sc_hvl__sdfrbp_1.pex.spice
* Created: Wed Sep  2 09:09:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%VNB 5 7 11
c148 11 0 1.72602e-20 $X=0.24 $Y=0
r149 7 11 0.000353423 $w=2.016e-05 $l=5.7e-08 $layer=MET1_cond $X=10.08 $Y=0.057
+ $X2=10.08 $Y2=0
r150 5 11 0.442857 $w=1.7e-07 $l=3.57e-06 $layer=mcon $count=21 $X=19.92 $Y=0
+ $X2=19.92 $Y2=0
r151 5 11 0.442857 $w=1.7e-07 $l=3.57e-06 $layer=mcon $count=21 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%VPB 4 6 14
r210 10 14 0.442857 $w=1.7e-07 $l=3.57e-06 $layer=mcon $count=21 $X=19.92
+ $Y=4.07 $X2=19.92 $Y2=4.07
r211 9 14 1283.94 $w=1.68e-07 $l=1.968e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=19.92 $Y2=4.07
r212 9 10 0.442857 $w=1.7e-07 $l=3.57e-06 $layer=mcon $count=21 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r213 6 10 0.000353423 $w=2.016e-05 $l=5.7e-08 $layer=MET1_cond $X=10.08 $Y=4.013
+ $X2=10.08 $Y2=4.07
r214 4 14 8.66667 $w=1.7e-07 $l=1.99625e-05 $layer=licon1_NTAP_notbjt $count=21
+ $X=0 $Y=3.985 $X2=19.92 $Y2=4.07
r215 4 9 8.66667 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=21
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%SCE 3 7 10 13 17 25 26 28 30 33 36 37 41
+ 43 44 48 55 59 63
c125 33 0 7.00078e-20 $X=2.875 $Y=2.75
c126 25 0 1.16047e-19 $X=1.515 $Y=0.35
r127 59 61 5.31017 $w=5.9e-07 $l=6.5e-08 $layer=POLY_cond $X=3.765 $Y=1.507
+ $X2=3.83 $Y2=1.507
r128 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.765
+ $Y=1.365 $X2=3.765 $Y2=1.365
r129 44 60 7.24547 $w=5.18e-07 $l=3.15e-07 $layer=LI1_cond $X=4.08 $Y=1.535
+ $X2=3.765 $Y2=1.535
r130 43 60 3.79525 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.6 $Y=1.535
+ $X2=3.765 $Y2=1.535
r131 43 63 8.49122 $w=5.18e-07 $l=1.15e-07 $layer=LI1_cond $X=3.6 $Y=1.535
+ $X2=3.485 $Y2=1.535
r132 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=2.83 $X2=1.6 $Y2=2.83
r133 37 40 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.64 $Y=2.75 $X2=1.64
+ $Y2=2.83
r134 34 55 131.991 $w=2.4e-07 $l=5.1e-07 $layer=POLY_cond $X=2.875 $Y=2.685
+ $X2=3.385 $Y2=2.685
r135 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.875
+ $Y=2.75 $X2=2.875 $Y2=2.75
r136 31 37 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.765 $Y=2.75
+ $X2=1.64 $Y2=2.75
r137 31 33 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=1.765 $Y=2.75
+ $X2=2.875 $Y2=2.75
r138 30 63 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=1.685 $Y=1.36
+ $X2=3.485 $Y2=1.36
r139 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.6 $Y=1.275
+ $X2=1.685 $Y2=1.36
r140 27 28 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.6 $Y=0.435
+ $X2=1.6 $Y2=1.275
r141 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.515 $Y=0.35
+ $X2=1.6 $Y2=0.435
r142 25 26 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.515 $Y=0.35
+ $X2=0.985 $Y2=0.35
r143 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.9 $Y=0.435
+ $X2=0.985 $Y2=0.35
r144 23 36 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.9 $Y=0.435 $X2=0.9
+ $Y2=1.295
r145 21 48 63.6685 $w=5e-07 $l=5.95e-07 $layer=POLY_cond $X=0.86 $Y=1.46
+ $X2=0.86 $Y2=0.865
r146 20 36 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.82 $Y=1.46
+ $X2=0.82 $Y2=1.295
r147 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.82
+ $Y=1.46 $X2=0.82 $Y2=1.46
r148 16 41 52.4329 $w=5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.11 $Y=2.865 $X2=1.6
+ $Y2=2.865
r149 16 17 5.30422 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.11 $Y=2.865
+ $X2=0.86 $Y2=2.865
r150 15 21 123.592 $w=5e-07 $l=1.155e-06 $layer=POLY_cond $X=0.86 $Y=2.615
+ $X2=0.86 $Y2=1.46
r151 15 17 20.4101 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.86 $Y=2.615
+ $X2=0.86 $Y2=2.865
r152 11 61 6.7465 $w=5e-07 $l=3.82e-07 $layer=POLY_cond $X=3.83 $Y=1.125
+ $X2=3.83 $Y2=1.507
r153 11 13 40.6622 $w=5e-07 $l=3.8e-07 $layer=POLY_cond $X=3.83 $Y=1.125
+ $X2=3.83 $Y2=0.745
r154 10 55 3.85076 $w=2.3e-07 $l=1.2e-07 $layer=POLY_cond $X=3.385 $Y=2.565
+ $X2=3.385 $Y2=2.685
r155 9 59 31.0441 $w=5.9e-07 $l=5.40582e-07 $layer=POLY_cond $X=3.385 $Y=1.89
+ $X2=3.765 $Y2=1.507
r156 9 10 188.33 $w=2.3e-07 $l=6.75e-07 $layer=POLY_cond $X=3.385 $Y=1.89
+ $X2=3.385 $Y2=2.565
r157 7 34 72.764 $w=5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.94 $Y=3.485 $X2=2.94
+ $Y2=2.805
r158 1 17 20.4101 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.86 $Y=3.115 $X2=0.86
+ $Y2=2.865
r159 1 3 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.86 $Y=3.115 $X2=0.86
+ $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%D 1 3 7 9 13
c39 7 0 1.16047e-19 $X=2.34 $Y=0.745
r40 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.165
+ $Y=1.71 $X2=2.165 $Y2=1.71
r41 9 13 11.3745 $w=5.08e-07 $l=4.85e-07 $layer=LI1_cond $X=1.68 $Y=1.88
+ $X2=2.165 $Y2=1.88
r42 5 12 52.538 $w=5e-07 $l=5.71839e-07 $layer=POLY_cond $X=2.34 $Y=1.165
+ $X2=2.285 $Y2=1.71
r43 5 7 44.9425 $w=5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.34 $Y=1.165 $X2=2.34
+ $Y2=0.745
r44 1 12 6.266 $w=5e-07 $l=8.83176e-08 $layer=POLY_cond $X=2.23 $Y=1.775
+ $X2=2.285 $Y2=1.71
r45 1 3 182.98 $w=5e-07 $l=1.71e-06 $layer=POLY_cond $X=2.23 $Y=1.775 $X2=2.23
+ $Y2=3.485
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%A_222_131# 1 2 9 13 15 18 19 24 28 30 32
+ 36 37 39 42 43 44 47 48 50 51 52
c135 43 0 1.78387e-19 $X=4.35 $Y=2.75
c136 9 0 8.22034e-20 $X=3.05 $Y=0.745
r137 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.515
+ $Y=2.41 $X2=4.515 $Y2=2.41
r138 45 47 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.515 $Y=2.665
+ $X2=4.515 $Y2=2.41
r139 43 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.35 $Y=2.75
+ $X2=4.515 $Y2=2.665
r140 43 44 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=4.35 $Y=2.75
+ $X2=3.44 $Y2=2.75
r141 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.355 $Y=2.665
+ $X2=3.44 $Y2=2.75
r142 41 42 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.355 $Y=2.485
+ $X2=3.355 $Y2=2.665
r143 40 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=2.4
+ $X2=2.895 $Y2=2.4
r144 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.27 $Y=2.4
+ $X2=3.355 $Y2=2.485
r145 39 40 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.27 $Y=2.4
+ $X2=3.06 $Y2=2.4
r146 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.895
+ $Y=1.79 $X2=2.895 $Y2=1.79
r147 34 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=2.315
+ $X2=2.895 $Y2=2.4
r148 34 36 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=2.895 $Y=2.315
+ $X2=2.895 $Y2=1.79
r149 33 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.335 $Y=2.4
+ $X2=1.25 $Y2=2.4
r150 32 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=2.4
+ $X2=2.895 $Y2=2.4
r151 32 33 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=2.73 $Y=2.4
+ $X2=1.335 $Y2=2.4
r152 28 51 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=1.29 $Y2=3.205
r153 28 30 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=1.29 $Y2=3.455
r154 26 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=2.485
+ $X2=1.25 $Y2=2.4
r155 26 51 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.25 $Y=2.485
+ $X2=1.25 $Y2=3.205
r156 22 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=2.315
+ $X2=1.25 $Y2=2.4
r157 22 24 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=1.25 $Y=2.315
+ $X2=1.25 $Y2=0.865
r158 21 48 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=4.515 $Y=2.77
+ $X2=4.515 $Y2=2.41
r159 18 37 31.6089 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.895 $Y=1.625
+ $X2=2.895 $Y2=1.79
r160 18 19 48.974 $w=2.6e-07 $l=2.05e-07 $layer=POLY_cond $X=2.93 $Y=1.625
+ $X2=2.93 $Y2=1.42
r161 13 21 32.941 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.43 $Y=3.02 $X2=4.43
+ $Y2=2.77
r162 13 15 49.7577 $w=5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.43 $Y=3.02
+ $X2=4.43 $Y2=3.485
r163 7 19 39.0276 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.05 $Y=1.17 $X2=3.05
+ $Y2=1.42
r164 7 9 45.4775 $w=5e-07 $l=4.25e-07 $layer=POLY_cond $X=3.05 $Y=1.17 $X2=3.05
+ $Y2=0.745
r165 2 30 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.11
+ $Y=3.245 $X2=1.25 $Y2=3.455
r166 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.11
+ $Y=0.655 $X2=1.25 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%SCD 1 3 6 7 9 13 15 16 21 25 30
c67 21 0 1.72602e-20 $X=4.54 $Y=0.745
c68 6 0 7.00078e-20 $X=3.72 $Y=3.015
r69 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.54
+ $Y=1.46 $X2=4.54 $Y2=1.46
r70 21 24 76.5092 $w=5e-07 $l=7.15e-07 $layer=POLY_cond $X=4.54 $Y=0.745
+ $X2=4.54 $Y2=1.46
r71 16 30 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.54 $Y=2.065 $X2=4.54
+ $Y2=1.975
r72 16 30 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=4.54 $Y=1.962
+ $X2=4.54 $Y2=1.975
r73 15 16 10.372 $w=3.28e-07 $l=2.97e-07 $layer=LI1_cond $X=4.54 $Y=1.665
+ $X2=4.54 $Y2=1.962
r74 15 25 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.54 $Y=1.665
+ $X2=4.54 $Y2=1.46
r75 13 29 45.5978 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=3.875 $Y=2.315
+ $X2=3.875 $Y2=2.56
r76 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.875
+ $Y=2.315 $X2=3.875 $Y2=2.315
r77 9 12 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.875 $Y=2.065
+ $X2=3.875 $Y2=2.315
r78 8 9 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.04 $Y=2.065
+ $X2=3.875 $Y2=2.065
r79 7 16 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.375 $Y=2.065
+ $X2=4.54 $Y2=2.065
r80 7 8 20.6414 $w=1.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.375 $Y=2.065
+ $X2=4.04 $Y2=2.065
r81 6 29 108.698 $w=2.6e-07 $l=4.55e-07 $layer=POLY_cond $X=3.84 $Y=3.015
+ $X2=3.84 $Y2=2.56
r82 1 6 39.0276 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.72 $Y=3.265 $X2=3.72
+ $Y2=3.015
r83 1 3 21.208 $w=5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.72 $Y=3.265 $X2=3.72
+ $Y2=3.485
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%CLK 3 7 9 12 13
r35 12 15 48.459 $w=6e-07 $l=5.25e-07 $layer=POLY_cond $X=6.15 $Y=2.015 $X2=6.15
+ $Y2=2.54
r36 12 14 23.9368 $w=6e-07 $l=2.5e-07 $layer=POLY_cond $X=6.15 $Y=2.015 $X2=6.15
+ $Y2=1.765
r37 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.035
+ $Y=2.015 $X2=6.035 $Y2=2.015
r38 9 13 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6.035 $Y=2.405
+ $X2=6.035 $Y2=2.015
r39 7 15 85.6047 $w=5e-07 $l=8e-07 $layer=POLY_cond $X=6.2 $Y=3.34 $X2=6.2
+ $Y2=2.54
r40 3 14 98.9805 $w=5e-07 $l=9.25e-07 $layer=POLY_cond $X=6.2 $Y=0.84 $X2=6.2
+ $Y2=1.765
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%A_1569_126# 1 2 7 9 12 16 18 19 20 22 25
+ 28 31 32 33 35 36 40 41 43 45 49 50 53 54 57 64 68
c187 68 0 1.02319e-19 $X=12.897 $Y=1.395
c188 57 0 9.36316e-20 $X=9.745 $Y=0.84
c189 54 0 3.39237e-20 $X=12.99 $Y=1.56
c190 49 0 6.67328e-20 $X=9.837 $Y=1.01
c191 33 0 1.3651e-19 $X=12.145 $Y=0.35
c192 25 0 2.48877e-20 $X=9.81 $Y=1.44
r193 54 68 15.9063 $w=5.55e-07 $l=1.65e-07 $layer=POLY_cond $X=12.897 $Y=1.56
+ $X2=12.897 $Y2=1.395
r194 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.99
+ $Y=1.56 $X2=12.99 $Y2=1.56
r195 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.52
+ $Y=2.57 $X2=8.52 $Y2=2.57
r196 45 47 3.28743 $w=6.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.255 $Y=2.39
+ $X2=8.255 $Y2=2.57
r197 41 64 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=14.105 $Y=2.39
+ $X2=14.105 $Y2=2.925
r198 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.185
+ $Y=2.39 $X2=14.185 $Y2=2.39
r199 38 40 127.545 $w=1.68e-07 $l=1.955e-06 $layer=LI1_cond $X=14.185 $Y=0.435
+ $X2=14.185 $Y2=2.39
r200 37 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.995 $Y=0.35
+ $X2=12.91 $Y2=0.35
r201 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.1 $Y=0.35
+ $X2=14.185 $Y2=0.435
r202 36 37 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=14.1 $Y=0.35
+ $X2=12.995 $Y2=0.35
r203 35 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.91 $Y=1.475
+ $X2=12.91 $Y2=1.56
r204 34 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.91 $Y=0.435
+ $X2=12.91 $Y2=0.35
r205 34 35 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=12.91 $Y=0.435
+ $X2=12.91 $Y2=1.475
r206 32 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.825 $Y=0.35
+ $X2=12.91 $Y2=0.35
r207 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=12.825 $Y=0.35
+ $X2=12.145 $Y2=0.35
r208 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.06 $Y=0.435
+ $X2=12.145 $Y2=0.35
r209 30 31 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=12.06 $Y=0.435
+ $X2=12.06 $Y2=0.925
r210 29 49 3.11956 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=9.975 $Y=1.01
+ $X2=9.837 $Y2=1.01
r211 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.975 $Y=1.01
+ $X2=12.06 $Y2=0.925
r212 28 29 130.481 $w=1.68e-07 $l=2e-06 $layer=LI1_cond $X=11.975 $Y=1.01
+ $X2=9.975 $Y2=1.01
r213 26 57 64.2035 $w=5e-07 $l=6e-07 $layer=POLY_cond $X=9.745 $Y=1.44 $X2=9.745
+ $Y2=0.84
r214 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.81
+ $Y=1.44 $X2=9.81 $Y2=1.44
r215 23 49 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=9.837 $Y=1.095
+ $X2=9.837 $Y2=1.01
r216 23 25 14.4579 $w=2.73e-07 $l=3.45e-07 $layer=LI1_cond $X=9.837 $Y=1.095
+ $X2=9.837 $Y2=1.44
r217 22 49 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=9.837 $Y=0.925
+ $X2=9.837 $Y2=1.01
r218 21 22 20.5344 $w=2.73e-07 $l=4.9e-07 $layer=LI1_cond $X=9.837 $Y=0.435
+ $X2=9.837 $Y2=0.925
r219 19 21 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=9.7 $Y=0.35
+ $X2=9.837 $Y2=0.435
r220 19 20 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=9.7 $Y=0.35
+ $X2=8.15 $Y2=0.35
r221 18 45 8.15664 $w=6.68e-07 $l=2.99339e-07 $layer=LI1_cond $X=8.027 $Y=2.225
+ $X2=8.255 $Y2=2.39
r222 18 43 57.8573 $w=2.43e-07 $l=1.23e-06 $layer=LI1_cond $X=8.027 $Y=2.225
+ $X2=8.027 $Y2=0.995
r223 14 43 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=8.025 $Y=0.87
+ $X2=8.025 $Y2=0.995
r224 14 16 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=8.025 $Y=0.87
+ $X2=8.025 $Y2=0.83
r225 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.025 $Y=0.435
+ $X2=8.15 $Y2=0.35
r226 13 16 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=8.025 $Y=0.435
+ $X2=8.025 $Y2=0.83
r227 12 68 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=12.87 $Y=0.91
+ $X2=12.87 $Y2=1.395
r228 7 48 47.5716 $w=6.67e-07 $l=6.8815e-07 $layer=POLY_cond $X=8.83 $Y=3.185
+ $X2=8.675 $Y2=2.57
r229 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.83 $Y=3.185 $X2=8.83
+ $Y2=3.505
r230 2 45 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.93
+ $Y=2.245 $X2=8.07 $Y2=2.39
r231 1 16 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=7.845
+ $Y=0.63 $X2=7.985 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%A_1290_126# 1 2 9 12 14 16 18 20 23 27 29
+ 30 33 35 39 43 45 47 50 51 52 55 58 60 66 67 71 75 76 85
c216 55 0 3.39237e-20 $X=13.055 $Y=2.26
c217 23 0 7.48103e-20 $X=9.61 $Y=3.505
c218 16 0 9.16205e-20 $X=8.965 $Y=1.125
r219 75 76 21.4018 $w=5.85e-07 $l=2.2e-07 $layer=POLY_cond $X=7.637 $Y=1.345
+ $X2=7.637 $Y2=1.125
r220 71 73 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.21 $Y=1.96
+ $X2=12.21 $Y2=2.26
r221 67 81 7.02564 $w=4.95e-07 $l=6.5e-08 $layer=POLY_cond $X=9.675 $Y=2.232
+ $X2=9.61 $Y2=2.232
r222 66 69 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=9.675 $Y=2.17
+ $X2=9.675 $Y2=2.4
r223 66 67 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.675
+ $Y=2.17 $X2=9.675 $Y2=2.17
r224 61 78 25.5174 $w=5.85e-07 $l=2.65e-07 $layer=POLY_cond $X=7.637 $Y=1.51
+ $X2=7.637 $Y2=1.775
r225 61 75 15.0906 $w=5.85e-07 $l=1.65e-07 $layer=POLY_cond $X=7.637 $Y=1.51
+ $X2=7.637 $Y2=1.345
r226 60 63 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.53 $Y=1.51 $X2=7.53
+ $Y2=1.59
r227 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.53
+ $Y=1.51 $X2=7.53 $Y2=1.51
r228 56 85 14.1765 $w=5.27e-07 $l=1.55e-07 $layer=POLY_cond $X=13.055 $Y=2.16
+ $X2=13.21 $Y2=2.16
r229 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.055
+ $Y=2.26 $X2=13.055 $Y2=2.26
r230 53 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.295 $Y=2.26
+ $X2=12.21 $Y2=2.26
r231 53 55 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=12.295 $Y=2.26
+ $X2=13.055 $Y2=2.26
r232 51 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.125 $Y=1.96
+ $X2=12.21 $Y2=1.96
r233 51 52 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=12.125 $Y=1.96
+ $X2=11.595 $Y2=1.96
r234 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.51 $Y=2.045
+ $X2=11.595 $Y2=1.96
r235 49 50 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=11.51 $Y=2.045
+ $X2=11.51 $Y2=2.315
r236 48 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.84 $Y=2.4
+ $X2=9.675 $Y2=2.4
r237 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.425 $Y=2.4
+ $X2=11.51 $Y2=2.315
r238 47 48 103.406 $w=1.68e-07 $l=1.585e-06 $layer=LI1_cond $X=11.425 $Y=2.4
+ $X2=9.84 $Y2=2.4
r239 46 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.675 $Y=1.59
+ $X2=6.59 $Y2=1.59
r240 45 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.365 $Y=1.59
+ $X2=7.53 $Y2=1.59
r241 45 46 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.365 $Y=1.59
+ $X2=6.675 $Y2=1.59
r242 41 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.59 $Y=1.675
+ $X2=6.59 $Y2=1.59
r243 41 43 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=6.59 $Y=1.675
+ $X2=6.59 $Y2=3.19
r244 37 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.59 $Y=1.505
+ $X2=6.59 $Y2=1.59
r245 37 39 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=6.59 $Y=1.505
+ $X2=6.59 $Y2=0.83
r246 33 36 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=13.745 $Y=0.745
+ $X2=13.745 $Y2=1.085
r247 30 85 47.2854 $w=5.27e-07 $l=6.97864e-07 $layer=POLY_cond $X=13.727
+ $Y=1.735 $X2=13.21 $Y2=2.16
r248 29 36 27.0046 $w=5.35e-07 $l=2.67e-07 $layer=POLY_cond $X=13.727 $Y=1.352
+ $X2=13.727 $Y2=1.085
r249 29 30 38.3021 $w=5.35e-07 $l=3.83e-07 $layer=POLY_cond $X=13.727 $Y=1.352
+ $X2=13.727 $Y2=1.735
r250 25 85 4.08967 $w=5e-07 $l=4.25e-07 $layer=POLY_cond $X=13.21 $Y=2.585
+ $X2=13.21 $Y2=2.16
r251 25 27 67.4137 $w=5e-07 $l=6.3e-07 $layer=POLY_cond $X=13.21 $Y=2.585
+ $X2=13.21 $Y2=3.215
r252 21 81 2.58818 $w=5e-07 $l=2.48e-07 $layer=POLY_cond $X=9.61 $Y=2.48
+ $X2=9.61 $Y2=2.232
r253 21 23 109.681 $w=5e-07 $l=1.025e-06 $layer=POLY_cond $X=9.61 $Y=2.48
+ $X2=9.61 $Y2=3.505
r254 20 81 55.1242 $w=4.95e-07 $l=5.1e-07 $layer=POLY_cond $X=9.1 $Y=2.232
+ $X2=9.61 $Y2=2.232
r255 19 35 20.6049 $w=4.35e-07 $l=2.6533e-07 $layer=POLY_cond $X=9.1 $Y=1.565
+ $X2=9 $Y2=1.345
r256 19 20 65.5021 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=9.1 $Y=1.565
+ $X2=9.1 $Y2=1.985
r257 16 35 20.6049 $w=4.35e-07 $l=2.36854e-07 $layer=POLY_cond $X=8.965 $Y=1.125
+ $X2=9 $Y2=1.345
r258 16 18 27.474 $w=5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.965 $Y=1.125
+ $X2=8.965 $Y2=0.84
r259 15 75 9.51117 $w=4.4e-07 $l=2.93e-07 $layer=POLY_cond $X=7.93 $Y=1.345
+ $X2=7.637 $Y2=1.345
r260 14 35 5.14175 $w=4.4e-07 $l=2.85e-07 $layer=POLY_cond $X=8.715 $Y=1.345
+ $X2=9 $Y2=1.345
r261 14 15 99.2229 $w=4.4e-07 $l=7.85e-07 $layer=POLY_cond $X=8.715 $Y=1.345
+ $X2=7.93 $Y2=1.345
r262 12 78 90.42 $w=5e-07 $l=8.45e-07 $layer=POLY_cond $X=7.68 $Y=2.62 $X2=7.68
+ $Y2=1.775
r263 9 76 27.474 $w=5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.595 $Y=0.84
+ $X2=7.595 $Y2=1.125
r264 2 43 600 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_PDIFF $count=1 $X=6.45
+ $Y=2.965 $X2=6.59 $Y2=3.19
r265 1 39 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=6.45
+ $Y=0.63 $X2=6.59 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%A_2014_537# 1 2 9 12 13 15 18 22 25 26 27
+ 30 34 35 37 39 41 43
c122 43 0 7.25359e-20 $X=10.455 $Y=0.84
r123 40 43 64.2035 $w=5e-07 $l=6e-07 $layer=POLY_cond $X=10.455 $Y=1.44
+ $X2=10.455 $Y2=0.84
r124 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.39
+ $Y=1.44 $X2=10.39 $Y2=1.44
r125 36 37 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=13.485 $Y=1.995
+ $X2=13.485 $Y2=2.525
r126 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.4 $Y=2.61
+ $X2=13.485 $Y2=2.525
r127 34 35 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=13.4 $Y=2.61
+ $X2=12.985 $Y2=2.61
r128 30 32 34.5733 $w=2.48e-07 $l=7.5e-07 $layer=LI1_cond $X=12.86 $Y=2.84
+ $X2=12.86 $Y2=3.59
r129 28 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.86 $Y=2.695
+ $X2=12.985 $Y2=2.61
r130 28 30 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=12.86 $Y=2.695
+ $X2=12.86 $Y2=2.84
r131 26 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.4 $Y=1.91
+ $X2=13.485 $Y2=1.995
r132 26 27 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=13.4 $Y=1.91
+ $X2=12.645 $Y2=1.91
r133 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.56 $Y=1.825
+ $X2=12.645 $Y2=1.91
r134 24 41 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=12.56 $Y=1.445
+ $X2=12.48 $Y2=1.36
r135 24 25 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=12.56 $Y=1.445
+ $X2=12.56 $Y2=1.825
r136 20 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.48 $Y=1.275
+ $X2=12.48 $Y2=1.36
r137 20 22 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=12.48 $Y=1.275
+ $X2=12.48 $Y2=0.7
r138 19 39 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=10.505 $Y=1.36
+ $X2=10.365 $Y2=1.36
r139 18 41 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.315 $Y=1.36
+ $X2=12.48 $Y2=1.36
r140 18 19 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=12.315 $Y=1.36
+ $X2=10.505 $Y2=1.36
r141 14 40 29.4266 $w=5e-07 $l=2.75e-07 $layer=POLY_cond $X=10.455 $Y=1.715
+ $X2=10.455 $Y2=1.44
r142 14 15 27.7985 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=10.455 $Y=1.715
+ $X2=10.455 $Y2=1.965
r143 12 13 54.55 $w=5e-07 $l=5e-07 $layer=POLY_cond $X=10.355 $Y=2.685
+ $X2=10.355 $Y2=3.185
r144 12 15 92.0531 $w=4.35e-07 $l=7.2e-07 $layer=POLY_cond $X=10.422 $Y=2.685
+ $X2=10.422 $Y2=1.965
r145 9 13 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.32 $Y=3.505
+ $X2=10.32 $Y2=3.185
r146 2 32 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=12.68
+ $Y=2.715 $X2=12.82 $Y2=3.59
r147 2 30 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=12.68
+ $Y=2.715 $X2=12.82 $Y2=2.84
r148 1 22 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=12.34
+ $Y=0.535 $X2=12.48 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%RESET_B 3 7 8 9 12 14 16 19 22 25 27 28 31
+ 32 33 34 43 48 51 54 56 62 63
c213 51 0 1.3651e-19 $X=11.165 $Y=0.84
c214 28 0 1.15308e-20 $X=15.6 $Y=2.035
c215 25 0 1.54595e-19 $X=15.24 $Y=1.765
c216 19 0 1.78387e-19 $X=5.292 $Y=3.165
r217 62 65 9.69479 $w=6e-07 $l=9.5e-08 $layer=POLY_cond $X=5.37 $Y=1.46 $X2=5.37
+ $Y2=1.555
r218 62 64 26.1661 $w=6e-07 $l=2.75e-07 $layer=POLY_cond $X=5.37 $Y=1.46
+ $X2=5.37 $Y2=1.185
r219 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.4
+ $Y=1.46 $X2=5.4 $Y2=1.46
r220 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=15.175
+ $Y=1.51 $X2=15.175 $Y2=1.51
r221 56 59 81.8595 $w=5e-07 $l=7.65e-07 $layer=POLY_cond $X=15.24 $Y=0.745
+ $X2=15.24 $Y2=1.51
r222 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.08
+ $Y=1.71 $X2=11.08 $Y2=1.71
r223 51 53 93.0951 $w=5e-07 $l=8.7e-07 $layer=POLY_cond $X=11.165 $Y=0.84
+ $X2=11.165 $Y2=1.71
r224 49 63 9.79577 $w=3.98e-07 $l=3.4e-07 $layer=LI1_cond $X=5.435 $Y=1.8
+ $X2=5.435 $Y2=1.46
r225 48 65 25.4529 $w=5.15e-07 $l=2.45e-07 $layer=POLY_cond $X=5.327 $Y=1.8
+ $X2=5.327 $Y2=1.555
r226 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.4
+ $Y=1.8 $X2=5.4 $Y2=1.8
r227 41 54 6.5667 $w=5.08e-07 $l=2.8e-07 $layer=LI1_cond $X=10.8 $Y=1.88
+ $X2=11.08 $Y2=1.88
r228 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r229 37 49 6.7706 $w=3.98e-07 $l=2.35e-07 $layer=LI1_cond $X=5.435 $Y=2.035
+ $X2=5.435 $Y2=1.8
r230 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r231 34 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.945 $Y=2.035
+ $X2=10.8 $Y2=2.035
r232 33 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.975 $Y=2.035
+ $X2=15.12 $Y2=2.035
r233 33 34 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=14.975 $Y=2.035
+ $X2=10.945 $Y2=2.035
r234 32 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r235 31 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r236 31 32 6.17573 $w=1.4e-07 $l=4.99e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=5.665 $Y2=2.035
r237 28 60 7.31415 $w=6.93e-07 $l=4.25e-07 $layer=LI1_cond $X=15.6 $Y=1.772
+ $X2=15.175 $Y2=1.772
r238 27 60 0.946537 $w=6.93e-07 $l=5.5e-08 $layer=LI1_cond $X=15.12 $Y=1.772
+ $X2=15.175 $Y2=1.772
r239 27 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=2.035
+ $X2=15.12 $Y2=2.035
r240 25 59 27.2865 $w=5e-07 $l=2.55e-07 $layer=POLY_cond $X=15.24 $Y=1.765
+ $X2=15.24 $Y2=1.51
r241 25 26 37.442 $w=4.57e-07 $l=5.70526e-07 $layer=POLY_cond $X=15.24 $Y=1.765
+ $X2=15.595 $Y2=2.185
r242 23 51 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=11.165 $Y=0.29
+ $X2=11.165 $Y2=0.84
r243 21 53 102.191 $w=5e-07 $l=9.55e-07 $layer=POLY_cond $X=11.165 $Y=2.665
+ $X2=11.165 $Y2=1.71
r244 21 22 47.3477 $w=5.65e-07 $l=5e-07 $layer=POLY_cond $X=11.132 $Y=2.665
+ $X2=11.132 $Y2=3.165
r245 18 48 89.8642 $w=5.15e-07 $l=8.65e-07 $layer=POLY_cond $X=5.327 $Y=2.665
+ $X2=5.327 $Y2=1.8
r246 18 19 51.9446 $w=5.15e-07 $l=5e-07 $layer=POLY_cond $X=5.292 $Y=2.665
+ $X2=5.292 $Y2=3.165
r247 14 26 0.633894 $w=5e-07 $l=4.2e-07 $layer=POLY_cond $X=15.595 $Y=2.605
+ $X2=15.595 $Y2=2.185
r248 14 16 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=15.595 $Y=2.605
+ $X2=15.595 $Y2=2.925
r249 12 22 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=11.1 $Y=3.505 $X2=11.1
+ $Y2=3.165
r250 8 23 38.6381 $w=1.5e-07 $l=2.85044e-07 $layer=POLY_cond $X=10.915 $Y=0.215
+ $X2=11.165 $Y2=0.29
r251 8 9 2689.46 $w=1.5e-07 $l=5.245e-06 $layer=POLY_cond $X=10.915 $Y=0.215
+ $X2=5.67 $Y2=0.215
r252 7 64 36.917 $w=5e-07 $l=3.45e-07 $layer=POLY_cond $X=5.42 $Y=0.84 $X2=5.42
+ $Y2=1.185
r253 4 9 38.6381 $w=1.5e-07 $l=2.85044e-07 $layer=POLY_cond $X=5.42 $Y=0.29
+ $X2=5.67 $Y2=0.215
r254 4 7 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.42 $Y=0.29 $X2=5.42
+ $Y2=0.84
r255 3 19 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.25 $Y=3.485 $X2=5.25
+ $Y2=3.165
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%A_1816_659# 1 2 3 12 16 19 22 24 26 28 32
+ 38 40 45
c120 38 0 7.25359e-20 $X=9.355 $Y=0.85
r121 44 45 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=12.09 $Y=2.335
+ $X2=12.43 $Y2=2.335
r122 35 38 4.09421 $w=3.78e-07 $l=1.35e-07 $layer=LI1_cond $X=9.22 $Y=0.805
+ $X2=9.355 $Y2=0.805
r123 33 44 24.6114 $w=5e-07 $l=2.3e-07 $layer=POLY_cond $X=11.86 $Y=2.335
+ $X2=12.09 $Y2=2.335
r124 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.86
+ $Y=2.39 $X2=11.86 $Y2=2.39
r125 30 41 13.588 $w=5.2e-07 $l=4.22788e-07 $layer=LI1_cond $X=11.86 $Y=2.665
+ $X2=11.635 $Y2=2.99
r126 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.86 $Y=2.665
+ $X2=11.86 $Y2=2.39
r127 26 41 2.24855 $w=5.2e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.55 $Y=3.075
+ $X2=11.635 $Y2=2.99
r128 26 28 11.4292 $w=4.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.55 $Y=3.075
+ $X2=11.55 $Y2=3.505
r129 25 40 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.385 $Y=2.99
+ $X2=9.26 $Y2=2.99
r130 24 41 7.40362 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=11.325 $Y=2.99
+ $X2=11.635 $Y2=2.99
r131 24 25 126.567 $w=1.68e-07 $l=1.94e-06 $layer=LI1_cond $X=11.325 $Y=2.99
+ $X2=9.385 $Y2=2.99
r132 20 40 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=9.26 $Y=3.075
+ $X2=9.26 $Y2=2.99
r133 20 22 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.26 $Y=3.075
+ $X2=9.26 $Y2=3.505
r134 19 40 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=9.22 $Y=2.905
+ $X2=9.26 $Y2=2.99
r135 18 35 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.22 $Y=0.995
+ $X2=9.22 $Y2=0.805
r136 18 19 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=9.22 $Y=0.995
+ $X2=9.22 $Y2=2.905
r137 14 45 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=12.43 $Y=2.585
+ $X2=12.43 $Y2=2.335
r138 14 16 67.4137 $w=5e-07 $l=6.3e-07 $layer=POLY_cond $X=12.43 $Y=2.585
+ $X2=12.43 $Y2=3.215
r139 10 44 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=12.09 $Y=2.085
+ $X2=12.09 $Y2=2.335
r140 10 12 125.732 $w=5e-07 $l=1.175e-06 $layer=POLY_cond $X=12.09 $Y=2.085
+ $X2=12.09 $Y2=0.91
r141 3 28 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.35
+ $Y=3.295 $X2=11.49 $Y2=3.505
r142 2 22 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=9.08
+ $Y=3.295 $X2=9.22 $Y2=3.505
r143 1 38 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=9.215
+ $Y=0.63 $X2=9.355 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%A_2841_81# 1 2 9 14 15 16 17 20 24 27 28
+ 29 31 32 36 39 40
c96 16 0 1.52211e-19 $X=14.492 $Y=1.565
r97 34 36 3.63929 $w=3.78e-07 $l=1.2e-07 $layer=LI1_cond $X=16.34 $Y=0.705
+ $X2=16.46 $Y2=0.705
r98 30 36 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=16.46 $Y=0.895
+ $X2=16.46 $Y2=0.705
r99 30 31 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=16.46 $Y=0.895
+ $X2=16.46 $Y2=1.835
r100 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=16.375 $Y=1.92
+ $X2=16.46 $Y2=1.835
r101 28 29 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=16.375 $Y=1.92
+ $X2=16.15 $Y2=1.92
r102 27 32 4.85493 $w=2.1e-07 $l=1.15278e-07 $layer=LI1_cond $X=16.065 $Y=2.3
+ $X2=16.025 $Y2=2.397
r103 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=16.065 $Y=2.005
+ $X2=16.15 $Y2=1.92
r104 26 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=16.065 $Y=2.005
+ $X2=16.065 $Y2=2.3
r105 22 32 4.85493 $w=2.1e-07 $l=9.8e-08 $layer=LI1_cond $X=16.025 $Y=2.495
+ $X2=16.025 $Y2=2.397
r106 22 24 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=16.025 $Y=2.495
+ $X2=16.025 $Y2=2.925
r107 20 40 21.1989 $w=5.65e-07 $l=2.15e-07 $layer=POLY_cond $X=14.847 $Y=2.39
+ $X2=14.847 $Y2=2.605
r108 20 39 37.0454 $w=5.65e-07 $l=1.65e-07 $layer=POLY_cond $X=14.847 $Y=2.39
+ $X2=14.847 $Y2=2.225
r109 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.965
+ $Y=2.39 $X2=14.965 $Y2=2.39
r110 17 32 1.61074 $w=1.95e-07 $l=1.25e-07 $layer=LI1_cond $X=15.9 $Y=2.397
+ $X2=16.025 $Y2=2.397
r111 17 19 53.1795 $w=1.93e-07 $l=9.35e-07 $layer=LI1_cond $X=15.9 $Y=2.397
+ $X2=14.965 $Y2=2.397
r112 16 39 196.992 $w=2.15e-07 $l=6.6e-07 $layer=POLY_cond $X=14.672 $Y=1.565
+ $X2=14.672 $Y2=2.225
r113 15 16 71.2322 $w=5e-07 $l=5e-07 $layer=POLY_cond $X=14.492 $Y=1.065
+ $X2=14.492 $Y2=1.565
r114 14 40 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=14.815 $Y=2.925
+ $X2=14.815 $Y2=2.605
r115 9 15 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=14.455 $Y=0.745
+ $X2=14.455 $Y2=1.065
r116 2 24 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=15.845
+ $Y=2.715 $X2=15.985 $Y2=2.925
r117 1 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=16.2
+ $Y=0.535 $X2=16.34 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%A_2624_107# 1 2 7 9 12 16 18 20 21 22 25
+ 29 31 32 34 36 40 43 44 47 48 49 55 57
c163 36 0 1.52211e-19 $X=13.75 $Y=1.21
c164 32 0 1.02319e-19 $X=13.3 $Y=1.125
c165 12 0 1.15308e-20 $X=16.375 $Y=2.925
r166 61 62 68.9134 $w=6.12e-07 $l=8.75e-07 $layer=POLY_cond $X=16.375 $Y=1.492
+ $X2=17.25 $Y2=1.492
r167 58 61 27.1716 $w=6.12e-07 $l=3.45e-07 $layer=POLY_cond $X=16.03 $Y=1.492
+ $X2=16.375 $Y2=1.492
r168 58 59 6.30065 $w=6.12e-07 $l=8e-08 $layer=POLY_cond $X=16.03 $Y=1.492
+ $X2=15.95 $Y2=1.492
r169 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=16.03
+ $Y=1.23 $X2=16.03 $Y2=1.23
r170 48 57 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.865 $Y=1.16
+ $X2=16.03 $Y2=1.16
r171 48 49 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=15.865 $Y=1.16
+ $X2=14.62 $Y2=1.16
r172 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.535 $Y=1.245
+ $X2=14.62 $Y2=1.16
r173 46 47 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=14.535 $Y=1.245
+ $X2=14.535 $Y2=2.875
r174 45 55 2.76166 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=13.92 $Y=2.96
+ $X2=13.677 $Y2=2.96
r175 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.45 $Y=2.96
+ $X2=14.535 $Y2=2.875
r176 44 45 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=14.45 $Y=2.96
+ $X2=13.92 $Y2=2.96
r177 43 55 3.70735 $w=2.5e-07 $l=1.95944e-07 $layer=LI1_cond $X=13.835 $Y=2.875
+ $X2=13.677 $Y2=2.96
r178 42 43 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=13.835 $Y=1.295
+ $X2=13.835 $Y2=2.875
r179 38 55 3.70735 $w=2.5e-07 $l=1.17346e-07 $layer=LI1_cond $X=13.6 $Y=3.045
+ $X2=13.677 $Y2=2.96
r180 38 40 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=13.6 $Y=3.045
+ $X2=13.6 $Y2=3.59
r181 37 53 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.425 $Y=1.21
+ $X2=13.3 $Y2=1.21
r182 36 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.75 $Y=1.21
+ $X2=13.835 $Y2=1.295
r183 36 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=13.75 $Y=1.21
+ $X2=13.425 $Y2=1.21
r184 32 53 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.3 $Y=1.125
+ $X2=13.3 $Y2=1.21
r185 32 34 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=13.3 $Y=1.125
+ $X2=13.3 $Y2=0.78
r186 27 31 21.2518 $w=5e-07 $l=3.5242e-07 $layer=POLY_cond $X=18.61 $Y=1.395
+ $X2=18.595 $Y2=1.74
r187 27 29 51.3628 $w=5e-07 $l=4.8e-07 $layer=POLY_cond $X=18.61 $Y=1.395
+ $X2=18.61 $Y2=0.915
r188 23 31 21.2518 $w=5e-07 $l=3.5242e-07 $layer=POLY_cond $X=18.58 $Y=2.085
+ $X2=18.595 $Y2=1.74
r189 23 25 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=18.58 $Y=2.085
+ $X2=18.58 $Y2=2.59
r190 21 31 4.61246 $w=5.25e-07 $l=3.03677e-07 $layer=POLY_cond $X=18.33 $Y=1.657
+ $X2=18.595 $Y2=1.74
r191 21 22 81.5283 $w=5.25e-07 $l=8e-07 $layer=POLY_cond $X=18.33 $Y=1.657
+ $X2=17.53 $Y2=1.657
r192 18 22 20.7987 $w=6.12e-07 $l=3.22102e-07 $layer=POLY_cond $X=17.28 $Y=1.492
+ $X2=17.53 $Y2=1.657
r193 18 62 2.36275 $w=6.12e-07 $l=3e-08 $layer=POLY_cond $X=17.28 $Y=1.492
+ $X2=17.25 $Y2=1.492
r194 18 20 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=17.28 $Y=1.395
+ $X2=17.28 $Y2=0.91
r195 14 62 7.59805 $w=5e-07 $l=4.28e-07 $layer=POLY_cond $X=17.25 $Y=1.92
+ $X2=17.25 $Y2=1.492
r196 14 16 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=17.25 $Y=1.92
+ $X2=17.25 $Y2=2.8
r197 10 61 7.59805 $w=5e-07 $l=4.28e-07 $layer=POLY_cond $X=16.375 $Y=1.92
+ $X2=16.375 $Y2=1.492
r198 10 12 107.541 $w=5e-07 $l=1.005e-06 $layer=POLY_cond $X=16.375 $Y=1.92
+ $X2=16.375 $Y2=2.925
r199 7 59 7.59805 $w=5e-07 $l=4.27e-07 $layer=POLY_cond $X=15.95 $Y=1.065
+ $X2=15.95 $Y2=1.492
r200 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=15.95 $Y=1.065 $X2=15.95
+ $Y2=0.745
r201 2 55 600 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_PDIFF $count=1 $X=13.46
+ $Y=2.715 $X2=13.6 $Y2=2.96
r202 2 40 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=13.46
+ $Y=2.715 $X2=13.6 $Y2=3.59
r203 1 53 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=13.12
+ $Y=0.535 $X2=13.26 $Y2=1.13
r204 1 34 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=13.12
+ $Y=0.535 $X2=13.26 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%A_3613_443# 1 2 9 13 17 21 25 26 28
r45 26 31 25.9337 $w=5.65e-07 $l=2.65e-07 $layer=POLY_cond $X=19.452 $Y=1.82
+ $X2=19.452 $Y2=2.085
r46 26 30 23.0928 $w=5.65e-07 $l=2.35e-07 $layer=POLY_cond $X=19.452 $Y=1.82
+ $X2=19.452 $Y2=1.585
r47 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=19.355
+ $Y=1.82 $X2=19.355 $Y2=1.82
r48 23 28 1.50311 $w=3.3e-07 $l=1.8e-07 $layer=LI1_cond $X=18.385 $Y=1.82
+ $X2=18.205 $Y2=1.82
r49 23 25 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=18.385 $Y=1.82
+ $X2=19.355 $Y2=1.82
r50 19 28 4.97762 $w=3.45e-07 $l=1.72337e-07 $layer=LI1_cond $X=18.19 $Y=1.985
+ $X2=18.205 $Y2=1.82
r51 19 21 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=18.19 $Y=1.985
+ $X2=18.19 $Y2=2.36
r52 15 28 4.97762 $w=3.45e-07 $l=1.65e-07 $layer=LI1_cond $X=18.205 $Y=1.655
+ $X2=18.205 $Y2=1.82
r53 15 17 23.6891 $w=3.58e-07 $l=7.4e-07 $layer=LI1_cond $X=18.205 $Y=1.655
+ $X2=18.205 $Y2=0.915
r54 13 30 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=19.485 $Y=1.08
+ $X2=19.485 $Y2=1.585
r55 9 31 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=19.475 $Y=2.965
+ $X2=19.475 $Y2=2.085
r56 2 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=18.065
+ $Y=2.215 $X2=18.19 $Y2=2.36
r57 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=18.095
+ $Y=0.705 $X2=18.22 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%VPWR 1 2 3 4 5 6 7 8 9 28 31 44 53 58 69
+ 74 81 90 103 111
c158 81 0 1.54595e-19 $X=15.205 $Y=2.925
r159 109 111 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=18.65 $Y=3.63
+ $X2=19.37 $Y2=3.63
r160 108 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=19.37 $Y=3.59
+ $X2=19.37 $Y2=3.59
r161 108 109 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=18.65 $Y=3.59
+ $X2=18.65 $Y2=3.59
r162 106 108 5.32947 $w=9.48e-07 $l=4.15e-07 $layer=LI1_cond $X=19.01 $Y=3.175
+ $X2=19.01 $Y2=3.59
r163 103 106 10.7232 $w=9.48e-07 $l=8.35e-07 $layer=LI1_cond $X=19.01 $Y=2.34
+ $X2=19.01 $Y2=3.175
r164 100 109 0.575858 $w=3.7e-07 $l=1.5e-06 $layer=MET1_cond $X=17.15 $Y=3.63
+ $X2=18.65 $Y2=3.63
r165 98 100 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=16.43 $Y=3.63
+ $X2=17.15 $Y2=3.63
r166 97 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.15 $Y=3.59
+ $X2=17.15 $Y2=3.59
r167 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.43 $Y=3.59
+ $X2=16.43 $Y2=3.59
r168 95 97 2.44 $w=9.23e-07 $l=1.85e-07 $layer=LI1_cond $X=16.792 $Y=3.405
+ $X2=16.792 $Y2=3.59
r169 93 95 4.94595 $w=9.23e-07 $l=3.75e-07 $layer=LI1_cond $X=16.792 $Y=3.03
+ $X2=16.792 $Y2=3.405
r170 90 93 10.0238 $w=9.23e-07 $l=7.6e-07 $layer=LI1_cond $X=16.792 $Y=2.27
+ $X2=16.792 $Y2=3.03
r171 87 98 0.310963 $w=3.7e-07 $l=8.1e-07 $layer=MET1_cond $X=15.62 $Y=3.63
+ $X2=16.43 $Y2=3.63
r172 85 87 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=14.9 $Y=3.63
+ $X2=15.62 $Y2=3.63
r173 84 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.62 $Y=3.59
+ $X2=15.62 $Y2=3.59
r174 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.9 $Y=3.59
+ $X2=14.9 $Y2=3.59
r175 81 84 8.81848 $w=9.18e-07 $l=6.65e-07 $layer=LI1_cond $X=15.26 $Y=2.925
+ $X2=15.26 $Y2=3.59
r176 78 85 0.948246 $w=3.7e-07 $l=2.47e-06 $layer=MET1_cond $X=12.43 $Y=3.63
+ $X2=14.9 $Y2=3.63
r177 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.43 $Y=3.59
+ $X2=12.43 $Y2=3.59
r178 74 77 8.31173 $w=5.88e-07 $l=4.1e-07 $layer=LI1_cond $X=12.25 $Y=3.18
+ $X2=12.25 $Y2=3.59
r179 71 78 0.641122 $w=3.7e-07 $l=1.67e-06 $layer=MET1_cond $X=10.76 $Y=3.63
+ $X2=12.43 $Y2=3.63
r180 69 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.76 $Y=3.59
+ $X2=10.76 $Y2=3.59
r181 65 69 16.0275 $w=4.98e-07 $l=6.7e-07 $layer=LI1_cond $X=10.04 $Y=3.505
+ $X2=10.71 $Y2=3.505
r182 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.29 $Y=3.59
+ $X2=7.29 $Y2=3.59
r183 58 61 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=7.29 $Y=2.37
+ $X2=7.29 $Y2=3.59
r184 55 62 0.537468 $w=3.7e-07 $l=1.4e-06 $layer=MET1_cond $X=5.89 $Y=3.63
+ $X2=7.29 $Y2=3.63
r185 53 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.89 $Y=3.59
+ $X2=5.89 $Y2=3.59
r186 50 55 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.17 $Y=3.63
+ $X2=5.89 $Y2=3.63
r187 49 53 18.9119 $w=3.88e-07 $l=6.4e-07 $layer=LI1_cond $X=5.17 $Y=3.56
+ $X2=5.81 $Y2=3.56
r188 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.17 $Y=3.59
+ $X2=5.17 $Y2=3.59
r189 46 50 0.687191 $w=3.7e-07 $l=1.79e-06 $layer=MET1_cond $X=3.38 $Y=3.63
+ $X2=5.17 $Y2=3.63
r190 44 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.38 $Y=3.59
+ $X2=3.38 $Y2=3.59
r191 41 46 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.66 $Y=3.63
+ $X2=3.38 $Y2=3.63
r192 40 44 20.8686 $w=3.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.66 $Y=3.55
+ $X2=3.33 $Y2=3.55
r193 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.66 $Y=3.59
+ $X2=2.66 $Y2=3.59
r194 37 41 0.675673 $w=3.7e-07 $l=1.76e-06 $layer=MET1_cond $X=0.9 $Y=3.63
+ $X2=2.66 $Y2=3.63
r195 35 37 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.18 $Y=3.63
+ $X2=0.9 $Y2=3.63
r196 34 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.9 $Y=3.59
+ $X2=0.9 $Y2=3.59
r197 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.18 $Y=3.59
+ $X2=0.18 $Y2=3.59
r198 31 34 1.84022 $w=8.93e-07 $l=1.35e-07 $layer=LI1_cond $X=0.537 $Y=3.455
+ $X2=0.537 $Y2=3.59
r199 28 71 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.04 $Y=3.63
+ $X2=10.76 $Y2=3.63
r200 28 62 1.05574 $w=3.7e-07 $l=2.75e-06 $layer=MET1_cond $X=10.04 $Y=3.63
+ $X2=7.29 $Y2=3.63
r201 28 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.04 $Y=3.59
+ $X2=10.04 $Y2=3.59
r202 9 106 300 $w=1.7e-07 $l=1.08e-06 $layer=licon1_PDIFF $count=2 $X=18.83
+ $Y=2.215 $X2=19.085 $Y2=3.175
r203 9 103 300 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=2 $X=18.83
+ $Y=2.215 $X2=19.085 $Y2=2.34
r204 8 95 600 $w=1.7e-07 $l=7.98906e-07 $layer=licon1_PDIFF $count=1 $X=16.625
+ $Y=2.715 $X2=16.86 $Y2=3.405
r205 8 93 600 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=1 $X=16.625
+ $Y=2.715 $X2=16.86 $Y2=3.03
r206 8 90 300 $w=1.7e-07 $l=5.50091e-07 $layer=licon1_PDIFF $count=2 $X=16.625
+ $Y=2.715 $X2=16.86 $Y2=2.27
r207 7 81 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=15.065
+ $Y=2.715 $X2=15.205 $Y2=2.925
r208 6 74 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=11.915
+ $Y=2.715 $X2=12.04 $Y2=3.18
r209 5 69 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=10.57
+ $Y=3.295 $X2=10.71 $Y2=3.505
r210 4 58 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=7.145
+ $Y=2.245 $X2=7.29 $Y2=2.37
r211 3 53 600 $w=1.7e-07 $l=4.14789e-07 $layer=licon1_PDIFF $count=1 $X=5.5
+ $Y=3.275 $X2=5.81 $Y2=3.52
r212 2 44 600 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=3.275 $X2=3.33 $Y2=3.51
r213 1 31 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=3.245 $X2=0.47 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%A_339_655# 1 2 3 4 5 16 17 18 22 25 26 29
+ 30 31 33 34 35 37 38 39 40 43 48 52 53 61
c176 61 0 9.36316e-20 $X=8.87 $Y=0.805
c177 40 0 7.48103e-20 $X=8.785 $Y=3.34
c178 18 0 8.22034e-20 $X=4.885 $Y=1.01
r179 59 61 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=8.575 $Y=0.805
+ $X2=8.87 $Y2=0.805
r180 53 56 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.44 $Y=3.34
+ $X2=8.44 $Y2=3.505
r181 48 50 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.44 $Y=0.765
+ $X2=3.44 $Y2=1.01
r182 42 61 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.87 $Y=0.995
+ $X2=8.87 $Y2=0.805
r183 42 43 147.444 $w=1.68e-07 $l=2.26e-06 $layer=LI1_cond $X=8.87 $Y=0.995
+ $X2=8.87 $Y2=3.255
r184 41 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.605 $Y=3.34
+ $X2=8.44 $Y2=3.34
r185 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.785 $Y=3.34
+ $X2=8.87 $Y2=3.255
r186 40 41 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.785 $Y=3.34
+ $X2=8.605 $Y2=3.34
r187 38 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.275 $Y=3.34
+ $X2=8.44 $Y2=3.34
r188 38 39 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=8.275 $Y=3.34
+ $X2=7.725 $Y2=3.34
r189 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.64 $Y=3.255
+ $X2=7.725 $Y2=3.34
r190 36 37 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=7.64 $Y=2.025
+ $X2=7.64 $Y2=3.255
r191 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.555 $Y=1.94
+ $X2=7.64 $Y2=2.025
r192 34 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.555 $Y=1.94
+ $X2=7.025 $Y2=1.94
r193 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.94 $Y=2.025
+ $X2=7.025 $Y2=1.94
r194 32 33 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=6.94 $Y=2.025
+ $X2=6.94 $Y2=3.635
r195 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.855 $Y=3.72
+ $X2=6.94 $Y2=3.635
r196 30 31 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.855 $Y=3.72
+ $X2=6.325 $Y2=3.72
r197 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.24 $Y=3.635
+ $X2=6.325 $Y2=3.72
r198 28 29 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.24 $Y=3.185
+ $X2=6.24 $Y2=3.635
r199 27 52 3.71787 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=5.055 $Y=3.1 $X2=4.855
+ $Y2=3.1
r200 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.155 $Y=3.1
+ $X2=6.24 $Y2=3.185
r201 26 27 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=6.155 $Y=3.1
+ $X2=5.055 $Y2=3.1
r202 25 52 2.43149 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.97 $Y=3.015
+ $X2=4.855 $Y2=3.1
r203 24 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.97 $Y=1.095
+ $X2=4.97 $Y2=3.015
r204 20 52 2.43149 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=4.78 $Y=3.185
+ $X2=4.855 $Y2=3.1
r205 20 22 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=4.78 $Y=3.185
+ $X2=4.78 $Y2=3.485
r206 19 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=1.01
+ $X2=3.44 $Y2=1.01
r207 18 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.885 $Y=1.01
+ $X2=4.97 $Y2=1.095
r208 18 19 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=4.885 $Y=1.01
+ $X2=3.605 $Y2=1.01
r209 17 46 13.1569 $w=3.57e-07 $l=4.82623e-07 $layer=LI1_cond $X=2.115 $Y=3.1
+ $X2=1.895 $Y2=3.485
r210 16 52 3.71787 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=4.655 $Y=3.1 $X2=4.855
+ $Y2=3.1
r211 16 17 165.711 $w=1.68e-07 $l=2.54e-06 $layer=LI1_cond $X=4.655 $Y=3.1
+ $X2=2.115 $Y2=3.1
r212 5 56 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=8.295
+ $Y=3.295 $X2=8.44 $Y2=3.505
r213 4 22 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.68
+ $Y=3.275 $X2=4.82 $Y2=3.485
r214 3 46 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=1.695
+ $Y=3.275 $X2=1.84 $Y2=3.485
r215 2 59 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=8.43
+ $Y=0.63 $X2=8.575 $Y2=0.85
r216 1 48 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=3.3
+ $Y=0.535 $X2=3.44 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%Q_N 1 2 7 8 9 10 11 12 13 22
r19 13 41 7.49088 $w=3.98e-07 $l=2.6e-07 $layer=LI1_cond $X=17.635 $Y=3.145
+ $X2=17.635 $Y2=3.405
r20 12 13 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=17.635 $Y=2.775
+ $X2=17.635 $Y2=3.145
r21 11 12 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=17.635 $Y=2.405
+ $X2=17.635 $Y2=2.775
r22 11 33 6.05033 $w=3.98e-07 $l=2.1e-07 $layer=LI1_cond $X=17.635 $Y=2.405
+ $X2=17.635 $Y2=2.195
r23 10 33 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=17.635 $Y=2.035
+ $X2=17.635 $Y2=2.195
r24 9 10 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=17.635 $Y=1.665
+ $X2=17.635 $Y2=2.035
r25 8 9 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=17.635 $Y=1.295
+ $X2=17.635 $Y2=1.665
r26 7 8 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=17.635 $Y=0.925
+ $X2=17.635 $Y2=1.295
r27 7 22 7.05871 $w=3.98e-07 $l=2.45e-07 $layer=LI1_cond $X=17.635 $Y=0.925
+ $X2=17.635 $Y2=0.68
r28 2 41 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=17.5
+ $Y=2.05 $X2=17.64 $Y2=3.405
r29 2 33 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=17.5
+ $Y=2.05 $X2=17.64 $Y2=2.195
r30 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=17.53
+ $Y=0.535 $X2=17.67 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%Q 1 2 7 8 9 10 11 12 13
r12 13 39 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=19.87 $Y=3.145
+ $X2=19.87 $Y2=3.59
r13 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=19.87 $Y=2.775
+ $X2=19.87 $Y2=3.145
r14 11 12 14.7445 $w=3.38e-07 $l=4.35e-07 $layer=LI1_cond $X=19.87 $Y=2.34
+ $X2=19.87 $Y2=2.775
r15 10 11 10.3381 $w=3.38e-07 $l=3.05e-07 $layer=LI1_cond $X=19.87 $Y=2.035
+ $X2=19.87 $Y2=2.34
r16 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=19.87 $Y=1.665
+ $X2=19.87 $Y2=2.035
r17 8 9 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=19.87 $Y=1.295
+ $X2=19.87 $Y2=1.665
r18 7 8 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=19.87 $Y=0.85
+ $X2=19.87 $Y2=1.295
r19 2 39 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=19.725
+ $Y=2.215 $X2=19.865 $Y2=3.59
r20 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=19.725
+ $Y=2.215 $X2=19.865 $Y2=2.34
r21 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=19.735
+ $Y=0.705 $X2=19.875 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%VGND 1 2 3 4 5 6 7 22 25 32 41 55 58 67 74
+ 78
r137 80 82 5.90737 $w=9.48e-07 $l=4.6e-07 $layer=LI1_cond $X=19.04 $Y=0.85
+ $X2=19.04 $Y2=1.31
r138 75 78 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=18.68 $Y=0.44
+ $X2=19.4 $Y2=0.44
r139 74 80 4.75158 $w=9.48e-07 $l=3.7e-07 $layer=LI1_cond $X=19.04 $Y=0.48
+ $X2=19.04 $Y2=0.85
r140 74 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=19.4 $Y=0.48
+ $X2=19.4 $Y2=0.48
r141 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=18.68 $Y=0.48
+ $X2=18.68 $Y2=0.48
r142 68 75 0.579697 $w=3.7e-07 $l=1.51e-06 $layer=MET1_cond $X=17.17 $Y=0.44
+ $X2=18.68 $Y2=0.44
r143 67 71 4.5135 $w=5.28e-07 $l=2e-07 $layer=LI1_cond $X=16.99 $Y=0.48
+ $X2=16.99 $Y2=0.68
r144 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.17 $Y=0.48
+ $X2=17.17 $Y2=0.48
r145 62 68 0.723662 $w=3.7e-07 $l=1.885e-06 $layer=MET1_cond $X=15.285 $Y=0.44
+ $X2=17.17 $Y2=0.44
r146 59 62 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=14.565 $Y=0.44
+ $X2=15.285 $Y2=0.44
r147 58 64 3.27474 $w=9.48e-07 $l=2.55e-07 $layer=LI1_cond $X=14.925 $Y=0.48
+ $X2=14.925 $Y2=0.735
r148 58 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.285 $Y=0.48
+ $X2=15.285 $Y2=0.48
r149 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.565 $Y=0.48
+ $X2=14.565 $Y2=0.48
r150 53 59 1.13636 $w=3.7e-07 $l=2.96e-06 $layer=MET1_cond $X=11.605 $Y=0.44
+ $X2=14.565 $Y2=0.44
r151 52 55 1.06146 $w=3.78e-07 $l=3.5e-08 $layer=LI1_cond $X=11.605 $Y=0.555
+ $X2=11.64 $Y2=0.555
r152 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.605 $Y=0.48
+ $X2=11.605 $Y2=0.48
r153 49 53 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.885 $Y=0.44
+ $X2=11.605 $Y2=0.44
r154 48 52 21.8358 $w=3.78e-07 $l=7.2e-07 $layer=LI1_cond $X=10.885 $Y=0.555
+ $X2=11.605 $Y2=0.555
r155 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.885 $Y=0.48
+ $X2=10.885 $Y2=0.48
r156 41 45 5.27528 $w=8.48e-07 $l=3.5e-07 $layer=LI1_cond $X=7.295 $Y=0.48
+ $X2=7.295 $Y2=0.83
r157 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.555 $Y=0.48
+ $X2=7.555 $Y2=0.48
r158 36 42 0.554743 $w=3.7e-07 $l=1.445e-06 $layer=MET1_cond $X=6.11 $Y=0.44
+ $X2=7.555 $Y2=0.44
r159 33 36 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.39 $Y=0.44
+ $X2=6.11 $Y2=0.44
r160 32 38 4.49474 $w=9.48e-07 $l=3.5e-07 $layer=LI1_cond $X=5.75 $Y=0.48
+ $X2=5.75 $Y2=0.83
r161 32 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.11 $Y=0.48
+ $X2=6.11 $Y2=0.48
r162 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.39 $Y=0.48
+ $X2=5.39 $Y2=0.48
r163 26 33 1.86194 $w=3.7e-07 $l=4.85e-06 $layer=MET1_cond $X=0.54 $Y=0.44
+ $X2=5.39 $Y2=0.44
r164 25 29 8.44936 $w=5.43e-07 $l=3.85e-07 $layer=LI1_cond $X=0.362 $Y=0.48
+ $X2=0.362 $Y2=0.865
r165 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.54 $Y=0.48
+ $X2=0.54 $Y2=0.48
r166 22 49 0.309044 $w=3.7e-07 $l=8.05e-07 $layer=MET1_cond $X=10.08 $Y=0.44
+ $X2=10.885 $Y2=0.44
r167 22 42 0.969361 $w=3.7e-07 $l=2.525e-06 $layer=MET1_cond $X=10.08 $Y=0.44
+ $X2=7.555 $Y2=0.44
r168 7 82 182 $w=1.7e-07 $l=7.12881e-07 $layer=licon1_NDIFF $count=1 $X=18.86
+ $Y=0.705 $X2=19.095 $Y2=1.31
r169 7 80 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=18.86
+ $Y=0.705 $X2=19.095 $Y2=0.85
r170 6 71 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=16.765
+ $Y=0.535 $X2=16.89 $Y2=0.68
r171 5 64 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=14.705
+ $Y=0.535 $X2=14.845 $Y2=0.735
r172 4 55 182 $w=1.7e-07 $l=2.39531e-07 $layer=licon1_NDIFF $count=1 $X=11.415
+ $Y=0.63 $X2=11.64 $Y2=0.66
r173 3 45 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=7.06
+ $Y=0.63 $X2=7.205 $Y2=0.83
r174 2 38 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=5.67
+ $Y=0.63 $X2=5.81 $Y2=0.83
r175 1 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.325
+ $Y=0.655 $X2=0.47 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRBP_1%noxref_25 1 2 9 11 12 13
r31 13 16 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=4.93 $Y=0.35
+ $X2=4.93 $Y2=0.67
r32 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=0.35
+ $X2=4.93 $Y2=0.35
r33 11 12 172.888 $w=1.68e-07 $l=2.65e-06 $layer=LI1_cond $X=4.765 $Y=0.35
+ $X2=2.115 $Y2=0.35
r34 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.99 $Y=0.435
+ $X2=2.115 $Y2=0.35
r35 7 9 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=1.99 $Y=0.435 $X2=1.99
+ $Y2=0.745
r36 2 16 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=4.79
+ $Y=0.535 $X2=4.93 $Y2=0.67
r37 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.535 $X2=1.95 $Y2=0.745
.ends

