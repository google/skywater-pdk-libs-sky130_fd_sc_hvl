* File: sky130_fd_sc_hvl__dfrtp_1.spice
* Created: Wed Sep  2 09:05:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__dfrtp_1.pex.spice"
.subckt sky130_fd_sc_hvl__dfrtp_1  VNB VPB CLK RESET_B D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* RESET_B	RESET_B
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_CLK_M1016_g N_A_30_107#_M1016_s N_VNB_M1016_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1028 N_A_339_537#_M1028_d N_A_30_107#_M1028_g N_VGND_M1016_d N_VNB_M1016_b NHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1012 A_637_173# N_RESET_B_M1012_g N_VGND_M1012_s N_VNB_M1016_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250000 SB=250007 A=0.21 P=1.84 MULT=1
MM1014 N_A_452_632#_M1014_d N_D_M1014_g A_637_173# N_VNB_M1016_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250001 SB=250006 A=0.21 P=1.84 MULT=1
MM1008 N_A_921_632#_M1008_d N_A_30_107#_M1008_g N_A_452_632#_M1014_d
+ N_VNB_M1016_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0
+ M=1 R=0.84 SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1020 A_1091_173# N_A_339_537#_M1020_g N_A_921_632#_M1008_d N_VNB_M1016_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1003 A_1233_173# N_A_1119_506#_M1003_g A_1091_173# N_VNB_M1016_b NHV L=0.5
+ W=0.42 AD=0.04935 AS=0.0441 PD=0.655 PS=0.63 NRD=16.9632 NRS=13.566 M=1 R=0.84
+ SA=250003 SB=250004 A=0.21 P=1.84 MULT=1
MM1029 N_VGND_M1029_d N_RESET_B_M1029_g A_1233_173# N_VNB_M1016_b NHV L=0.5
+ W=0.42 AD=0.233962 AS=0.04935 PD=1.44667 PS=0.655 NRD=136.264 NRS=16.9632 M=1
+ R=0.84 SA=250004 SB=250003 A=0.21 P=1.84 MULT=1
MM1004 N_A_1119_506#_M1004_d N_A_921_632#_M1004_g N_VGND_M1029_d N_VNB_M1016_b
+ NHV L=0.5 W=0.75 AD=0.105 AS=0.417788 PD=1.03 PS=2.58333 NRD=0 NRS=12.1524 M=1
+ R=1.5 SA=250003 SB=250003 A=0.375 P=2.5 MULT=1
MM1017 N_A_1875_543#_M1017_d N_A_339_537#_M1017_g N_A_1119_506#_M1004_d
+ N_VNB_M1016_b NHV L=0.5 W=0.75 AD=0.197019 AS=0.105 PD=1.60256 PS=1.03
+ NRD=1.5162 NRS=0 M=1 R=1.5 SA=250004 SB=250002 A=0.375 P=2.5 MULT=1
MM1030 A_2089_107# N_A_30_107#_M1030_g N_A_1875_543#_M1017_d N_VNB_M1016_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.110331 PD=0.63 PS=0.897436 NRD=13.566 NRS=56.9886
+ M=1 R=0.84 SA=250003 SB=250002 A=0.21 P=1.84 MULT=1
MM1031 N_VGND_M1031_d N_A_2096_417#_M1031_g A_2089_107# N_VNB_M1016_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250004 SB=250002 A=0.21 P=1.84 MULT=1
MM1011 A_2387_107# N_RESET_B_M1011_g N_VGND_M1031_d N_VNB_M1016_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250005 SB=250001 A=0.21 P=1.84 MULT=1
MM1023 N_A_2096_417#_M1023_d N_A_1875_543#_M1023_g A_2387_107# N_VNB_M1016_b NHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250005 SB=250000 A=0.21 P=1.84 MULT=1
MM1015 N_VGND_M1015_d N_A_1875_543#_M1015_g N_A_2649_207#_M1015_s N_VNB_M1016_b
+ NHV L=0.5 W=0.42 AD=0.0933154 AS=0.1197 PD=0.822051 PS=1.41 NRD=31.2132 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1002 N_Q_M1002_d N_A_2649_207#_M1002_g N_VGND_M1015_d N_VNB_M1016_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.166635 PD=2.07 PS=1.46795 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1018 N_VPWR_M1018_d N_CLK_M1018_g N_A_30_107#_M1018_s N_VPB_M1018_b PHV L=0.5
+ W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1000 N_A_339_537#_M1000_d N_A_30_107#_M1000_g N_VPWR_M1018_d N_VPB_M1018_b PHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1024 N_VPWR_M1024_d N_RESET_B_M1024_g N_A_452_632#_M1024_s N_VPB_M1018_b PHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250004 A=0.21 P=1.84 MULT=1
MM1009 N_A_452_632#_M1009_d N_D_M1009_g N_VPWR_M1024_d N_VPB_M1018_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250001
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1001 N_A_921_632#_M1001_d N_A_339_537#_M1001_g N_A_452_632#_M1009_d
+ N_VPB_M1018_b PHV L=0.5 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0
+ M=1 R=0.84 SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1013 A_1077_632# N_A_30_107#_M1013_g N_A_921_632#_M1001_d N_VPB_M1018_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1026 N_VPWR_M1026_d N_A_1119_506#_M1026_g A_1077_632# N_VPB_M1018_b PHV L=0.5
+ W=0.42 AD=0.0756 AS=0.0441 PD=0.78 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250003 SB=250001 A=0.21 P=1.84 MULT=1
MM1006 N_A_921_632#_M1006_d N_RESET_B_M1006_g N_VPWR_M1026_d N_VPB_M1018_b PHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0756 PD=1.41 PS=0.78 NRD=0 NRS=36.3664 M=1 R=0.84
+ SA=250004 SB=250000 A=0.21 P=1.84 MULT=1
MM1022 N_A_1119_506#_M1022_d N_A_921_632#_M1022_g N_VPWR_M1022_s N_VPB_M1018_b
+ PHV L=0.5 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=2 SA=250000
+ SB=250002 A=0.5 P=3 MULT=1
MM1007 N_A_1875_543#_M1007_d N_A_30_107#_M1007_g N_A_1119_506#_M1022_d
+ N_VPB_M1018_b PHV L=0.5 W=1 AD=0.233239 AS=0.14 PD=1.96479 PS=1.28 NRD=0 NRS=0
+ M=1 R=2 SA=250001 SB=250001 A=0.5 P=3 MULT=1
MM1027 A_2054_543# N_A_339_537#_M1027_g N_A_1875_543#_M1007_d N_VPB_M1018_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0979606 PD=0.63 PS=0.825211 NRD=22.729 NRS=52.2958
+ M=1 R=0.84 SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1021 N_VPWR_M1021_d N_A_2096_417#_M1021_g A_2054_543# N_VPB_M1018_b PHV L=0.5
+ W=0.42 AD=0.08085 AS=0.0441 PD=0.805 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1005 N_A_2096_417#_M1005_d N_RESET_B_M1005_g N_VPWR_M1021_d N_VPB_M1018_b PHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.08085 PD=0.7 PS=0.805 NRD=0 NRS=47.75 M=1 R=0.84
+ SA=250003 SB=250001 A=0.21 P=1.84 MULT=1
MM1025 N_VPWR_M1025_d N_A_1875_543#_M1025_g N_A_2096_417#_M1005_d N_VPB_M1018_b
+ PHV L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250004 SB=250000 A=0.21 P=1.84 MULT=1
MM1019 N_VPWR_M1019_d N_A_1875_543#_M1019_g N_A_2649_207#_M1019_s N_VPB_M1018_b
+ PHV L=0.5 W=0.75 AD=0.16 AS=0.21375 PD=1.25 PS=2.07 NRD=24.1806 NRS=0 M=1
+ R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1010 N_Q_M1010_d N_A_2649_207#_M1010_g N_VPWR_M1019_d N_VPB_M1018_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.32 PD=3.53 PS=2.5 NRD=0 NRS=0 M=1 R=3 SA=250000 SB=250000
+ A=0.75 P=4 MULT=1
DX32_noxref N_VNB_M1016_b N_VPB_M1018_b NWDIODE A=41.652 P=37.24
*
.include "sky130_fd_sc_hvl__dfrtp_1.pxi.spice"
*
.ends
*
*
