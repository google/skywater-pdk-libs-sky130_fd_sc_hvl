* NGSPICE file created from sky130_fd_sc_hvl__dfrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
M1000 a_2412_107# RESET_B VGND VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.24515e+12p ps=1.148e+07u
M1001 a_2122_348# a_1900_107# a_2412_107# VNB nhv w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1002 a_1900_107# a_37_107# a_1176_466# VPB phv w=1e+06u l=500000u
+  ad=3.312e+11p pd=2.79e+06u as=2.8e+11p ps=2.56e+06u
M1003 a_350_107# a_37_107# VGND VNB nhv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1004 VPWR CLK a_37_107# VPB phv w=750000u l=500000u
+  ad=2.2032e+12p pd=1.785e+07u as=2.1375e+11p ps=2.07e+06u
M1005 a_2114_107# a_37_107# a_1900_107# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=3.219e+11p ps=2.64e+06u
M1006 a_978_608# a_37_107# a_509_608# VNB nhv w=420000u l=500000u
+  ad=1.869e+11p pd=1.73e+06u as=1.176e+11p ps=1.4e+06u
M1007 VGND a_2122_348# a_2114_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_509_608# D VPWR VPB phv w=420000u l=500000u
+  ad=2.373e+11p pd=2.81e+06u as=0p ps=0u
M1009 a_1176_466# a_978_608# VPWR VPB phv w=1e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Q a_2937_443# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=0p ps=0u
M1011 a_978_608# RESET_B VPWR VPB phv w=420000u l=500000u
+  ad=2.373e+11p pd=2.81e+06u as=0p ps=0u
M1012 VPWR a_1900_107# a_2122_348# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1013 a_728_173# RESET_B VGND VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1014 a_509_608# D a_728_173# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_2079_462# a_350_107# a_1900_107# VPB phv w=420000u l=500000u
+  ad=9.03e+10p pd=1.27e+06u as=0p ps=0u
M1016 a_1900_107# a_350_107# a_1176_466# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=2.1e+11p ps=2.06e+06u
M1017 Q_N a_1900_107# VGND VNB nhv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
M1018 VPWR RESET_B a_509_608# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1134_608# a_37_107# a_978_608# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1020 VGND CLK a_37_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1021 Q a_2937_443# VGND VNB nhv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
M1022 VPWR a_1176_466# a_1134_608# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q_N a_1900_107# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=0p ps=0u
M1024 VGND a_1900_107# a_2937_443# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1025 a_2122_348# RESET_B VPWR VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_350_107# a_37_107# VPWR VPB phv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
M1027 VPWR a_2122_348# a_2079_462# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1215_173# a_350_107# a_978_608# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1029 VGND RESET_B a_1357_173# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=9.66e+10p ps=1.3e+06u
M1030 a_978_608# a_350_107# a_509_608# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1357_173# a_1176_466# a_1215_173# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1176_466# a_978_608# VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_1900_107# a_2937_443# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=2.1375e+11p ps=2.07e+06u
.ends

