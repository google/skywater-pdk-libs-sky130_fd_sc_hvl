* File: sky130_fd_sc_hvl__sdfxtp_1.pex.spice
* Created: Fri Aug 28 09:40:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%VNB 5 7 11
c115 11 0 1.09283e-19 $X=0.24 $Y=0
c116 5 0 1.30116e-19 $X=-0.33 $Y=-0.265
r117 7 11 0.000478831 $w=1.488e-05 $l=5.7e-08 $layer=MET1_cond $X=7.44 $Y=0.057
+ $X2=7.44 $Y2=0
r118 5 11 0.6 $w=1.7e-07 $l=2.635e-06 $layer=mcon $count=15 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r119 5 11 0.6 $w=1.7e-07 $l=2.635e-06 $layer=mcon $count=15 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%VPB 4 6 14
r136 10 14 0.6 $w=1.7e-07 $l=2.635e-06 $layer=mcon $count=15 $X=14.64 $Y=4.07
+ $X2=14.64 $Y2=4.07
r137 9 14 939.465 $w=1.68e-07 $l=1.44e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=14.64 $Y2=4.07
r138 9 10 0.6 $w=1.7e-07 $l=2.635e-06 $layer=mcon $count=15 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r139 6 10 0.000478831 $w=1.488e-05 $l=5.7e-08 $layer=MET1_cond $X=7.44 $Y=4.013
+ $X2=7.44 $Y2=4.07
r140 4 14 11.7419 $w=1.7e-07 $l=1.46824e-05 $layer=licon1_NTAP_notbjt $count=15
+ $X=0 $Y=3.985 $X2=14.64 $Y2=4.07
r141 4 9 11.7419 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=15
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%SCE 3 6 7 9 10 12 16 20 23 24 25 30 35 39
+ 48
c73 30 0 2.82364e-20 $X=2.95 $Y=0.745
r74 35 38 53.5029 $w=5.25e-07 $l=5.25e-07 $layer=POLY_cond $X=0.692 $Y=1.565
+ $X2=0.692 $Y2=2.09
r75 35 37 19.0243 $w=5.25e-07 $l=1.85e-07 $layer=POLY_cond $X=0.692 $Y=1.565
+ $X2=0.692 $Y2=1.38
r76 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.77
+ $Y=1.565 $X2=0.77 $Y2=1.565
r77 25 48 8.99479 $w=5.78e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.735
+ $X2=1.795 $Y2=1.735
r78 25 39 3.60886 $w=5.78e-07 $l=1.75e-07 $layer=LI1_cond $X=1.68 $Y=1.735
+ $X2=1.505 $Y2=1.735
r79 24 39 6.28972 $w=5.78e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=1.735
+ $X2=1.505 $Y2=1.735
r80 24 36 8.86748 $w=5.78e-07 $l=4.3e-07 $layer=LI1_cond $X=1.2 $Y=1.735
+ $X2=0.77 $Y2=1.735
r81 23 36 1.0311 $w=5.78e-07 $l=5e-08 $layer=LI1_cond $X=0.72 $Y=1.735 $X2=0.77
+ $Y2=1.735
r82 21 30 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.95 $Y=1.25 $X2=2.95
+ $Y2=0.745
r83 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.885
+ $Y=1.25 $X2=2.885 $Y2=1.25
r84 18 20 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=2.885 $Y=1.855
+ $X2=2.885 $Y2=1.25
r85 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.72 $Y=1.94
+ $X2=2.885 $Y2=1.855
r86 16 48 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=2.72 $Y=1.94
+ $X2=1.795 $Y2=1.94
r87 10 12 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.465 $Y=2.855
+ $X2=1.465 $Y2=3.175
r88 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.685 $Y=2.855 $X2=0.685
+ $Y2=3.175
r89 6 10 105.139 $w=3.53e-07 $l=8.86228e-07 $layer=POLY_cond $X=0.695 $Y=2.605
+ $X2=1.465 $Y2=2.855
r90 6 7 1.36544 $w=3.53e-07 $l=1e-08 $layer=POLY_cond $X=0.695 $Y=2.605
+ $X2=0.685 $Y2=2.605
r91 6 38 27.2659 $w=5.2e-07 $l=2.65e-07 $layer=POLY_cond $X=0.695 $Y=2.355
+ $X2=0.695 $Y2=2.09
r92 3 37 67.9487 $w=5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.68 $Y=0.745 $X2=0.68
+ $Y2=1.38
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%D 3 6 9 11 12 13 14 15 16 24
c45 16 0 2.82364e-20 $X=2.64 $Y=2.405
c46 9 0 3.21713e-20 $X=2.175 $Y=3.175
r47 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.635
+ $Y=2.29 $X2=1.635 $Y2=2.29
r48 22 24 12.2886 $w=4.04e-07 $l=1.03e-07 $layer=POLY_cond $X=1.532 $Y=2.355
+ $X2=1.635 $Y2=2.355
r49 15 16 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=2.362
+ $X2=2.64 $Y2=2.362
r50 14 15 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.362
+ $X2=2.16 $Y2=2.362
r51 14 25 1.64635 $w=3.13e-07 $l=4.5e-08 $layer=LI1_cond $X=1.68 $Y=2.362
+ $X2=1.635 $Y2=2.362
r52 13 25 15.9147 $w=3.13e-07 $l=4.35e-07 $layer=LI1_cond $X=1.2 $Y=2.362
+ $X2=1.635 $Y2=2.362
r53 12 13 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=2.362 $X2=1.2
+ $Y2=2.362
r54 7 24 64.4257 $w=4.04e-07 $l=7.00999e-07 $layer=POLY_cond $X=2.175 $Y=2.725
+ $X2=1.635 $Y2=2.355
r55 7 9 48.1527 $w=5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.175 $Y=2.725 $X2=2.175
+ $Y2=3.175
r56 6 22 5.95965 $w=3.55e-07 $l=3.7e-07 $layer=POLY_cond $X=1.532 $Y=1.985
+ $X2=1.532 $Y2=2.355
r57 6 11 65.0188 $w=3.55e-07 $l=4e-07 $layer=POLY_cond $X=1.532 $Y=1.985
+ $X2=1.532 $Y2=1.585
r58 1 11 31.3249 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.46 $Y=1.335 $X2=1.46
+ $Y2=1.585
r59 1 3 63.1335 $w=5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.46 $Y=1.335 $X2=1.46
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%A_30_593# 1 2 7 9 12 16 20 22 26 28 31
r64 29 31 2.47603 $w=5.84e-07 $l=3e-08 $layer=POLY_cond $X=2.14 $Y=1.525
+ $X2=2.17 $Y2=1.525
r65 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.14
+ $Y=1.25 $X2=2.14 $Y2=1.25
r66 23 26 3.35233 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.455 $Y=1.18
+ $X2=0.29 $Y2=1.18
r67 22 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=1.18
+ $X2=2.14 $Y2=1.18
r68 22 23 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=1.975 $Y=1.18
+ $X2=0.455 $Y2=1.18
r69 18 26 3.22182 $w=2.92e-07 $l=1.0225e-07 $layer=LI1_cond $X=0.252 $Y=1.265
+ $X2=0.29 $Y2=1.18
r70 18 20 86.3202 $w=2.53e-07 $l=1.91e-06 $layer=LI1_cond $X=0.252 $Y=1.265
+ $X2=0.252 $Y2=3.175
r71 14 26 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=0.29 $Y=1.095
+ $X2=0.29 $Y2=1.18
r72 14 16 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.29 $Y=1.095
+ $X2=0.29 $Y2=0.745
r73 10 31 64.7894 $w=5.84e-07 $l=1.09413e-06 $layer=POLY_cond $X=2.955 $Y=2.265
+ $X2=2.17 $Y2=1.525
r74 10 12 97.3754 $w=5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.955 $Y=2.265
+ $X2=2.955 $Y2=3.175
r75 7 31 6.50804 $w=5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.17 $Y=1.065 $X2=2.17
+ $Y2=1.525
r76 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.17 $Y=1.065 $X2=2.17
+ $Y2=0.745
r77 2 20 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.965 $X2=0.295 $Y2=3.175
r78 1 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.535 $X2=0.29 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%SCD 3 7 12 13 16 18
r42 16 19 53.8061 $w=5.35e-07 $l=5.35e-07 $layer=POLY_cond $X=3.682 $Y=2.3
+ $X2=3.682 $Y2=2.835
r43 16 18 18.8041 $w=5.35e-07 $l=1.85e-07 $layer=POLY_cond $X=3.682 $Y=2.3
+ $X2=3.682 $Y2=2.115
r44 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.765
+ $Y=2.3 $X2=3.765 $Y2=2.3
r45 13 17 6.85027 $w=5.48e-07 $l=3.15e-07 $layer=LI1_cond $X=4.08 $Y=2.49
+ $X2=3.765 $Y2=2.49
r46 12 18 56.7131 $w=5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.7 $Y=1.585 $X2=3.7
+ $Y2=2.115
r47 11 12 49.5398 $w=5.4e-07 $l=5e-07 $layer=POLY_cond $X=3.68 $Y=1.085 $X2=3.68
+ $Y2=1.585
r48 7 19 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.665 $Y=3.175 $X2=3.665
+ $Y2=2.835
r49 3 11 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.66 $Y=0.745 $X2=3.66
+ $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%CLK 3 6 8 11 13
r35 11 14 48.459 $w=6e-07 $l=5.25e-07 $layer=POLY_cond $X=4.49 $Y=1.26 $X2=4.49
+ $Y2=1.785
r36 11 13 18.1407 $w=6e-07 $l=1.85e-07 $layer=POLY_cond $X=4.49 $Y=1.26 $X2=4.49
+ $Y2=1.075
r37 8 11 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.51 $Y=1.26
+ $X2=4.51 $Y2=1.26
r38 6 14 166.394 $w=5e-07 $l=1.555e-06 $layer=POLY_cond $X=4.54 $Y=3.34 $X2=4.54
+ $Y2=1.785
r39 3 13 31.812 $w=5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.44 $Y=0.745 $X2=4.44
+ $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%A_1204_107# 1 2 7 9 12 16 20 24 26 27 28
+ 29 33 34 39 41 42 45 49 51 53 55 61
c148 55 0 1.09283e-19 $X=7.98 $Y=0.745
c149 41 0 2.13081e-20 $X=10.045 $Y=1.34
c150 34 0 1.4382e-19 $X=7.935 $Y=0.35
c151 16 0 1.58977e-19 $X=11.26 $Y=2.925
r152 61 62 83.177 $w=4.52e-07 $l=7.8e-07 $layer=POLY_cond $X=10.48 $Y=1.71
+ $X2=11.26 $Y2=1.71
r153 49 52 7.26135 $w=3.63e-07 $l=1.25e-07 $layer=LI1_cond $X=7.142 $Y=2.39
+ $X2=7.142 $Y2=2.515
r154 49 51 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=7.142 $Y=2.39
+ $X2=7.142 $Y2=2.225
r155 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.125
+ $Y=2.39 $X2=7.125 $Y2=2.39
r156 46 61 28.792 $w=4.52e-07 $l=2.7e-07 $layer=POLY_cond $X=10.21 $Y=1.71
+ $X2=10.48 $Y2=1.71
r157 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.21
+ $Y=1.61 $X2=10.21 $Y2=1.61
r158 43 45 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=10.17 $Y=1.425
+ $X2=10.17 $Y2=1.61
r159 41 43 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.045 $Y=1.34
+ $X2=10.17 $Y2=1.425
r160 41 42 119.717 $w=1.68e-07 $l=1.835e-06 $layer=LI1_cond $X=10.045 $Y=1.34
+ $X2=8.21 $Y2=1.34
r161 40 55 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.98 $Y=1.25 $X2=7.98
+ $Y2=0.745
r162 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.045
+ $Y=1.25 $X2=8.045 $Y2=1.25
r163 37 42 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=8.072 $Y=1.255
+ $X2=8.21 $Y2=1.34
r164 37 39 0.209535 $w=2.73e-07 $l=5e-09 $layer=LI1_cond $X=8.072 $Y=1.255
+ $X2=8.072 $Y2=1.25
r165 36 39 34.1542 $w=2.73e-07 $l=8.15e-07 $layer=LI1_cond $X=8.072 $Y=0.435
+ $X2=8.072 $Y2=1.25
r166 35 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.245 $Y=0.35
+ $X2=7.16 $Y2=0.35
r167 34 36 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=7.935 $Y=0.35
+ $X2=8.072 $Y2=0.435
r168 34 35 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.935 $Y=0.35
+ $X2=7.245 $Y2=0.35
r169 33 52 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=7.24 $Y=3.335
+ $X2=7.24 $Y2=2.515
r170 30 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.16 $Y=0.435
+ $X2=7.16 $Y2=0.35
r171 30 51 116.781 $w=1.68e-07 $l=1.79e-06 $layer=LI1_cond $X=7.16 $Y=0.435
+ $X2=7.16 $Y2=2.225
r172 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.155 $Y=3.42
+ $X2=7.24 $Y2=3.335
r173 28 29 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.155 $Y=3.42
+ $X2=6.425 $Y2=3.42
r174 26 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.075 $Y=0.35
+ $X2=7.16 $Y2=0.35
r175 26 27 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=7.075 $Y=0.35
+ $X2=6.325 $Y2=0.35
r176 22 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.26 $Y=3.335
+ $X2=6.425 $Y2=3.42
r177 22 24 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=6.26 $Y=3.335
+ $X2=6.26 $Y2=3.11
r178 18 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.16 $Y=0.435
+ $X2=6.325 $Y2=0.35
r179 18 20 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.16 $Y=0.435
+ $X2=6.16 $Y2=0.745
r180 14 62 0.360583 $w=5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.26 $Y=1.995
+ $X2=11.26 $Y2=1.71
r181 14 16 99.5155 $w=5e-07 $l=9.3e-07 $layer=POLY_cond $X=11.26 $Y=1.995
+ $X2=11.26 $Y2=2.925
r182 10 61 0.360583 $w=5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.48 $Y=1.425
+ $X2=10.48 $Y2=1.71
r183 10 12 72.764 $w=5e-07 $l=6.8e-07 $layer=POLY_cond $X=10.48 $Y=1.425
+ $X2=10.48 $Y2=0.745
r184 7 50 18.6365 $w=6.31e-07 $l=2.47538e-07 $layer=POLY_cond $X=7.2 $Y=2.605
+ $X2=7.13 $Y2=2.39
r185 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.2 $Y=2.605 $X2=7.2
+ $Y2=2.925
r186 2 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.12
+ $Y=2.965 $X2=6.26 $Y2=3.11
r187 1 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.02
+ $Y=0.535 $X2=6.16 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%A_938_107# 1 2 7 9 11 15 19 23 26 27 28 29
+ 30 33 40 44 45 46 48 49 53 57 61 63 66 68 70 75 81 84 91
c192 91 0 5.71718e-20 $X=7.98 $Y=1.725
c193 84 0 1.16941e-19 $X=11.3 $Y=0.745
c194 68 0 3.33405e-19 $X=10.405 $Y=2.4
r195 90 91 63.3997 $w=5.93e-07 $l=7.8e-07 $layer=POLY_cond $X=7.2 $Y=1.725
+ $X2=7.98 $Y2=1.725
r196 73 88 28.7947 $w=7e-07 $l=3.99349e-07 $layer=POLY_cond $X=5.77 $Y=1.275
+ $X2=5.687 $Y2=1.635
r197 70 71 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.405 $Y=3.24
+ $X2=10.405 $Y2=3.41
r198 66 81 88.2799 $w=5e-07 $l=8.25e-07 $layer=POLY_cond $X=10.365 $Y=2.39
+ $X2=10.365 $Y2=3.215
r199 65 68 4.66986 $w=1.88e-07 $l=8e-08 $layer=LI1_cond $X=10.325 $Y=2.4
+ $X2=10.405 $Y2=2.4
r200 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.325
+ $Y=2.39 $X2=10.325 $Y2=2.39
r201 62 73 2.67515 $w=5e-07 $l=2.5e-08 $layer=POLY_cond $X=5.77 $Y=1.25 $X2=5.77
+ $Y2=1.275
r202 62 75 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.77 $Y=1.25 $X2=5.77
+ $Y2=0.745
r203 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.705
+ $Y=1.25 $X2=5.705 $Y2=1.25
r204 57 59 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=4.845 $Y=0.745
+ $X2=4.845 $Y2=0.975
r205 54 84 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=11.3 $Y=1.25 $X2=11.3
+ $Y2=0.745
r206 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.355
+ $Y=1.25 $X2=11.355 $Y2=1.25
r207 51 53 118.019 $w=1.93e-07 $l=2.075e-06 $layer=LI1_cond $X=11.352 $Y=3.325
+ $X2=11.352 $Y2=1.25
r208 50 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.49 $Y=3.41
+ $X2=10.405 $Y2=3.41
r209 49 51 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=11.255 $Y=3.41
+ $X2=11.352 $Y2=3.325
r210 49 50 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=11.255 $Y=3.41
+ $X2=10.49 $Y2=3.41
r211 48 70 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=10.405 $Y=3.155
+ $X2=10.405 $Y2=3.24
r212 47 68 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=10.405 $Y=2.495
+ $X2=10.405 $Y2=2.4
r213 47 48 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=10.405 $Y=2.495
+ $X2=10.405 $Y2=3.155
r214 45 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.32 $Y=3.24
+ $X2=10.405 $Y2=3.24
r215 45 46 137.658 $w=1.68e-07 $l=2.11e-06 $layer=LI1_cond $X=10.32 $Y=3.24
+ $X2=8.21 $Y2=3.24
r216 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.125 $Y=3.155
+ $X2=8.21 $Y2=3.24
r217 44 63 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=8.125 $Y=3.155
+ $X2=8.125 $Y2=2.495
r218 41 91 5.28331 $w=5.93e-07 $l=6.5e-08 $layer=POLY_cond $X=8.045 $Y=1.725
+ $X2=7.98 $Y2=1.725
r219 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.045
+ $Y=2.05 $X2=8.045 $Y2=2.05
r220 38 63 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.045 $Y=2.33
+ $X2=8.045 $Y2=2.495
r221 38 40 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=8.045 $Y=2.33
+ $X2=8.045 $Y2=2.05
r222 34 88 45.79 $w=7e-07 $l=6.65e-07 $layer=POLY_cond $X=5.687 $Y=2.3 $X2=5.687
+ $Y2=1.635
r223 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.44
+ $Y=2.3 $X2=5.44 $Y2=2.3
r224 31 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.44 $Y=2.595
+ $X2=5.44 $Y2=2.3
r225 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.275 $Y=2.68
+ $X2=5.44 $Y2=2.595
r226 29 30 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.275 $Y=2.68
+ $X2=5.095 $Y2=2.68
r227 27 61 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=1.24
+ $X2=5.705 $Y2=1.24
r228 27 28 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.54 $Y=1.24
+ $X2=5.025 $Y2=1.24
r229 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.94 $Y=1.155
+ $X2=5.025 $Y2=1.24
r230 26 59 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.94 $Y=1.155
+ $X2=4.94 $Y2=0.975
r231 21 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.93 $Y=2.765
+ $X2=5.095 $Y2=2.68
r232 21 23 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.93 $Y=2.765
+ $X2=4.93 $Y2=3.11
r233 17 91 6.8647 $w=5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.98 $Y=2.175 $X2=7.98
+ $Y2=1.725
r234 17 19 80.2544 $w=5e-07 $l=7.5e-07 $layer=POLY_cond $X=7.98 $Y=2.175
+ $X2=7.98 $Y2=2.925
r235 13 90 6.8647 $w=5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.2 $Y=1.275 $X2=7.2
+ $Y2=1.725
r236 13 15 56.7131 $w=5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.2 $Y=1.275 $X2=7.2
+ $Y2=0.745
r237 12 88 2.14911 $w=7.2e-07 $l=4.33e-07 $layer=POLY_cond $X=6.12 $Y=1.635
+ $X2=5.687 $Y2=1.635
r238 11 90 18.3784 $w=7.2e-07 $l=2.91548e-07 $layer=POLY_cond $X=6.95 $Y=1.635
+ $X2=7.2 $Y2=1.725
r239 11 12 59.2726 $w=7.2e-07 $l=8.3e-07 $layer=POLY_cond $X=6.95 $Y=1.635
+ $X2=6.12 $Y2=1.635
r240 7 34 40.8447 $w=7e-07 $l=6.19782e-07 $layer=POLY_cond $X=5.87 $Y=2.835
+ $X2=5.687 $Y2=2.3
r241 7 9 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.87 $Y=2.835 $X2=5.87
+ $Y2=3.34
r242 2 23 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.79
+ $Y=2.965 $X2=4.93 $Y2=3.11
r243 1 57 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.69
+ $Y=0.535 $X2=4.83 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%A_1688_81# 1 2 9 12 16 17 20 22 27 29 30
+ 32 34 35 36 38 39 42
c86 30 0 1.30116e-19 $X=10.14 $Y=0.99
c87 29 0 1.16941e-19 $X=10.475 $Y=0.99
c88 17 0 1.0179e-19 $X=8.705 $Y=1.565
c89 16 0 1.4382e-19 $X=8.705 $Y=1.065
c90 12 0 1.22988e-19 $X=8.69 $Y=2.925
r91 38 39 9.33524 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=9.975 $Y=2.865
+ $X2=9.975 $Y2=2.675
r92 35 43 54.2411 $w=5.3e-07 $l=5.35e-07 $layer=POLY_cond $X=8.705 $Y=2.05
+ $X2=8.705 $Y2=2.585
r93 35 42 18.909 $w=5.3e-07 $l=1.85e-07 $layer=POLY_cond $X=8.705 $Y=2.05
+ $X2=8.705 $Y2=1.865
r94 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.785
+ $Y=2.05 $X2=8.785 $Y2=2.05
r95 31 32 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=10.56 $Y=1.075
+ $X2=10.56 $Y2=1.955
r96 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.475 $Y=0.99
+ $X2=10.56 $Y2=1.075
r97 29 30 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.475 $Y=0.99
+ $X2=10.14 $Y2=0.99
r98 28 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.98 $Y=2.04
+ $X2=9.895 $Y2=2.04
r99 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.475 $Y=2.04
+ $X2=10.56 $Y2=1.955
r100 27 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=10.475 $Y=2.04
+ $X2=9.98 $Y2=2.04
r101 25 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.895 $Y=2.125
+ $X2=9.895 $Y2=2.04
r102 25 39 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=9.895 $Y=2.125
+ $X2=9.895 $Y2=2.675
r103 22 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.975 $Y=0.905
+ $X2=10.14 $Y2=0.99
r104 22 24 2.95758 $w=3.3e-07 $l=8e-08 $layer=LI1_cond $X=9.975 $Y=0.905
+ $X2=9.975 $Y2=0.825
r105 21 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.95 $Y=2.04
+ $X2=8.785 $Y2=2.04
r106 20 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.81 $Y=2.04
+ $X2=9.895 $Y2=2.04
r107 20 21 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=9.81 $Y=2.04
+ $X2=8.95 $Y2=2.04
r108 17 42 32.1018 $w=5e-07 $l=3e-07 $layer=POLY_cond $X=8.72 $Y=1.565 $X2=8.72
+ $Y2=1.865
r109 16 17 50.4745 $w=5.3e-07 $l=5e-07 $layer=POLY_cond $X=8.705 $Y=1.065
+ $X2=8.705 $Y2=1.565
r110 12 43 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=8.69 $Y=2.925 $X2=8.69
+ $Y2=2.585
r111 9 16 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.69 $Y=0.745 $X2=8.69
+ $Y2=1.065
r112 2 38 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=9.835
+ $Y=2.715 $X2=9.975 $Y2=2.865
r113 1 24 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=9.835
+ $Y=0.535 $X2=9.975 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%A_1490_107# 1 2 8 11 13 17 21 24 25 27 31
c75 27 0 1.74428e-19 $X=9.585 $Y=0.91
c76 21 0 1.0179e-19 $X=7.59 $Y=0.765
c77 13 0 7.79532e-21 $X=7.59 $Y=2.925
c78 11 0 1.15193e-19 $X=7.63 $Y=2.8
r79 21 23 8.73685 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=7.59 $Y=0.765
+ $X2=7.59 $Y2=0.995
r80 18 31 163.184 $w=5e-07 $l=1.525e-06 $layer=POLY_cond $X=9.585 $Y=1.69
+ $X2=9.585 $Y2=3.215
r81 18 27 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=9.585 $Y=1.69
+ $X2=9.585 $Y2=0.91
r82 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.52
+ $Y=1.69 $X2=9.52 $Y2=1.69
r83 15 24 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.755 $Y=1.69
+ $X2=7.63 $Y2=1.69
r84 15 17 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=7.755 $Y=1.69
+ $X2=9.52 $Y2=1.69
r85 11 25 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=7.63 $Y=2.8
+ $X2=7.63 $Y2=2.675
r86 11 13 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=7.63 $Y=2.8
+ $X2=7.63 $Y2=2.925
r87 9 24 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=7.59 $Y=1.775
+ $X2=7.63 $Y2=1.69
r88 9 25 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=7.59 $Y=1.775 $X2=7.59
+ $Y2=2.675
r89 8 24 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.63 $Y=1.605 $X2=7.63
+ $Y2=1.69
r90 8 23 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=7.63 $Y=1.605
+ $X2=7.63 $Y2=0.995
r91 2 13 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.45
+ $Y=2.715 $X2=7.59 $Y2=2.925
r92 1 21 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=7.45
+ $Y=0.535 $X2=7.59 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%A_2352_81# 1 2 9 13 17 21 23 24 27 31 33
+ 35 40 41
c93 23 0 1.49663e-19 $X=13.965 $Y=1.8
r94 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.53
+ $Y=1.85 $X2=13.53 $Y2=1.85
r95 42 44 7.22199 $w=4.73e-07 $l=2.8e-07 $layer=LI1_cond $X=13.39 $Y=1.57
+ $X2=13.39 $Y2=1.85
r96 41 50 50.2236 $w=5.7e-07 $l=5.25e-07 $layer=POLY_cond $X=12.045 $Y=1.65
+ $X2=12.045 $Y2=2.175
r97 41 49 18.3095 $w=5.7e-07 $l=1.85e-07 $layer=POLY_cond $X=12.045 $Y=1.65
+ $X2=12.045 $Y2=1.465
r98 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.145
+ $Y=1.65 $X2=12.145 $Y2=1.65
r99 35 37 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=13.275 $Y=2.86
+ $X2=13.275 $Y2=3.57
r100 33 44 5.38397 $w=4.73e-07 $l=2.14942e-07 $layer=LI1_cond $X=13.275 $Y=2.015
+ $X2=13.39 $Y2=1.85
r101 33 35 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=13.275 $Y=2.015
+ $X2=13.275 $Y2=2.86
r102 29 42 3.32055 $w=4.73e-07 $l=1.51658e-07 $layer=LI1_cond $X=13.275 $Y=1.485
+ $X2=13.39 $Y2=1.57
r103 29 31 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=13.275 $Y=1.485
+ $X2=13.275 $Y2=0.68
r104 28 40 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.31 $Y=1.57
+ $X2=12.145 $Y2=1.57
r105 27 42 6.80958 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=13.11 $Y=1.57
+ $X2=13.39 $Y2=1.57
r106 27 28 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=13.11 $Y=1.57
+ $X2=12.31 $Y2=1.57
r107 23 45 40.8312 $w=5.7e-07 $l=4.35e-07 $layer=POLY_cond $X=13.965 $Y=1.8
+ $X2=13.53 $Y2=1.8
r108 23 24 3.45798 $w=5.7e-07 $l=2.5e-07 $layer=POLY_cond $X=13.965 $Y=1.8
+ $X2=14.215 $Y2=1.8
r109 19 24 22.7291 $w=5e-07 $l=2.85e-07 $layer=POLY_cond $X=14.215 $Y=2.085
+ $X2=14.215 $Y2=1.8
r110 19 21 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=14.215 $Y=2.085
+ $X2=14.215 $Y2=2.965
r111 15 24 22.7291 $w=5e-07 $l=2.85e-07 $layer=POLY_cond $X=14.215 $Y=1.515
+ $X2=14.215 $Y2=1.8
r112 15 17 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=14.215 $Y=1.515
+ $X2=14.215 $Y2=1.01
r113 13 50 80.2544 $w=5e-07 $l=7.5e-07 $layer=POLY_cond $X=12.01 $Y=2.925
+ $X2=12.01 $Y2=2.175
r114 9 49 77.0442 $w=5e-07 $l=7.2e-07 $layer=POLY_cond $X=12.01 $Y=0.745
+ $X2=12.01 $Y2=1.465
r115 2 37 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=13.135
+ $Y=2.715 $X2=13.275 $Y2=3.57
r116 2 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.135
+ $Y=2.715 $X2=13.275 $Y2=2.86
r117 1 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.135
+ $Y=0.535 $X2=13.275 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%A_2123_543# 1 2 9 13 18 19 20 22 23 24 27
+ 28 33
c96 27 0 1.49663e-19 $X=12.765 $Y=2.01
r97 31 33 4.96245 $w=4.68e-07 $l=1.95e-07 $layer=LI1_cond $X=10.755 $Y=2.91
+ $X2=10.95 $Y2=2.91
r98 28 37 56.0721 $w=5.55e-07 $l=5.75e-07 $layer=POLY_cond $X=12.857 $Y=2.01
+ $X2=12.857 $Y2=2.585
r99 28 36 18.4754 $w=5.55e-07 $l=1.85e-07 $layer=POLY_cond $X=12.857 $Y=2.01
+ $X2=12.857 $Y2=1.825
r100 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.765
+ $Y=2.01 $X2=12.765 $Y2=2.01
r101 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=12.765 $Y=2.345
+ $X2=12.765 $Y2=2.01
r102 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.6 $Y=2.43
+ $X2=12.765 $Y2=2.345
r103 23 24 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=12.6 $Y=2.43 $X2=11.8
+ $Y2=2.43
r104 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.715 $Y=2.345
+ $X2=11.8 $Y2=2.43
r105 21 22 109.604 $w=1.68e-07 $l=1.68e-06 $layer=LI1_cond $X=11.715 $Y=0.665
+ $X2=11.715 $Y2=2.345
r106 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.63 $Y=0.58
+ $X2=11.715 $Y2=0.665
r107 19 20 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=11.63 $Y=0.58
+ $X2=11.075 $Y2=0.58
r108 16 33 4.43409 $w=2.5e-07 $l=2.35e-07 $layer=LI1_cond $X=10.95 $Y=2.675
+ $X2=10.95 $Y2=2.91
r109 16 18 88.9686 $w=2.48e-07 $l=1.93e-06 $layer=LI1_cond $X=10.95 $Y=2.675
+ $X2=10.95 $Y2=0.745
r110 15 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.95 $Y=0.665
+ $X2=11.075 $Y2=0.58
r111 15 18 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=10.95 $Y=0.665
+ $X2=10.95 $Y2=0.745
r112 13 37 67.4137 $w=5e-07 $l=6.3e-07 $layer=POLY_cond $X=12.885 $Y=3.215
+ $X2=12.885 $Y2=2.585
r113 9 36 97.9104 $w=5e-07 $l=9.15e-07 $layer=POLY_cond $X=12.885 $Y=0.91
+ $X2=12.885 $Y2=1.825
r114 2 31 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=10.615
+ $Y=2.715 $X2=10.755 $Y2=2.91
r115 1 18 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=10.73
+ $Y=0.535 $X2=10.91 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%VPWR 1 2 3 4 5 6 19 22 31 42 54 58 69 74
r93 72 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.675 $Y=3.59
+ $X2=14.675 $Y2=3.59
r94 69 72 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=14.495 $Y=2.36
+ $X2=14.495 $Y2=3.57
r95 66 74 0.714064 $w=3.7e-07 $l=1.86e-06 $layer=MET1_cond $X=12.815 $Y=3.63
+ $X2=14.675 $Y2=3.63
r96 64 66 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=12.095 $Y=3.63
+ $X2=12.815 $Y2=3.63
r97 63 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.815 $Y=3.59
+ $X2=12.815 $Y2=3.59
r98 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.095 $Y=3.59
+ $X2=12.095 $Y2=3.59
r99 61 63 4.81579 $w=9.48e-07 $l=3.75e-07 $layer=LI1_cond $X=12.455 $Y=3.215
+ $X2=12.455 $Y2=3.59
r100 58 61 4.55895 $w=9.48e-07 $l=3.55e-07 $layer=LI1_cond $X=12.455 $Y=2.86
+ $X2=12.455 $Y2=3.215
r101 55 64 0.856109 $w=3.7e-07 $l=2.23e-06 $layer=MET1_cond $X=9.865 $Y=3.63
+ $X2=12.095 $Y2=3.63
r102 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.865 $Y=3.62
+ $X2=9.865 $Y2=3.62
r103 50 55 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=9.145 $Y=3.63
+ $X2=9.865 $Y2=3.63
r104 49 54 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=9.145 $Y=3.63
+ $X2=9.865 $Y2=3.63
r105 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.145 $Y=3.62
+ $X2=9.145 $Y2=3.62
r106 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.79 $Y=3.59
+ $X2=5.79 $Y2=3.59
r107 42 45 9.73081 $w=5.88e-07 $l=4.8e-07 $layer=LI1_cond $X=5.61 $Y=3.11
+ $X2=5.61 $Y2=3.59
r108 39 46 0.506755 $w=3.7e-07 $l=1.32e-06 $layer=MET1_cond $X=4.47 $Y=3.63
+ $X2=5.79 $Y2=3.63
r109 37 39 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.75 $Y=3.63
+ $X2=4.47 $Y2=3.63
r110 36 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.47 $Y=3.59
+ $X2=4.47 $Y2=3.59
r111 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.75 $Y=3.59
+ $X2=3.75 $Y2=3.59
r112 34 36 0.256842 $w=9.48e-07 $l=2e-08 $layer=LI1_cond $X=4.11 $Y=3.57
+ $X2=4.11 $Y2=3.59
r113 31 34 5.90737 $w=9.48e-07 $l=4.6e-07 $layer=LI1_cond $X=4.11 $Y=3.11
+ $X2=4.11 $Y2=3.57
r114 28 37 0.76973 $w=3.7e-07 $l=2.005e-06 $layer=MET1_cond $X=1.745 $Y=3.63
+ $X2=3.75 $Y2=3.63
r115 26 28 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.025 $Y=3.63
+ $X2=1.745 $Y2=3.63
r116 25 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.745 $Y=3.59
+ $X2=1.745 $Y2=3.59
r117 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.025 $Y=3.59
+ $X2=1.025 $Y2=3.59
r118 22 25 5.32947 $w=9.48e-07 $l=4.15e-07 $layer=LI1_cond $X=1.385 $Y=3.175
+ $X2=1.385 $Y2=3.59
r119 19 50 0.654559 $w=3.7e-07 $l=1.705e-06 $layer=MET1_cond $X=7.44 $Y=3.63
+ $X2=9.145 $Y2=3.63
r120 19 46 0.633444 $w=3.7e-07 $l=1.65e-06 $layer=MET1_cond $X=7.44 $Y=3.63
+ $X2=5.79 $Y2=3.63
r121 6 72 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=14.465
+ $Y=2.215 $X2=14.605 $Y2=3.57
r122 6 69 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=14.465
+ $Y=2.215 $X2=14.605 $Y2=2.36
r123 5 61 300 $w=1.7e-07 $l=6.06218e-07 $layer=licon1_PDIFF $count=2 $X=12.26
+ $Y=2.715 $X2=12.495 $Y2=3.215
r124 5 58 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=12.26
+ $Y=2.715 $X2=12.495 $Y2=2.86
r125 4 49 600 $w=1.7e-07 $l=9.94359e-07 $layer=licon1_PDIFF $count=1 $X=8.94
+ $Y=2.715 $X2=9.195 $Y2=3.59
r126 3 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=5.355
+ $Y=2.965 $X2=5.48 $Y2=3.11
r127 2 34 600 $w=1.7e-07 $l=7.12881e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=2.965 $X2=4.15 $Y2=3.57
r128 2 31 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=2.965 $X2=4.15 $Y2=3.11
r129 1 22 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=2.965 $X2=1.075 $Y2=3.175
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%A_484_107# 1 2 3 4 13 15 18 20 21 24 28 32
+ 37 39 42 44 45
c96 44 0 3.58637e-20 $X=6.81 $Y=2.925
c97 15 0 3.21713e-20 $X=3.23 $Y=3.01
r98 44 45 10.5766 $w=3.63e-07 $l=2.3e-07 $layer=LI1_cond $X=6.792 $Y=2.925
+ $X2=6.792 $Y2=2.695
r99 39 41 9.43019 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=6.73 $Y=0.765
+ $X2=6.73 $Y2=0.995
r100 32 35 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=3.01
+ $X2=2.565 $Y2=3.175
r101 28 30 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.745
+ $X2=2.56 $Y2=0.83
r102 25 42 4.65272 $w=1.92e-07 $l=9.58123e-08 $layer=LI1_cond $X=6.695 $Y=2.035
+ $X2=6.672 $Y2=1.95
r103 25 45 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=6.695 $Y=2.035
+ $X2=6.695 $Y2=2.695
r104 24 42 4.65272 $w=1.92e-07 $l=8.5e-08 $layer=LI1_cond $X=6.672 $Y=1.865
+ $X2=6.672 $Y2=1.95
r105 24 41 46.6337 $w=2.13e-07 $l=8.7e-07 $layer=LI1_cond $X=6.672 $Y=1.865
+ $X2=6.672 $Y2=0.995
r106 22 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.4 $Y=1.95
+ $X2=3.315 $Y2=1.95
r107 21 42 1.79375 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=6.565 $Y=1.95
+ $X2=6.672 $Y2=1.95
r108 21 22 206.487 $w=1.68e-07 $l=3.165e-06 $layer=LI1_cond $X=6.565 $Y=1.95
+ $X2=3.4 $Y2=1.95
r109 19 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=2.035
+ $X2=3.315 $Y2=1.95
r110 19 20 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.315 $Y=2.035
+ $X2=3.315 $Y2=2.925
r111 18 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=1.865
+ $X2=3.315 $Y2=1.95
r112 17 18 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.315 $Y=0.915
+ $X2=3.315 $Y2=1.865
r113 16 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=3.01
+ $X2=2.565 $Y2=3.01
r114 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.23 $Y=3.01
+ $X2=3.315 $Y2=2.925
r115 15 16 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.23 $Y=3.01 $X2=2.73
+ $Y2=3.01
r116 14 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0.83
+ $X2=2.56 $Y2=0.83
r117 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.23 $Y=0.83
+ $X2=3.315 $Y2=0.915
r118 13 14 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.23 $Y=0.83
+ $X2=2.725 $Y2=0.83
r119 4 44 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=6.685
+ $Y=2.715 $X2=6.81 $Y2=2.925
r120 3 35 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=2.965 $X2=2.565 $Y2=3.175
r121 2 39 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=6.585
+ $Y=0.535 $X2=6.73 $Y2=0.765
r122 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.42
+ $Y=0.535 $X2=2.56 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%Q 1 2 9 13 18 20 21 22 23
r38 22 23 20.1154 $w=2.73e-07 $l=4.8e-07 $layer=LI1_cond $X=14.16 $Y=1.642
+ $X2=14.64 $Y2=1.642
r39 20 21 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=13.84 $Y=2.36
+ $X2=13.84 $Y2=2.195
r40 17 22 5.86698 $w=2.73e-07 $l=1.4e-07 $layer=LI1_cond $X=14.02 $Y=1.642
+ $X2=14.16 $Y2=1.642
r41 17 18 1.20952 $w=2.75e-07 $l=4.9368e-07 $layer=LI1_cond $X=14.02 $Y=1.642
+ $X2=13.66 $Y2=1.325
r42 15 18 5.32718 $w=2.65e-07 $l=5.76325e-07 $layer=LI1_cond $X=13.935 $Y=1.78
+ $X2=13.66 $Y2=1.325
r43 15 21 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=13.935 $Y=1.78
+ $X2=13.935 $Y2=2.195
r44 11 20 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=13.84 $Y=2.375
+ $X2=13.84 $Y2=2.36
r45 11 13 38.2547 $w=3.58e-07 $l=1.195e-06 $layer=LI1_cond $X=13.84 $Y=2.375
+ $X2=13.84 $Y2=3.57
r46 7 18 5.32718 $w=2.65e-07 $l=1.8e-07 $layer=LI1_cond $X=13.84 $Y=1.325
+ $X2=13.66 $Y2=1.325
r47 7 9 17.4467 $w=3.58e-07 $l=5.45e-07 $layer=LI1_cond $X=13.84 $Y=1.325
+ $X2=13.84 $Y2=0.78
r48 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=13.7
+ $Y=2.215 $X2=13.825 $Y2=2.36
r49 2 13 300 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_PDIFF $count=2 $X=13.7
+ $Y=2.215 $X2=13.825 $Y2=3.57
r50 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=13.7
+ $Y=0.635 $X2=13.825 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXTP_1%VGND 1 2 3 4 5 6 19 28 32 41 48 57 68 69
r106 68 72 6.08175 $w=5.88e-07 $l=3e-07 $layer=LI1_cond $X=14.495 $Y=0.48
+ $X2=14.495 $Y2=0.78
r107 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.675 $Y=0.48
+ $X2=14.675 $Y2=0.48
r108 63 65 5.90737 $w=9.48e-07 $l=4.6e-07 $layer=LI1_cond $X=12.455 $Y=0.68
+ $X2=12.455 $Y2=1.14
r109 61 69 0.714064 $w=3.7e-07 $l=1.86e-06 $layer=MET1_cond $X=12.815 $Y=0.44
+ $X2=14.675 $Y2=0.44
r110 58 61 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=12.095 $Y=0.44
+ $X2=12.815 $Y2=0.44
r111 57 63 2.56842 $w=9.48e-07 $l=2e-07 $layer=LI1_cond $X=12.455 $Y=0.48
+ $X2=12.455 $Y2=0.68
r112 57 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.815 $Y=0.48
+ $X2=12.815 $Y2=0.48
r113 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.095 $Y=0.48
+ $X2=12.095 $Y2=0.48
r114 52 58 0.990476 $w=3.7e-07 $l=2.58e-06 $layer=MET1_cond $X=9.515 $Y=0.44
+ $X2=12.095 $Y2=0.44
r115 49 52 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.795 $Y=0.44
+ $X2=9.515 $Y2=0.44
r116 48 54 4.43053 $w=9.48e-07 $l=3.45e-07 $layer=LI1_cond $X=9.155 $Y=0.48
+ $X2=9.155 $Y2=0.825
r117 48 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.515 $Y=0.48
+ $X2=9.515 $Y2=0.48
r118 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.795 $Y=0.48
+ $X2=8.795 $Y2=0.48
r119 41 45 5.37222 $w=5.88e-07 $l=2.65e-07 $layer=LI1_cond $X=5.51 $Y=0.48
+ $X2=5.51 $Y2=0.745
r120 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.69 $Y=0.48
+ $X2=5.69 $Y2=0.48
r121 36 42 0.497158 $w=3.7e-07 $l=1.295e-06 $layer=MET1_cond $X=4.395 $Y=0.44
+ $X2=5.69 $Y2=0.44
r122 33 36 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.675 $Y=0.44
+ $X2=4.395 $Y2=0.44
r123 32 38 3.57238 $w=9.03e-07 $l=2.65e-07 $layer=LI1_cond $X=4.032 $Y=0.48
+ $X2=4.032 $Y2=0.745
r124 32 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.395 $Y=0.48
+ $X2=4.395 $Y2=0.48
r125 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.675 $Y=0.48
+ $X2=3.675 $Y2=0.48
r126 29 33 0.742857 $w=3.7e-07 $l=1.935e-06 $layer=MET1_cond $X=1.74 $Y=0.44
+ $X2=3.675 $Y2=0.44
r127 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.74 $Y=0.48
+ $X2=1.74 $Y2=0.48
r128 26 28 14.5704 $w=5.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.07 $Y=0.64
+ $X2=1.74 $Y2=0.64
r129 23 29 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.02 $Y=0.44
+ $X2=1.74 $Y2=0.44
r130 22 26 1.08734 $w=5.48e-07 $l=5e-08 $layer=LI1_cond $X=1.02 $Y=0.64 $X2=1.07
+ $Y2=0.64
r131 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.02 $Y=0.48
+ $X2=1.02 $Y2=0.48
r132 19 49 0.520192 $w=3.7e-07 $l=1.355e-06 $layer=MET1_cond $X=7.44 $Y=0.44
+ $X2=8.795 $Y2=0.44
r133 19 42 0.671834 $w=3.7e-07 $l=1.75e-06 $layer=MET1_cond $X=7.44 $Y=0.44
+ $X2=5.69 $Y2=0.44
r134 6 72 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.465
+ $Y=0.635 $X2=14.605 $Y2=0.78
r135 5 65 182 $w=1.7e-07 $l=7.12881e-07 $layer=licon1_NDIFF $count=1 $X=12.26
+ $Y=0.535 $X2=12.495 $Y2=1.14
r136 5 63 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=12.26
+ $Y=0.535 $X2=12.495 $Y2=0.68
r137 4 54 182 $w=1.7e-07 $l=3.97555e-07 $layer=licon1_NDIFF $count=1 $X=8.94
+ $Y=0.535 $X2=9.195 $Y2=0.825
r138 3 45 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.255
+ $Y=0.535 $X2=5.38 $Y2=0.745
r139 2 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.91
+ $Y=0.535 $X2=4.05 $Y2=0.745
r140 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.535 $X2=1.07 $Y2=0.745
.ends

