* File: sky130_fd_sc_hvl__buf_2.pex.spice
* Created: Fri Aug 28 09:33:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__BUF_2%VNB 5 7 11 25
r21 7 25 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0.058
r22 7 11 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0
r23 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r24 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_2%VPB 4 6 14 21
r23 10 21 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=4.07
+ $X2=1.68 $Y2=4.013
r24 10 14 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=4.07
+ $X2=3.12 $Y2=4.07
r25 9 14 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=3.12 $Y2=4.07
r26 9 10 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r27 6 21 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=4.012
+ $X2=1.68 $Y2=4.013
r28 4 14 52 $w=1.7e-07 $l=3.16221e-06 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=3.12 $Y2=4.07
r29 4 9 52 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_2%A_129_279# 1 2 7 9 10 12 15 17 19 20 24 28 30
+ 36 40
r56 37 38 1.65068 $w=5.84e-07 $l=2e-08 $layer=POLY_cond $X=0.895 $Y=1.75
+ $X2=0.915 $Y2=1.75
r57 34 40 1.65068 $w=5.84e-07 $l=2e-08 $layer=POLY_cond $X=1.715 $Y=1.75
+ $X2=1.695 $Y2=1.75
r58 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.715
+ $Y=1.59 $X2=1.715 $Y2=1.59
r59 30 33 3.12527 $w=2.93e-07 $l=8e-08 $layer=LI1_cond $X=1.717 $Y=1.51
+ $X2=1.717 $Y2=1.59
r60 26 36 3.58051 $w=2.6e-07 $l=8.9861e-08 $layer=LI1_cond $X=3.125 $Y=1.425
+ $X2=3.115 $Y2=1.51
r61 26 28 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=3.125 $Y=1.425
+ $X2=3.125 $Y2=1.075
r62 22 36 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=1.595
+ $X2=3.115 $Y2=1.51
r63 22 24 31.7989 $w=2.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.115 $Y=1.595
+ $X2=3.115 $Y2=2.34
r64 21 30 3.96227 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.865 $Y=1.51
+ $X2=1.717 $Y2=1.51
r65 20 36 2.90867 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.98 $Y=1.51
+ $X2=3.115 $Y2=1.51
r66 20 21 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=2.98 $Y=1.51
+ $X2=1.865 $Y2=1.51
r67 17 40 6.50804 $w=5e-07 $l=3.55e-07 $layer=POLY_cond $X=1.695 $Y=1.395
+ $X2=1.695 $Y2=1.75
r68 17 19 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.695 $Y=1.395
+ $X2=1.695 $Y2=0.91
r69 13 40 1.65068 $w=5.84e-07 $l=2e-08 $layer=POLY_cond $X=1.675 $Y=1.75
+ $X2=1.695 $Y2=1.75
r70 13 38 62.726 $w=5.84e-07 $l=7.6e-07 $layer=POLY_cond $X=1.675 $Y=1.75
+ $X2=0.915 $Y2=1.75
r71 13 15 114.496 $w=5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.675 $Y=1.895
+ $X2=1.675 $Y2=2.965
r72 10 38 6.50804 $w=5e-07 $l=3.55e-07 $layer=POLY_cond $X=0.915 $Y=1.395
+ $X2=0.915 $Y2=1.75
r73 10 12 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.915 $Y=1.395
+ $X2=0.915 $Y2=0.91
r74 7 37 6.50804 $w=5e-07 $l=3.55e-07 $layer=POLY_cond $X=0.895 $Y=2.105
+ $X2=0.895 $Y2=1.75
r75 7 9 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.895 $Y=2.105 $X2=0.895
+ $Y2=2.965
r76 2 24 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.925
+ $Y=2.215 $X2=3.065 $Y2=2.34
r77 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.865 $X2=3.085 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_2%A 3 6 7 8 12 14 15
r24 12 15 22.1214 $w=5.2e-07 $l=2.15e-07 $layer=POLY_cond $X=2.685 $Y=1.89
+ $X2=2.685 $Y2=2.105
r25 12 14 50.9307 $w=5.2e-07 $l=4.95e-07 $layer=POLY_cond $X=2.685 $Y=1.89
+ $X2=2.685 $Y2=1.395
r26 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.89 $X2=2.61 $Y2=1.89
r27 8 13 1.00212 $w=3.43e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=1.947 $X2=2.61
+ $Y2=1.947
r28 7 13 15.0319 $w=3.43e-07 $l=4.5e-07 $layer=LI1_cond $X=2.16 $Y=1.947
+ $X2=2.61 $Y2=1.947
r29 6 14 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.695 $Y=1.075 $X2=2.695
+ $Y2=1.395
r30 3 15 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.675 $Y=2.59 $X2=2.675
+ $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_2%VPWR 1 2 7 10 20 28
r24 25 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.715 $Y=3.59
+ $X2=2.715 $Y2=3.59
r25 23 25 3.904 $w=1.248e-06 $l=4e-07 $layer=LI1_cond $X=2.175 $Y=3.19 $X2=2.175
+ $Y2=3.59
r26 20 23 7.8568 $w=1.248e-06 $l=8.05e-07 $layer=LI1_cond $X=2.175 $Y=2.385
+ $X2=2.175 $Y2=3.19
r27 14 17 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.195 $Y=3.63
+ $X2=0.915 $Y2=3.63
r28 13 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.915 $Y=3.59
+ $X2=0.915 $Y2=3.59
r29 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.195 $Y=3.59
+ $X2=0.195 $Y2=3.59
r30 10 13 16.3979 $w=9.28e-07 $l=1.25e-06 $layer=LI1_cond $X=0.555 $Y=2.34
+ $X2=0.555 $Y2=3.59
r31 7 28 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=1.635 $Y=3.63
+ $X2=2.715 $Y2=3.63
r32 7 17 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.635 $Y=3.63
+ $X2=0.915 $Y2=3.63
r33 7 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.635 $Y=3.59
+ $X2=1.635 $Y2=3.59
r34 2 23 300 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=2 $X=1.925
+ $Y=2.215 $X2=2.065 $Y2=3.19
r35 2 20 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=1.925
+ $Y=2.215 $X2=2.065 $Y2=2.385
r36 1 13 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.36
+ $Y=2.215 $X2=0.505 $Y2=3.59
r37 1 10 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.36
+ $Y=2.215 $X2=0.505 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_2%X 1 2 9 15 17 18 19
r26 18 19 21.8964 $w=2.28e-07 $l=4.37e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=1.157 $Y2=1.665
r27 17 18 24.051 $w=2.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.72 $Y2=1.665
r28 13 19 6.59134 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.305 $Y=1.55
+ $X2=1.2 $Y2=1.55
r29 13 15 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=1.305 $Y=1.55
+ $X2=1.305 $Y2=0.66
r30 9 11 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=1.285 $Y=2.34
+ $X2=1.285 $Y2=3.59
r31 7 19 6.59134 $w=1.7e-07 $l=2.69165e-07 $layer=LI1_cond $X=1.285 $Y=1.78
+ $X2=1.2 $Y2=1.55
r32 7 9 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.285 $Y=1.78
+ $X2=1.285 $Y2=2.34
r33 2 11 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=2.215 $X2=1.285 $Y2=3.59
r34 2 9 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=2.215 $X2=1.285 $Y2=2.34
r35 1 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.165
+ $Y=0.535 $X2=1.305 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_2%VGND 1 2 7 10 19 23
r24 25 27 4.88 $w=1.248e-06 $l=5e-07 $layer=LI1_cond $X=2.195 $Y=0.66 $X2=2.195
+ $Y2=1.16
r25 19 25 1.7568 $w=1.248e-06 $l=1.8e-07 $layer=LI1_cond $X=2.195 $Y=0.48
+ $X2=2.195 $Y2=0.66
r26 19 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.735 $Y=0.48
+ $X2=2.735 $Y2=0.48
r27 11 14 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.205 $Y=0.44
+ $X2=0.925 $Y2=0.44
r28 10 16 2.31158 $w=9.48e-07 $l=1.8e-07 $layer=LI1_cond $X=0.565 $Y=0.48
+ $X2=0.565 $Y2=0.66
r29 10 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.925 $Y=0.48
+ $X2=0.925 $Y2=0.48
r30 10 11 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.205 $Y=0.48
+ $X2=0.205 $Y2=0.48
r31 7 23 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=1.655 $Y=0.44
+ $X2=2.735 $Y2=0.44
r32 7 14 0.280251 $w=3.7e-07 $l=7.3e-07 $layer=MET1_cond $X=1.655 $Y=0.44
+ $X2=0.925 $Y2=0.44
r33 7 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.655 $Y=0.48
+ $X2=1.655 $Y2=0.48
r34 2 27 182 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.535 $X2=2.085 $Y2=1.16
r35 2 25 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.535 $X2=2.085 $Y2=0.66
r36 1 16 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.38
+ $Y=0.535 $X2=0.525 $Y2=0.66
.ends

