* NGSPICE file created from sky130_fd_sc_hvl__buf_4.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__buf_4 A VGND VNB VPB VPWR X
M1000 VGND a_149_81# X VNB nhv w=750000u l=500000u
+  ad=6.3375e+11p pd=6.19e+06u as=4.2e+11p ps=4.12e+06u
M1001 a_149_81# A VPWR VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=1.2675e+12p ps=1.069e+07u
M1002 VGND a_149_81# X VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_149_81# VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_149_81# X VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=8.4e+11p ps=7.12e+06u
M1005 X a_149_81# VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_149_81# X VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_149_81# A VGND VNB nhv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
M1008 X a_149_81# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_149_81# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends

