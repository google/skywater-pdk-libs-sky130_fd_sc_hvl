* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdlxtp_1 D GATE SCD SCE VGND VNB VPB VPWR Q
X0 a_1724_593# a_1678_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 a_1480_107# a_944_107# a_1636_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_489_107# SCE a_645_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_1678_81# a_1480_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 a_489_107# a_30_587# a_660_587# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X5 a_489_107# a_1214_107# a_1480_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 VGND D a_347_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_1480_107# a_1214_107# a_1724_593# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR a_944_107# a_1214_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X9 a_489_107# a_944_107# a_1480_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X10 VPWR SCE a_362_587# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 VPWR a_1480_107# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X12 VPWR GATE a_944_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X13 a_1636_107# a_1678_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 VGND GATE a_944_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_944_107# a_1214_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 a_660_587# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X17 a_645_107# SCD VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X18 a_30_587# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X19 a_30_587# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 a_347_107# a_30_587# a_489_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X21 a_1678_81# a_1480_107# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 VGND a_1480_107# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X23 a_362_587# D a_489_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
.ends
