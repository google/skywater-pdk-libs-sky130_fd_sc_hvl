# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hvl__sdfsbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  20.16000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.845000 2.305000 2.355000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.498750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.700000 0.495000 20.035000 1.325000 ;
        RECT 19.700000 2.355000 20.035000 3.435000 ;
        RECT 19.805000 1.325000 20.035000 2.355000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.611250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.405000 0.495000 17.785000 3.735000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 0.810000 3.690000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.495000 2.955000 1.665000 ;
        RECT 0.605000 1.665000 1.795000 2.165000 ;
        RECT 2.680000 1.095000 2.955000 1.495000 ;
        RECT 2.680000 1.665000 2.955000 1.765000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.205000 1.210000 12.355000 1.380000 ;
        RECT 12.185000 0.265000 14.170000 0.435000 ;
        RECT 12.185000 0.435000 12.355000 1.210000 ;
        RECT 14.000000 0.435000 14.170000 1.425000 ;
        RECT 14.000000 1.425000 14.845000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.380000 1.180000 4.710000 2.150000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.665000 0.365000 1.615000 0.915000 ;
    END
    PORT
      LAYER li1 ;
        RECT 10.545000 0.365000 11.495000 1.030000 ;
    END
    PORT
      LAYER li1 ;
        RECT 14.350000 0.365000 15.300000 1.245000 ;
    END
    PORT
      LAYER li1 ;
        RECT 16.240000 0.365000 17.190000 1.325000 ;
    END
    PORT
      LAYER li1 ;
        RECT 18.535000 0.365000 19.485000 1.325000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.870000 0.365000 4.760000 0.995000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.370000 0.365000 5.960000 1.020000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.410000 0.365000 9.360000 0.960000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 20.160000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 20.160000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 20.160000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 20.160000 4.155000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 20.160000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.640000 2.885000 1.590000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 10.955000 3.350000 11.905000 3.755000 ;
    END
    PORT
      LAYER li1 ;
        RECT 13.500000 2.875000 14.450000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 16.240000 2.195000 17.190000 3.735000 ;
    END
    PORT
      LAYER li1 ;
        RECT 18.535000 2.355000 19.485000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.415000 2.805000 4.305000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.695000 2.400000 5.865000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.615000 2.960000 9.565000 3.705000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 20.160000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.130000 0.495000  0.485000 1.095000 ;
      RECT  0.130000 1.095000  2.300000 1.315000 ;
      RECT  0.130000 1.315000  0.300000 2.535000 ;
      RECT  0.130000 2.535000  2.885000 2.705000 ;
      RECT  0.130000 2.705000  0.460000 3.305000 ;
      RECT  2.400000 2.885000  3.235000 3.055000 ;
      RECT  2.400000 3.055000  2.730000 3.305000 ;
      RECT  2.425000 0.495000  2.755000 0.745000 ;
      RECT  2.425000 0.745000  3.305000 0.915000 ;
      RECT  2.635000 2.015000  2.885000 2.535000 ;
      RECT  3.065000 2.455000  4.655000 2.625000 ;
      RECT  3.065000 2.625000  3.235000 2.885000 ;
      RECT  3.135000 0.915000  3.305000 2.455000 ;
      RECT  4.485000 2.625000  4.655000 3.635000 ;
      RECT  4.485000 3.635000  5.515000 3.805000 ;
      RECT  4.835000 2.805000  5.165000 3.455000 ;
      RECT  4.940000 0.515000  5.190000 1.700000 ;
      RECT  4.940000 1.700000  6.065000 1.870000 ;
      RECT  4.940000 1.870000  5.165000 2.805000 ;
      RECT  5.345000 2.050000  6.215000 2.220000 ;
      RECT  5.345000 2.220000  5.515000 3.635000 ;
      RECT  5.735000 1.200000  6.065000 1.700000 ;
      RECT  6.045000 2.220000  6.215000 3.390000 ;
      RECT  6.045000 3.390000  7.295000 3.560000 ;
      RECT  6.190000 0.265000  8.220000 0.435000 ;
      RECT  6.190000 0.435000  6.565000 1.020000 ;
      RECT  6.395000 1.020000  6.565000 2.290000 ;
      RECT  6.395000 2.290000  6.645000 3.210000 ;
      RECT  6.760000 0.615000  7.010000 1.060000 ;
      RECT  6.840000 1.060000  7.010000 2.740000 ;
      RECT  6.840000 2.740000  7.295000 3.390000 ;
      RECT  7.190000 0.435000  7.360000 2.290000 ;
      RECT  7.190000 2.290000  7.520000 2.560000 ;
      RECT  7.540000 0.640000  7.870000 1.060000 ;
      RECT  7.700000 1.060000  7.870000 1.910000 ;
      RECT  7.700000 1.910000 11.645000 2.080000 ;
      RECT  7.700000 2.080000  7.995000 3.240000 ;
      RECT  8.050000 0.435000  8.220000 1.150000 ;
      RECT  8.050000 1.150000  8.325000 1.560000 ;
      RECT  8.050000 1.560000 12.530000 1.730000 ;
      RECT  8.200000 2.290000  8.530000 2.610000 ;
      RECT  8.200000 2.610000  9.915000 2.780000 ;
      RECT  8.910000 1.140000  9.910000 1.380000 ;
      RECT  8.910000 2.260000 10.425000 2.430000 ;
      RECT  9.580000 0.515000  9.910000 1.140000 ;
      RECT  9.745000 2.780000  9.915000 3.170000 ;
      RECT  9.745000 3.170000 10.775000 3.340000 ;
      RECT 10.095000 2.430000 10.425000 2.990000 ;
      RECT 10.605000 3.000000 12.335000 3.170000 ;
      RECT 11.315000 2.080000 11.645000 2.555000 ;
      RECT 12.025000 2.125000 13.405000 2.295000 ;
      RECT 12.025000 2.295000 12.335000 3.000000 ;
      RECT 12.200000 1.730000 12.530000 1.875000 ;
      RECT 12.515000 2.525000 15.300000 2.695000 ;
      RECT 12.515000 2.695000 12.845000 3.755000 ;
      RECT 12.655000 0.615000 13.755000 0.785000 ;
      RECT 12.655000 0.785000 12.985000 1.325000 ;
      RECT 13.165000 1.415000 13.405000 2.125000 ;
      RECT 13.585000 0.785000 13.755000 1.825000 ;
      RECT 13.585000 1.825000 15.545000 1.995000 ;
      RECT 13.585000 1.995000 13.755000 2.525000 ;
      RECT 13.935000 2.175000 16.060000 2.345000 ;
      RECT 14.970000 2.695000 15.300000 3.175000 ;
      RECT 15.215000 1.425000 15.545000 1.825000 ;
      RECT 15.685000 2.345000 16.060000 2.675000 ;
      RECT 15.730000 0.825000 16.060000 2.175000 ;
      RECT 18.025000 0.825000 18.355000 1.505000 ;
      RECT 18.025000 1.505000 19.575000 1.675000 ;
      RECT 18.025000 1.675000 18.355000 3.185000 ;
      RECT 19.245000 1.675000 19.575000 2.175000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.670000  3.505000  0.840000 3.675000 ;
      RECT  0.695000  0.395000  0.865000 0.565000 ;
      RECT  1.030000  3.505000  1.200000 3.675000 ;
      RECT  1.055000  0.395000  1.225000 0.565000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.390000  3.505000  1.560000 3.675000 ;
      RECT  1.415000  0.395000  1.585000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.415000  3.505000  3.585000 3.675000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.775000  3.505000  3.945000 3.675000 ;
      RECT  3.870000  0.395000  4.040000 0.565000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.135000  3.505000  4.305000 3.675000 ;
      RECT  4.230000  0.395000  4.400000 0.565000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.590000  0.395000  4.760000 0.565000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.400000  0.395000  5.570000 0.565000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.695000  3.505000  5.865000 3.675000 ;
      RECT  5.760000  0.395000  5.930000 0.565000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.440000  0.395000  8.610000 0.565000 ;
      RECT  8.645000  3.505000  8.815000 3.675000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.800000  0.395000  8.970000 0.565000 ;
      RECT  9.005000  3.505000  9.175000 3.675000 ;
      RECT  9.160000  0.395000  9.330000 0.565000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.365000  3.505000  9.535000 3.675000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.575000  0.395000 10.745000 0.565000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.935000  0.395000 11.105000 0.565000 ;
      RECT 10.985000  3.505000 11.155000 3.675000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.295000  0.395000 11.465000 0.565000 ;
      RECT 11.345000  3.505000 11.515000 3.675000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 11.705000  3.505000 11.875000 3.675000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.530000  3.505000 13.700000 3.675000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.890000  3.505000 14.060000 3.675000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.250000  3.505000 14.420000 3.675000 ;
      RECT 14.380000  0.395000 14.550000 0.565000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.740000  0.395000 14.910000 0.565000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.100000  0.395000 15.270000 0.565000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.270000  0.395000 16.440000 0.565000 ;
      RECT 16.270000  3.505000 16.440000 3.675000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.630000  0.395000 16.800000 0.565000 ;
      RECT 16.630000  3.505000 16.800000 3.675000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 16.990000  0.395000 17.160000 0.565000 ;
      RECT 16.990000  3.505000 17.160000 3.675000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.985000 18.085000 4.155000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.985000 18.565000 4.155000 ;
      RECT 18.565000  0.395000 18.735000 0.565000 ;
      RECT 18.565000  3.505000 18.735000 3.675000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  3.985000 19.045000 4.155000 ;
      RECT 18.925000  0.395000 19.095000 0.565000 ;
      RECT 18.925000  3.505000 19.095000 3.675000 ;
      RECT 19.285000  0.395000 19.455000 0.565000 ;
      RECT 19.285000  3.505000 19.455000 3.675000 ;
      RECT 19.355000 -0.085000 19.525000 0.085000 ;
      RECT 19.355000  3.985000 19.525000 4.155000 ;
      RECT 19.835000 -0.085000 20.005000 0.085000 ;
      RECT 19.835000  3.985000 20.005000 4.155000 ;
  END
END sky130_fd_sc_hvl__sdfsbp_1
