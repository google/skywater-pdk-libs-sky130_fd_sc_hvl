* File: sky130_fd_sc_hvl__a21o_1.pxi.spice
* Created: Wed Sep  2 09:03:09 2020
* 
x_PM_SKY130_FD_SC_HVL__A21O_1%VNB N_VNB_M1001_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__A21O_1%VNB
x_PM_SKY130_FD_SC_HVL__A21O_1%VPB N_VPB_M1002_b VPB N_VPB_c_29_p VPB
+ PM_SKY130_FD_SC_HVL__A21O_1%VPB
x_PM_SKY130_FD_SC_HVL__A21O_1%A_83_283# N_A_83_283#_M1000_d N_A_83_283#_M1004_s
+ N_A_83_283#_M1002_g N_A_83_283#_M1001_g N_A_83_283#_c_79_n N_A_83_283#_c_80_n
+ N_A_83_283#_c_83_n N_A_83_283#_c_71_n N_A_83_283#_c_73_n N_A_83_283#_c_96_p
+ N_A_83_283#_c_74_n N_A_83_283#_c_86_n N_A_83_283#_c_75_n
+ PM_SKY130_FD_SC_HVL__A21O_1%A_83_283#
x_PM_SKY130_FD_SC_HVL__A21O_1%B1 N_B1_M1004_g N_B1_M1000_g B1 B1 B1 N_B1_c_134_n
+ PM_SKY130_FD_SC_HVL__A21O_1%B1
x_PM_SKY130_FD_SC_HVL__A21O_1%A1 N_A1_M1003_g N_A1_M1006_g A1 A1 N_A1_c_168_n
+ PM_SKY130_FD_SC_HVL__A21O_1%A1
x_PM_SKY130_FD_SC_HVL__A21O_1%A2 N_A2_M1007_g N_A2_M1005_g A2 N_A2_c_200_n
+ PM_SKY130_FD_SC_HVL__A21O_1%A2
x_PM_SKY130_FD_SC_HVL__A21O_1%X N_X_M1001_s N_X_M1002_s X X X X X X X
+ N_X_c_224_n X PM_SKY130_FD_SC_HVL__A21O_1%X
x_PM_SKY130_FD_SC_HVL__A21O_1%VPWR N_VPWR_M1002_d N_VPWR_M1003_d VPWR
+ N_VPWR_c_239_n N_VPWR_c_242_n N_VPWR_c_245_n PM_SKY130_FD_SC_HVL__A21O_1%VPWR
x_PM_SKY130_FD_SC_HVL__A21O_1%A_469_443# N_A_469_443#_M1004_d
+ N_A_469_443#_M1005_d N_A_469_443#_c_280_n N_A_469_443#_c_273_n
+ N_A_469_443#_c_287_n N_A_469_443#_c_276_n N_A_469_443#_c_277_n
+ PM_SKY130_FD_SC_HVL__A21O_1%A_469_443#
x_PM_SKY130_FD_SC_HVL__A21O_1%VGND N_VGND_M1001_d N_VGND_M1007_d VGND
+ N_VGND_c_302_n N_VGND_c_304_n N_VGND_c_306_n PM_SKY130_FD_SC_HVL__A21O_1%VGND
cc_1 N_VNB_M1001_b N_A_83_283#_M1001_g 0.0505391f $X=-0.33 $Y=-0.265 $X2=0.765
+ $Y2=0.91
cc_2 N_VNB_c_2_p N_A_83_283#_M1001_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.765 $Y2=0.91
cc_3 N_VNB_M1001_b N_A_83_283#_c_71_n 0.00864253f $X=-0.33 $Y=-0.265 $X2=2.515
+ $Y2=0.66
cc_4 N_VNB_c_2_p N_A_83_283#_c_71_n 6.32535e-19 $X=0.24 $Y=0 $X2=2.515 $Y2=0.66
cc_5 N_VNB_M1001_b N_A_83_283#_c_73_n 0.010476f $X=-0.33 $Y=-0.265 $X2=2.54
+ $Y2=1.93
cc_6 N_VNB_M1001_b N_A_83_283#_c_74_n 0.0639452f $X=-0.33 $Y=-0.265 $X2=0.73
+ $Y2=1.89
cc_7 N_VNB_M1001_b N_A_83_283#_c_75_n 9.64347e-19 $X=-0.33 $Y=-0.265 $X2=2.555
+ $Y2=1.325
cc_8 N_VNB_M1001_b N_B1_M1000_g 0.0472256f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=2.085
cc_9 N_VNB_c_2_p N_B1_M1000_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=2.085
cc_10 N_VNB_M1001_b B1 0.0220362f $X=-0.33 $Y=-0.265 $X2=0.765 $Y2=1.415
cc_11 N_VNB_M1001_b N_B1_c_134_n 0.0549302f $X=-0.33 $Y=-0.265 $X2=0.895
+ $Y2=2.015
cc_12 N_VNB_M1001_b N_A1_M1006_g 0.0423107f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=2.085
cc_13 N_VNB_c_2_p N_A1_M1006_g 9.54195e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=2.085
cc_14 N_VNB_M1001_b A1 0.00490455f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_15 N_VNB_M1001_b N_A1_c_168_n 0.0415612f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_16 N_VNB_M1001_b N_A2_M1007_g 0.0432009f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_17 N_VNB_M1001_b N_A2_c_200_n 0.0842466f $X=-0.33 $Y=-0.265 $X2=1.62
+ $Y2=2.015
cc_18 N_VNB_M1001_b X 0.04072f $X=-0.33 $Y=-0.265 $X2=0.665 $Y2=2.965
cc_19 N_VNB_M1001_b N_X_c_224_n 0.036911f $X=-0.33 $Y=-0.265 $X2=1.87 $Y2=2.015
cc_20 N_VNB_c_2_p N_X_c_224_n 8.15548e-19 $X=0.24 $Y=0 $X2=1.87 $Y2=2.015
cc_21 N_VNB_M1001_b N_VGND_c_302_n 0.0913413f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_22 N_VNB_c_2_p N_VGND_c_302_n 0.00456362f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_23 N_VNB_M1001_b N_VGND_c_304_n 0.101038f $X=-0.33 $Y=-0.265 $X2=2.555
+ $Y2=1.2
cc_24 N_VNB_c_2_p N_VGND_c_304_n 0.00371223f $X=0.24 $Y=0 $X2=2.555 $Y2=1.2
cc_25 N_VNB_M1001_b N_VGND_c_306_n 0.0796948f $X=-0.33 $Y=-0.265 $X2=2.555
+ $Y2=0.66
cc_26 N_VNB_c_2_p N_VGND_c_306_n 0.461892f $X=0.24 $Y=0 $X2=2.555 $Y2=0.66
cc_27 N_VPB_M1002_b N_A_83_283#_M1002_g 0.0459774f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=2.965
cc_28 VPB N_A_83_283#_M1002_g 0.00970178f $X=0 $Y=3.955 $X2=0.665 $Y2=2.965
cc_29 N_VPB_c_29_p N_A_83_283#_M1002_g 0.0152133f $X=4.08 $Y=4.07 $X2=0.665
+ $Y2=2.965
cc_30 N_VPB_M1002_b N_A_83_283#_c_79_n 0.0198329f $X=-0.33 $Y=1.885 $X2=1.62
+ $Y2=2.015
cc_31 N_VPB_M1002_b N_A_83_283#_c_80_n 0.00550143f $X=-0.33 $Y=1.885 $X2=1.705
+ $Y2=2.34
cc_32 VPB N_A_83_283#_c_80_n 8.01732e-19 $X=0 $Y=3.955 $X2=1.705 $Y2=2.34
cc_33 N_VPB_c_29_p N_A_83_283#_c_80_n 0.0130099f $X=4.08 $Y=4.07 $X2=1.705
+ $Y2=2.34
cc_34 N_VPB_M1002_b N_A_83_283#_c_83_n 0.00577499f $X=-0.33 $Y=1.885 $X2=2.455
+ $Y2=2.015
cc_35 N_VPB_M1002_b N_A_83_283#_c_73_n 9.62171e-19 $X=-0.33 $Y=1.885 $X2=2.54
+ $Y2=1.93
cc_36 N_VPB_M1002_b N_A_83_283#_c_74_n 0.0273841f $X=-0.33 $Y=1.885 $X2=0.73
+ $Y2=1.89
cc_37 N_VPB_M1002_b N_A_83_283#_c_86_n 0.00243745f $X=-0.33 $Y=1.885 $X2=1.745
+ $Y2=2.015
cc_38 N_VPB_M1002_b N_B1_M1004_g 0.0559675f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_39 VPB N_B1_M1004_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_40 N_VPB_c_29_p N_B1_M1004_g 0.0191024f $X=4.08 $Y=4.07 $X2=0 $Y2=0
cc_41 N_VPB_M1002_b N_B1_c_134_n 0.00459079f $X=-0.33 $Y=1.885 $X2=0.895
+ $Y2=2.015
cc_42 N_VPB_M1002_b N_A1_M1003_g 0.0499699f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_43 VPB N_A1_M1003_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_44 N_VPB_c_29_p N_A1_M1003_g 0.0158814f $X=4.08 $Y=4.07 $X2=0 $Y2=0
cc_45 N_VPB_M1002_b N_A1_c_168_n 0.00364711f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_46 N_VPB_M1002_b N_A2_M1005_g 0.0423641f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=2.085
cc_47 VPB N_A2_M1005_g 0.00970178f $X=0 $Y=3.955 $X2=0.665 $Y2=2.085
cc_48 N_VPB_c_29_p N_A2_M1005_g 0.0152133f $X=4.08 $Y=4.07 $X2=0.665 $Y2=2.085
cc_49 N_VPB_M1002_b N_A2_c_200_n 0.0418279f $X=-0.33 $Y=1.885 $X2=1.62 $Y2=2.015
cc_50 N_VPB_M1002_b X 0.0689552f $X=-0.33 $Y=1.885 $X2=0.665 $Y2=2.965
cc_51 VPB X 7.36921e-19 $X=0 $Y=3.955 $X2=0.665 $Y2=2.965
cc_52 N_VPB_c_29_p X 0.0120479f $X=4.08 $Y=4.07 $X2=0.665 $Y2=2.965
cc_53 N_VPB_M1002_b N_VPWR_c_239_n 0.027227f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_239_n 0.00339916f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_55 N_VPB_c_29_p N_VPWR_c_239_n 0.0459763f $X=4.08 $Y=4.07 $X2=0 $Y2=0
cc_56 N_VPB_M1002_b N_VPWR_c_242_n 0.00125033f $X=-0.33 $Y=1.885 $X2=1.745
+ $Y2=3.59
cc_57 VPB N_VPWR_c_242_n 0.00406397f $X=0 $Y=3.955 $X2=1.745 $Y2=3.59
cc_58 N_VPB_c_29_p N_VPWR_c_242_n 0.047451f $X=4.08 $Y=4.07 $X2=1.745 $Y2=3.59
cc_59 N_VPB_M1002_b N_VPWR_c_245_n 0.051634f $X=-0.33 $Y=1.885 $X2=2.515
+ $Y2=0.66
cc_60 VPB N_VPWR_c_245_n 0.458616f $X=0 $Y=3.955 $X2=2.515 $Y2=0.66
cc_61 N_VPB_c_29_p N_VPWR_c_245_n 0.0205091f $X=4.08 $Y=4.07 $X2=2.515 $Y2=0.66
cc_62 N_VPB_M1002_b N_A_469_443#_c_273_n 0.00124586f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=2.965
cc_63 VPB N_A_469_443#_c_273_n 0.00108855f $X=0 $Y=3.955 $X2=0.665 $Y2=2.965
cc_64 N_VPB_c_29_p N_A_469_443#_c_273_n 0.0171423f $X=4.08 $Y=4.07 $X2=0.665
+ $Y2=2.965
cc_65 N_VPB_M1002_b N_A_469_443#_c_276_n 0.0126063f $X=-0.33 $Y=1.885 $X2=0.765
+ $Y2=0.91
cc_66 N_VPB_M1002_b N_A_469_443#_c_277_n 0.0427929f $X=-0.33 $Y=1.885 $X2=1.62
+ $Y2=2.015
cc_67 VPB N_A_469_443#_c_277_n 7.36921e-19 $X=0 $Y=3.955 $X2=1.62 $Y2=2.015
cc_68 N_VPB_c_29_p N_A_469_443#_c_277_n 0.0120479f $X=4.08 $Y=4.07 $X2=1.62
+ $Y2=2.015
cc_69 N_A_83_283#_c_80_n N_B1_M1004_g 0.0487214f $X=1.705 $Y=2.34 $X2=0 $Y2=0
cc_70 N_A_83_283#_c_83_n N_B1_M1004_g 0.0384413f $X=2.455 $Y=2.015 $X2=0 $Y2=0
cc_71 N_A_83_283#_c_73_n N_B1_M1004_g 3.28406e-19 $X=2.54 $Y=1.93 $X2=0 $Y2=0
cc_72 N_A_83_283#_c_86_n N_B1_M1004_g 0.00500482f $X=1.745 $Y=2.015 $X2=0 $Y2=0
cc_73 N_A_83_283#_c_71_n N_B1_M1000_g 0.00134412f $X=2.515 $Y=0.66 $X2=0 $Y2=0
cc_74 N_A_83_283#_c_73_n N_B1_M1000_g 0.0101668f $X=2.54 $Y=1.93 $X2=0 $Y2=0
cc_75 N_A_83_283#_c_79_n B1 0.0397632f $X=1.62 $Y=2.015 $X2=0.24 $Y2=0
cc_76 N_A_83_283#_c_83_n B1 0.0269463f $X=2.455 $Y=2.015 $X2=0.24 $Y2=0
cc_77 N_A_83_283#_c_73_n B1 0.0185907f $X=2.54 $Y=1.93 $X2=0.24 $Y2=0
cc_78 N_A_83_283#_c_96_p B1 0.00186129f $X=0.73 $Y=1.89 $X2=0.24 $Y2=0
cc_79 N_A_83_283#_c_74_n B1 0.012296f $X=0.73 $Y=1.89 $X2=0.24 $Y2=0
cc_80 N_A_83_283#_c_86_n B1 0.0205804f $X=1.745 $Y=2.015 $X2=0.24 $Y2=0
cc_81 N_A_83_283#_c_83_n N_B1_c_134_n 0.00147531f $X=2.455 $Y=2.015 $X2=4.08
+ $Y2=0
cc_82 N_A_83_283#_c_83_n N_A1_M1003_g 0.00601391f $X=2.455 $Y=2.015 $X2=0 $Y2=0
cc_83 N_A_83_283#_c_71_n N_A1_M1006_g 0.0121186f $X=2.515 $Y=0.66 $X2=0 $Y2=0
cc_84 N_A_83_283#_c_73_n N_A1_M1006_g 0.00231767f $X=2.54 $Y=1.93 $X2=0 $Y2=0
cc_85 N_A_83_283#_c_75_n N_A1_M1006_g 0.00360345f $X=2.555 $Y=1.325 $X2=0 $Y2=0
cc_86 N_A_83_283#_c_73_n A1 0.0250925f $X=2.54 $Y=1.93 $X2=0.24 $Y2=0
cc_87 N_A_83_283#_c_73_n N_A1_c_168_n 0.00789878f $X=2.54 $Y=1.93 $X2=0 $Y2=0
cc_88 N_A_83_283#_c_75_n N_A1_c_168_n 0.00158354f $X=2.555 $Y=1.325 $X2=0 $Y2=0
cc_89 N_A_83_283#_c_71_n N_A2_M1007_g 2.95342e-19 $X=2.515 $Y=0.66 $X2=0 $Y2=0
cc_90 N_A_83_283#_M1001_g X 0.00372574f $X=0.765 $Y=0.91 $X2=0 $Y2=0
cc_91 N_A_83_283#_c_96_p X 0.0251954f $X=0.73 $Y=1.89 $X2=0 $Y2=0
cc_92 N_A_83_283#_c_74_n X 0.0354347f $X=0.73 $Y=1.89 $X2=0 $Y2=0
cc_93 N_A_83_283#_M1001_g N_X_c_224_n 0.00491044f $X=0.765 $Y=0.91 $X2=2.16
+ $Y2=0.058
cc_94 N_A_83_283#_M1002_g N_VPWR_c_239_n 0.0740873f $X=0.665 $Y=2.965 $X2=0.24
+ $Y2=0
cc_95 N_A_83_283#_c_79_n N_VPWR_c_239_n 0.0409507f $X=1.62 $Y=2.015 $X2=0.24
+ $Y2=0
cc_96 N_A_83_283#_c_80_n N_VPWR_c_239_n 0.115906f $X=1.705 $Y=2.34 $X2=0.24
+ $Y2=0
cc_97 N_A_83_283#_c_96_p N_VPWR_c_239_n 0.0253593f $X=0.73 $Y=1.89 $X2=0.24
+ $Y2=0
cc_98 N_A_83_283#_c_74_n N_VPWR_c_239_n 5.72841e-19 $X=0.73 $Y=1.89 $X2=0.24
+ $Y2=0
cc_99 N_A_83_283#_M1004_s N_VPWR_c_245_n 0.00254395f $X=1.56 $Y=2.215 $X2=0
+ $Y2=0
cc_100 N_A_83_283#_M1002_g N_VPWR_c_245_n 0.00914225f $X=0.665 $Y=2.965 $X2=0
+ $Y2=0
cc_101 N_A_83_283#_c_80_n N_VPWR_c_245_n 0.0333758f $X=1.705 $Y=2.34 $X2=0 $Y2=0
cc_102 N_A_83_283#_c_80_n N_A_469_443#_c_280_n 0.00602838f $X=1.705 $Y=2.34
+ $X2=0 $Y2=0
cc_103 N_A_83_283#_c_83_n N_A_469_443#_c_280_n 0.0204505f $X=2.455 $Y=2.015
+ $X2=0 $Y2=0
cc_104 N_A_83_283#_c_80_n N_A_469_443#_c_273_n 0.0390137f $X=1.705 $Y=2.34 $X2=0
+ $Y2=0
cc_105 N_A_83_283#_M1001_g N_VGND_c_302_n 0.0626596f $X=0.765 $Y=0.91 $X2=0.24
+ $Y2=0
cc_106 N_A_83_283#_c_79_n N_VGND_c_302_n 0.00562458f $X=1.62 $Y=2.015 $X2=0.24
+ $Y2=0
cc_107 N_A_83_283#_c_71_n N_VGND_c_302_n 0.0363808f $X=2.515 $Y=0.66 $X2=0.24
+ $Y2=0
cc_108 N_A_83_283#_c_96_p N_VGND_c_302_n 0.0102284f $X=0.73 $Y=1.89 $X2=0.24
+ $Y2=0
cc_109 N_A_83_283#_c_71_n N_VGND_c_304_n 0.0602248f $X=2.515 $Y=0.66 $X2=2.16
+ $Y2=0.058
cc_110 N_A_83_283#_M1000_d N_VGND_c_306_n 0.00221032f $X=2.375 $Y=0.535 $X2=0
+ $Y2=0
cc_111 N_A_83_283#_M1001_g N_VGND_c_306_n 0.00877352f $X=0.765 $Y=0.91 $X2=0
+ $Y2=0
cc_112 N_A_83_283#_c_71_n N_VGND_c_306_n 0.0243019f $X=2.515 $Y=0.66 $X2=0 $Y2=0
cc_113 N_B1_M1004_g N_A1_M1003_g 0.0246535f $X=2.095 $Y=2.965 $X2=0 $Y2=0
cc_114 N_B1_M1000_g N_A1_M1006_g 0.0169538f $X=2.125 $Y=0.91 $X2=0 $Y2=0
cc_115 N_B1_c_134_n N_A1_c_168_n 0.0248252f $X=2.03 $Y=1.63 $X2=0 $Y2=0
cc_116 N_B1_M1004_g N_VPWR_c_239_n 0.00310247f $X=2.095 $Y=2.965 $X2=0.24 $Y2=0
cc_117 N_B1_M1004_g N_VPWR_c_242_n 4.09987e-19 $X=2.095 $Y=2.965 $X2=0 $Y2=0
cc_118 N_B1_M1004_g N_VPWR_c_245_n 0.0270666f $X=2.095 $Y=2.965 $X2=0 $Y2=0
cc_119 N_B1_M1004_g N_A_469_443#_c_280_n 0.00496865f $X=2.095 $Y=2.965 $X2=0
+ $Y2=0
cc_120 N_B1_M1004_g N_A_469_443#_c_273_n 0.033158f $X=2.095 $Y=2.965 $X2=0 $Y2=0
cc_121 N_B1_M1000_g N_VGND_c_302_n 0.0738326f $X=2.125 $Y=0.91 $X2=0.24 $Y2=0
cc_122 B1 N_VGND_c_302_n 0.0934977f $X=2.075 $Y=1.58 $X2=0.24 $Y2=0
cc_123 N_B1_c_134_n N_VGND_c_302_n 9.0518e-19 $X=2.03 $Y=1.63 $X2=0.24 $Y2=0
cc_124 N_B1_M1000_g N_VGND_c_304_n 5.31178e-19 $X=2.125 $Y=0.91 $X2=2.16
+ $Y2=0.058
cc_125 N_B1_M1000_g N_VGND_c_306_n 0.00778503f $X=2.125 $Y=0.91 $X2=0 $Y2=0
cc_126 N_A1_M1006_g N_A2_M1007_g 0.0512415f $X=2.905 $Y=0.91 $X2=0 $Y2=0
cc_127 N_A1_M1003_g N_A2_M1005_g 0.0350141f $X=2.875 $Y=2.965 $X2=0 $Y2=0
cc_128 A1 A2 0.0249551f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A1_M1003_g N_A2_c_200_n 0.0122151f $X=2.875 $Y=2.965 $X2=0 $Y2=0
cc_130 A1 N_A2_c_200_n 0.0319267f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_131 N_A1_c_168_n N_A2_c_200_n 0.0512415f $X=2.97 $Y=1.67 $X2=0 $Y2=0
cc_132 N_A1_M1003_g N_VPWR_c_242_n 0.0524065f $X=2.875 $Y=2.965 $X2=0 $Y2=0
cc_133 N_A1_M1003_g N_VPWR_c_245_n 0.0101395f $X=2.875 $Y=2.965 $X2=0 $Y2=0
cc_134 N_A1_M1003_g N_A_469_443#_c_280_n 0.00163016f $X=2.875 $Y=2.965 $X2=0
+ $Y2=0
cc_135 N_A1_M1003_g N_A_469_443#_c_273_n 0.0263827f $X=2.875 $Y=2.965 $X2=0
+ $Y2=0
cc_136 N_A1_M1003_g N_A_469_443#_c_287_n 0.035834f $X=2.875 $Y=2.965 $X2=0.24
+ $Y2=0
cc_137 A1 N_A_469_443#_c_287_n 0.0293072f $X=3.515 $Y=1.58 $X2=0.24 $Y2=0
cc_138 N_A1_M1006_g N_VGND_c_302_n 7.32521e-19 $X=2.905 $Y=0.91 $X2=0.24 $Y2=0
cc_139 N_A1_M1006_g N_VGND_c_304_n 0.0548534f $X=2.905 $Y=0.91 $X2=2.16
+ $Y2=0.058
cc_140 A1 N_VGND_c_304_n 0.066717f $X=3.515 $Y=1.58 $X2=2.16 $Y2=0.058
cc_141 N_A1_M1006_g N_VGND_c_306_n 0.0108828f $X=2.905 $Y=0.91 $X2=0 $Y2=0
cc_142 N_A2_M1005_g N_VPWR_c_242_n 0.0573033f $X=3.655 $Y=2.965 $X2=0 $Y2=0
cc_143 N_A2_M1005_g N_VPWR_c_245_n 0.00853278f $X=3.655 $Y=2.965 $X2=0 $Y2=0
cc_144 N_A2_M1005_g N_A_469_443#_c_287_n 0.0360481f $X=3.655 $Y=2.965 $X2=0.24
+ $Y2=0
cc_145 A2 N_A_469_443#_c_287_n 0.00125889f $X=3.995 $Y=1.58 $X2=0.24 $Y2=0
cc_146 N_A2_M1005_g N_A_469_443#_c_276_n 9.14118e-19 $X=3.655 $Y=2.965 $X2=0
+ $Y2=0
cc_147 A2 N_A_469_443#_c_276_n 0.0113262f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A2_c_200_n N_A_469_443#_c_276_n 0.00831897f $X=4.03 $Y=1.67 $X2=0 $Y2=0
cc_149 N_A2_M1005_g N_A_469_443#_c_277_n 0.00179384f $X=3.655 $Y=2.965 $X2=0
+ $Y2=0
cc_150 N_A2_M1007_g N_VGND_c_304_n 0.0775946f $X=3.615 $Y=0.91 $X2=2.16
+ $Y2=0.058
cc_151 A2 N_VGND_c_304_n 0.0221192f $X=3.995 $Y=1.58 $X2=2.16 $Y2=0.058
cc_152 N_A2_c_200_n N_VGND_c_304_n 0.00976072f $X=4.03 $Y=1.67 $X2=2.16
+ $Y2=0.058
cc_153 X N_VPWR_c_239_n 0.0607971f $X=0.155 $Y=1.21 $X2=0.24 $Y2=0
cc_154 N_X_M1002_s N_VPWR_c_245_n 0.00221032f $X=0.15 $Y=2.215 $X2=0 $Y2=0
cc_155 X N_VPWR_c_245_n 0.0341921f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_156 N_X_c_224_n N_VGND_c_302_n 0.0364892f $X=0.375 $Y=0.66 $X2=0.24 $Y2=0
cc_157 N_X_M1001_s N_VGND_c_306_n 0.00221032f $X=0.23 $Y=0.535 $X2=0 $Y2=0
cc_158 N_X_c_224_n N_VGND_c_306_n 0.0350118f $X=0.375 $Y=0.66 $X2=0 $Y2=0
cc_159 N_VPWR_c_245_n N_A_469_443#_M1005_d 0.00221032f $X=3.665 $Y=3.59 $X2=0
+ $Y2=0
cc_160 N_VPWR_c_242_n N_A_469_443#_c_273_n 0.0808879f $X=3.265 $Y=2.715 $X2=0.24
+ $Y2=4.07
cc_161 N_VPWR_c_245_n N_A_469_443#_c_273_n 0.04111f $X=3.665 $Y=3.59 $X2=0.24
+ $Y2=4.07
cc_162 N_VPWR_M1003_d N_A_469_443#_c_287_n 0.00462521f $X=3.125 $Y=2.215 $X2=0
+ $Y2=0
cc_163 N_VPWR_c_242_n N_A_469_443#_c_287_n 0.0614519f $X=3.265 $Y=2.715 $X2=0
+ $Y2=0
cc_164 N_VPWR_c_242_n N_A_469_443#_c_277_n 0.0467807f $X=3.265 $Y=2.715 $X2=4.08
+ $Y2=4.07
cc_165 N_VPWR_c_245_n N_A_469_443#_c_277_n 0.0341921f $X=3.665 $Y=3.59 $X2=4.08
+ $Y2=4.07
