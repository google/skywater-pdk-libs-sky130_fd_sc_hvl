* File: sky130_fd_sc_hvl__lsbufhv2lv_1.pex.spice
* Created: Fri Aug 28 09:36:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%VNB 9 11 12 23 35 43 50
r70 35 50 2.30978 $w=2.3e-07 $l=3.6e-06 $layer=MET1_cond $X=7.92 $Y=8.14
+ $X2=4.32 $Y2=8.14
r71 23 43 2.30978 $w=2.3e-07 $l=3.6e-06 $layer=MET1_cond $X=7.92 $Y=0 $X2=4.32
+ $Y2=0
r72 12 50 0.153985 $w=2.3e-07 $l=2.4e-07 $layer=MET1_cond $X=4.08 $Y=8.14
+ $X2=4.32 $Y2=8.14
r73 12 29 2.46376 $w=2.3e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=8.14
+ $X2=0.24 $Y2=8.14
r74 11 43 0.153985 $w=2.3e-07 $l=2.4e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.32
+ $Y2=0
r75 11 17 2.46376 $w=2.3e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=0.24
+ $Y2=0
r76 9 35 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=7.92 $Y=8.14
+ $X2=7.92 $Y2=8.14
r77 9 29 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=0.24 $Y=8.14
+ $X2=0.24 $Y2=8.14
r78 9 23 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r79 9 17 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%VPB 7 8 11 14 20 21 29
r55 21 29 2.30978 $w=2.3e-07 $l=3.6e-06 $layer=MET1_cond $X=7.92 $Y=4.07
+ $X2=4.32 $Y2=4.07
r56 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=4.07
+ $X2=7.92 $Y2=4.07
r57 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=4.07
+ $X2=0.72 $Y2=4.07
r58 11 29 0.153985 $w=2.3e-07 $l=2.4e-07 $layer=MET1_cond $X=4.08 $Y=4.07
+ $X2=4.32 $Y2=4.07
r59 11 15 2.15579 $w=2.3e-07 $l=3.36e-06 $layer=MET1_cond $X=4.08 $Y=4.07
+ $X2=0.72 $Y2=4.07
r60 8 20 91 $w=1.7e-07 $l=6.3107e-07 $layer=licon1_NTAP_notbjt $count=2 $X=7.33
+ $Y=3.985 $X2=7.92 $Y2=4.07
r61 7 14 91 $w=1.7e-07 $l=7.61315e-07 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=0.72 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%LVPWR 1 2 10 14 16 18 22 29 36
r69 29 36 0.179425 $w=2.85e-07 $l=3.6e-07 $layer=MET1_cond $X=4.605 $Y=3.162
+ $X2=4.245 $Y2=3.162
r70 25 31 7.15962 $w=8.52e-07 $l=5e-07 $layer=LI1_cond $X=4.265 $Y=3.08
+ $X2=4.265 $Y2=3.58
r71 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.605 $Y=3.19
+ $X2=4.605 $Y2=3.19
r72 25 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.245 $Y=3.19
+ $X2=4.245 $Y2=3.19
r73 22 36 0.0822366 $w=2.85e-07 $l=1.65e-07 $layer=MET1_cond $X=4.08 $Y=3.162
+ $X2=4.245 $Y2=3.162
r74 18 20 35.427 $w=2.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.265 $Y=4.42
+ $X2=4.265 $Y2=5.25
r75 16 31 13.4189 $w=8.52e-07 $l=5.05e-07 $layer=LI1_cond $X=4.265 $Y=4.085
+ $X2=4.265 $Y2=3.58
r76 16 18 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.265 $Y=4.085
+ $X2=4.265 $Y2=4.42
r77 12 25 6.25931 $w=8.52e-07 $l=5e-09 $layer=LI1_cond $X=4.265 $Y=3.075
+ $X2=4.265 $Y2=3.08
r78 12 14 35.2135 $w=2.68e-07 $l=8.25e-07 $layer=LI1_cond $X=4.265 $Y=3.075
+ $X2=4.265 $Y2=2.25
r79 10 31 60.6667 $w=1.7e-07 $l=9.46546e-07 $layer=licon1_NTAP_notbjt $count=3
+ $X=3.71 $Y=3.495 $X2=4.615 $Y2=3.58
r80 10 31 60.6667 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=3
+ $X=3.71 $Y=3.495 $X2=3.915 $Y2=3.58
r81 2 20 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=4.125
+ $Y=4.275 $X2=4.265 $Y2=5.25
r82 2 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.125
+ $Y=4.275 $X2=4.265 $Y2=4.42
r83 1 25 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=4.125
+ $Y=2.105 $X2=4.265 $Y2=3.08
r84 1 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.125
+ $Y=2.105 $X2=4.265 $Y2=2.25
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A_30_1337# 1 2 7 9 12 13 15 16 18 20
+ 21 23 24 26 28 32 33 36 38 39 40 43 48 49 52
r98 51 53 4.88897 $w=7.98e-07 $l=3.27e-07 $layer=LI1_cond $X=1.35 $Y=6.07
+ $X2=1.35 $Y2=6.397
r99 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.61
+ $Y=6.07 $X2=1.61 $Y2=6.07
r100 48 51 5.3076 $w=7.98e-07 $l=3.55e-07 $layer=LI1_cond $X=1.35 $Y=5.715
+ $X2=1.35 $Y2=6.07
r101 48 49 7.8342 $w=7.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=5.715
+ $X2=1.35 $Y2=5.55
r102 45 49 101.456 $w=2.78e-07 $l=2.465e-06 $layer=LI1_cond $X=1.61 $Y=3.085
+ $X2=1.61 $Y2=5.55
r103 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.135
+ $Y=2.96 $X2=1.135 $Y2=2.96
r104 40 45 6.84494 $w=2.5e-07 $l=1.92614e-07 $layer=LI1_cond $X=1.47 $Y=2.96
+ $X2=1.61 $Y2=3.085
r105 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.47 $Y=2.96
+ $X2=1.135 $Y2=2.96
r106 38 53 5.52441 $w=3.55e-07 $l=4e-07 $layer=LI1_cond $X=0.95 $Y=6.397
+ $X2=1.35 $Y2=6.397
r107 38 39 17.2055 $w=3.53e-07 $l=5.3e-07 $layer=LI1_cond $X=0.95 $Y=6.397
+ $X2=0.42 $Y2=6.397
r108 34 39 7.08698 $w=3.55e-07 $l=2.32237e-07 $layer=LI1_cond $X=0.295 $Y=6.575
+ $X2=0.42 $Y2=6.397
r109 34 36 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=0.295 $Y=6.575
+ $X2=0.295 $Y2=6.895
r110 31 52 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=1.61 $Y=6.46
+ $X2=1.61 $Y2=6.07
r111 31 32 8.21244 $w=4.15e-07 $l=1.16619e-07 $layer=POLY_cond $X=1.61 $Y=6.46
+ $X2=1.695 $Y2=6.535
r112 30 43 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.935 $Y=2.96
+ $X2=1.135 $Y2=2.96
r113 29 30 6.42064 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.685 $Y=2.96
+ $X2=0.935 $Y2=2.96
r114 26 28 43.38 $w=5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.255 $Y=6.61 $X2=3.255
+ $Y2=7.06
r115 25 33 80.3333 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.725 $Y=6.535
+ $X2=2.475 $Y2=6.535
r116 24 26 38.6381 $w=1.5e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.005 $Y=6.535
+ $X2=3.255 $Y2=6.61
r117 24 25 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.005 $Y=6.535
+ $X2=2.725 $Y2=6.535
r118 21 33 7.23 $w=5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.475 $Y=6.61 $X2=2.475
+ $Y2=6.535
r119 21 23 43.38 $w=5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.475 $Y=6.61 $X2=2.475
+ $Y2=7.06
r120 18 33 7.23 $w=5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.475 $Y=6.46 $X2=2.475
+ $Y2=6.535
r121 18 20 43.38 $w=5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.475 $Y=6.46 $X2=2.475
+ $Y2=6.01
r122 17 32 20.4038 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.945 $Y=6.535
+ $X2=1.695 $Y2=6.535
r123 16 33 80.3333 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.225 $Y=6.535
+ $X2=2.475 $Y2=6.535
r124 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.225 $Y=6.535
+ $X2=1.945 $Y2=6.535
r125 13 32 8.21244 $w=4.15e-07 $l=7.5e-08 $layer=POLY_cond $X=1.695 $Y=6.61
+ $X2=1.695 $Y2=6.535
r126 13 15 43.38 $w=5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.695 $Y=6.61 $X2=1.695
+ $Y2=7.06
r127 9 12 126.267 $w=5e-07 $l=1.18e-06 $layer=POLY_cond $X=0.685 $Y=1.245
+ $X2=0.685 $Y2=2.425
r128 7 29 45.6147 $w=5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.685 $Y=2.515
+ $X2=0.685 $Y2=2.96
r129 7 12 9.63053 $w=5e-07 $l=9e-08 $layer=POLY_cond $X=0.685 $Y=2.515 $X2=0.685
+ $Y2=2.425
r130 2 48 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=5.505 $X2=1.075 $Y2=5.715
r131 1 36 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=6.685 $X2=0.295 $Y2=6.895
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A 1 3 5 9 10 11 12 16
r27 12 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.135
+ $Y=5.035 $X2=1.135 $Y2=5.035
r28 11 12 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.72 $Y=5.035
+ $X2=1.135 $Y2=5.035
r29 10 16 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.935 $Y=5.035
+ $X2=1.135 $Y2=5.035
r30 7 10 26.9851 $w=3.3e-07 $l=2.29063e-07 $layer=POLY_cond $X=0.782 $Y=5.2
+ $X2=0.935 $Y2=5.035
r31 7 9 34.4187 $w=3.05e-07 $l=1.75e-07 $layer=POLY_cond $X=0.782 $Y=5.2
+ $X2=0.782 $Y2=5.375
r32 3 5 126.267 $w=5e-07 $l=1.18e-06 $layer=POLY_cond $X=0.685 $Y=5.715
+ $X2=0.685 $Y2=6.895
r33 1 9 34.832 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.685 $Y=5.625 $X2=0.685
+ $Y2=5.375
r34 1 3 9.63053 $w=5e-07 $l=9e-08 $layer=POLY_cond $X=0.685 $Y=5.625 $X2=0.685
+ $Y2=5.715
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A_30_207# 1 2 9 11 13 17 19 23 25 26
+ 29 34 36
r51 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.61
+ $Y=1.73 $X2=1.61 $Y2=1.73
r52 34 36 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=1.597 $Y=1.73
+ $X2=1.61 $Y2=1.73
r53 33 34 18.2296 $w=3.28e-07 $l=5.22e-07 $layer=LI1_cond $X=1.075 $Y=1.73
+ $X2=1.597 $Y2=1.73
r54 27 33 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=1.075 $Y=1.895
+ $X2=1.075 $Y2=1.73
r55 27 29 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=1.075 $Y=1.895
+ $X2=1.075 $Y2=2.425
r56 25 33 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.95 $Y=1.73
+ $X2=1.075 $Y2=1.73
r57 25 26 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.95 $Y=1.73
+ $X2=0.42 $Y2=1.73
r58 21 26 6.98653 $w=3.3e-07 $l=2.18746e-07 $layer=LI1_cond $X=0.295 $Y=1.565
+ $X2=0.42 $Y2=1.73
r59 21 23 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=0.295 $Y=1.565
+ $X2=0.295 $Y2=1.245
r60 17 19 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.475 $Y=2.5
+ $X2=2.475 $Y2=3.55
r61 11 37 105.552 $w=3.95e-07 $l=8.65e-07 $layer=POLY_cond $X=2.475 $Y=1.942
+ $X2=1.61 $Y2=1.942
r62 11 17 55.6431 $w=5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.475 $Y=1.98
+ $X2=2.475 $Y2=2.5
r63 11 13 60.9934 $w=5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.475 $Y=1.65
+ $X2=2.475 $Y2=1.08
r64 9 37 60.9934 $w=5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.695 $Y=1.08 $X2=1.695
+ $Y2=1.65
r65 2 29 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=2.215 $X2=1.075 $Y2=2.425
r66 1 23 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=1.035 $X2=0.295 $Y2=1.245
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A_389_1337# 1 2 3 4 15 19 23 24 26 29
+ 31 35 38 41 42 45
r74 43 45 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=4.695 $Y=2.78
+ $X2=5.045 $Y2=2.78
r75 40 45 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.045 $Y=2.905
+ $X2=5.045 $Y2=2.78
r76 40 41 124.003 $w=2.48e-07 $l=2.69e-06 $layer=LI1_cond $X=5.045 $Y=2.905
+ $X2=5.045 $Y2=5.595
r77 36 43 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=4.695 $Y=2.655
+ $X2=4.695 $Y2=2.78
r78 36 38 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=4.695 $Y=2.655
+ $X2=4.695 $Y2=2.25
r79 35 47 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=4.22 $Y=5.72
+ $X2=4.05 $Y2=5.72
r80 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.22
+ $Y=5.72 $X2=4.22 $Y2=5.72
r81 32 42 1.88208 $w=2.5e-07 $l=2.6e-07 $layer=LI1_cond $X=3.81 $Y=5.72 $X2=3.55
+ $Y2=5.72
r82 32 34 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=3.81 $Y=5.72
+ $X2=4.22 $Y2=5.72
r83 31 41 6.81649 $w=2.5e-07 $l=1.76777e-07 $layer=LI1_cond $X=4.92 $Y=5.72
+ $X2=5.045 $Y2=5.595
r84 31 34 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=4.92 $Y=5.72 $X2=4.22
+ $Y2=5.72
r85 27 42 4.55795 $w=2.9e-07 $l=1.65831e-07 $layer=LI1_cond $X=3.645 $Y=5.845
+ $X2=3.55 $Y2=5.72
r86 27 29 34.3987 $w=3.28e-07 $l=9.85e-07 $layer=LI1_cond $X=3.645 $Y=5.845
+ $X2=3.645 $Y2=6.83
r87 26 42 4.55795 $w=2.9e-07 $l=1.8735e-07 $layer=LI1_cond $X=3.415 $Y=5.595
+ $X2=3.55 $Y2=5.72
r88 25 26 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=3.415 $Y=5.445
+ $X2=3.415 $Y2=5.595
r89 23 25 6.81649 $w=2.5e-07 $l=1.76777e-07 $layer=LI1_cond $X=3.29 $Y=5.32
+ $X2=3.415 $Y2=5.445
r90 23 24 47.9416 $w=2.48e-07 $l=1.04e-06 $layer=LI1_cond $X=3.29 $Y=5.32
+ $X2=2.25 $Y2=5.32
r91 19 21 36.6686 $w=3.28e-07 $l=1.05e-06 $layer=LI1_cond $X=2.085 $Y=5.78
+ $X2=2.085 $Y2=6.83
r92 17 24 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=2.085 $Y=5.445
+ $X2=2.25 $Y2=5.32
r93 17 19 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.085 $Y=5.445
+ $X2=2.085 $Y2=5.78
r94 13 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.05 $Y=5.555
+ $X2=4.05 $Y2=5.72
r95 13 15 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=4.05 $Y=5.555
+ $X2=4.05 $Y2=4.835
r96 4 38 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.555
+ $Y=2.105 $X2=4.695 $Y2=2.25
r97 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.505
+ $Y=6.685 $X2=3.645 $Y2=6.83
r98 2 19 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.96
+ $Y=5.635 $X2=2.085 $Y2=5.78
r99 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=6.685 $X2=2.085 $Y2=6.83
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A_389_141# 1 2 3 4 14 15 16 19 23 27
+ 30 34 40 41 48 50 54
r84 48 53 4.04821 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=3.835 $Y=4.595
+ $X2=3.835 $Y2=4.425
r85 48 50 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=3.835 $Y=4.595
+ $X2=3.835 $Y2=5.25
r86 47 54 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.335 $Y=4.43
+ $X2=3.17 $Y2=4.43
r87 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.335
+ $Y=4.43 $X2=3.335 $Y2=4.43
r88 44 54 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.995 $Y=4.43
+ $X2=3.17 $Y2=4.43
r89 43 46 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.995 $Y=4.425
+ $X2=3.335 $Y2=4.425
r90 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.995
+ $Y=4.43 $X2=2.995 $Y2=4.43
r91 41 43 25.2521 $w=3.38e-07 $l=7.45e-07 $layer=LI1_cond $X=2.25 $Y=4.425
+ $X2=2.995 $Y2=4.425
r92 40 53 2.97663 $w=3.4e-07 $l=1.25e-07 $layer=LI1_cond $X=3.71 $Y=4.425
+ $X2=3.835 $Y2=4.425
r93 40 46 12.7108 $w=3.38e-07 $l=3.75e-07 $layer=LI1_cond $X=3.71 $Y=4.425
+ $X2=3.335 $Y2=4.425
r94 37 39 36.6686 $w=3.28e-07 $l=1.05e-06 $layer=LI1_cond $X=2.085 $Y=2.27
+ $X2=2.085 $Y2=3.32
r95 34 37 49.59 $w=3.28e-07 $l=1.42e-06 $layer=LI1_cond $X=2.085 $Y=0.85
+ $X2=2.085 $Y2=2.27
r96 32 41 6.81847 $w=3.4e-07 $l=2.38642e-07 $layer=LI1_cond $X=2.085 $Y=4.255
+ $X2=2.25 $Y2=4.425
r97 32 39 32.6526 $w=3.28e-07 $l=9.35e-07 $layer=LI1_cond $X=2.085 $Y=4.255
+ $X2=2.085 $Y2=3.32
r98 29 30 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.05 $Y=1.8 $X2=4.48
+ $Y2=1.8
r99 25 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.48 $Y=1.965
+ $X2=4.48 $Y2=1.8
r100 25 27 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=4.48 $Y=1.965
+ $X2=4.48 $Y2=2.665
r101 21 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.05 $Y=1.965
+ $X2=4.05 $Y2=1.8
r102 21 23 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=4.05 $Y=1.965
+ $X2=4.05 $Y2=2.665
r103 17 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.05 $Y=1.635
+ $X2=4.05 $Y2=1.8
r104 17 19 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.05 $Y=1.635
+ $X2=4.05 $Y2=1.125
r105 15 29 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.975 $Y=1.8
+ $X2=4.05 $Y2=1.8
r106 15 16 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=3.975 $Y=1.8
+ $X2=3.5 $Y2=1.8
r107 14 47 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.335 $Y=4.265
+ $X2=3.335 $Y2=4.43
r108 13 16 26.9307 $w=3.3e-07 $l=2.33345e-07 $layer=POLY_cond $X=3.335 $Y=1.965
+ $X2=3.5 $Y2=1.8
r109 13 14 402.181 $w=3.3e-07 $l=2.3e-06 $layer=POLY_cond $X=3.335 $Y=1.965
+ $X2=3.335 $Y2=4.265
r110 4 53 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=4.275 $X2=3.835 $Y2=4.42
r111 4 50 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=4.275 $X2=3.835 $Y2=5.25
r112 3 39 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.96
+ $Y=3.175 $X2=2.085 $Y2=3.32
r113 2 37 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.96
+ $Y=2.125 $X2=2.085 $Y2=2.27
r114 1 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=0.705 $X2=2.085 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%VPWR 1 2 9 13 15 16 22 28 35 41
r67 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.605 $Y=4.58
+ $X2=0.605 $Y2=4.58
r68 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.605 $Y=3.56
+ $X2=0.605 $Y2=3.56
r69 16 41 0.0921373 $w=3.7e-07 $l=2.4e-07 $layer=MET1_cond $X=4.08 $Y=4.51
+ $X2=4.32 $Y2=4.51
r70 16 29 1.33407 $w=3.7e-07 $l=3.475e-06 $layer=MET1_cond $X=4.08 $Y=4.51
+ $X2=0.605 $Y2=4.51
r71 15 35 0.0921373 $w=3.7e-07 $l=2.4e-07 $layer=MET1_cond $X=4.08 $Y=3.63
+ $X2=4.32 $Y2=3.63
r72 15 23 1.33407 $w=3.7e-07 $l=3.475e-06 $layer=MET1_cond $X=4.08 $Y=3.63
+ $X2=0.605 $Y2=3.63
r73 11 28 15.5329 $w=2.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.295 $Y=4.58
+ $X2=0.605 $Y2=4.58
r74 11 13 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=0.295 $Y=4.695
+ $X2=0.295 $Y2=5.715
r75 7 22 15.5329 $w=2.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.295 $Y=3.56
+ $X2=0.605 $Y2=3.56
r76 7 9 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=0.295 $Y=3.445
+ $X2=0.295 $Y2=2.425
r77 2 13 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=5.505 $X2=0.295 $Y2=5.715
r78 1 9 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.215 $X2=0.295 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%X 1 2 7 8 9 10 11 12 20
r15 12 37 7.68008 $w=4.73e-07 $l=3.05e-07 $layer=LI1_cond $X=3.722 $Y=2.775
+ $X2=3.722 $Y2=3.08
r16 11 12 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.722 $Y=2.405
+ $X2=3.722 $Y2=2.775
r17 11 31 3.90299 $w=4.73e-07 $l=1.55e-07 $layer=LI1_cond $X=3.722 $Y=2.405
+ $X2=3.722 $Y2=2.25
r18 10 31 5.41383 $w=4.73e-07 $l=2.15e-07 $layer=LI1_cond $X=3.722 $Y=2.035
+ $X2=3.722 $Y2=2.25
r19 9 10 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.722 $Y=1.665
+ $X2=3.722 $Y2=2.035
r20 8 9 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.722 $Y=1.295
+ $X2=3.722 $Y2=1.665
r21 7 8 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.722 $Y=0.925
+ $X2=3.722 $Y2=1.295
r22 7 20 0.629515 $w=4.73e-07 $l=2.5e-08 $layer=LI1_cond $X=3.722 $Y=0.925
+ $X2=3.722 $Y2=0.9
r23 2 37 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=2.105 $X2=3.835 $Y2=3.08
r24 2 31 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=2.105 $X2=3.835 $Y2=2.25
r25 1 20 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=3.71
+ $Y=0.755 $X2=3.835 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%VGND 1 2 3 4 5 6 7 8 25 26 30 37 44 53
+ 64 65 75 83
r66 65 75 0.109413 $w=3.7e-07 $l=2.85e-07 $layer=MET1_cond $X=4.605 $Y=0.44
+ $X2=4.32 $Y2=0.44
r67 64 68 7.90628 $w=5.88e-07 $l=3.9e-07 $layer=LI1_cond $X=4.425 $Y=0.51
+ $X2=4.425 $Y2=0.9
r68 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.605 $Y=0.51
+ $X2=4.605 $Y2=0.51
r69 59 61 21.2861 $w=5.88e-07 $l=1.05e-06 $layer=LI1_cond $X=2.865 $Y=2.27
+ $X2=2.865 $Y2=3.32
r70 57 59 28.787 $w=5.88e-07 $l=1.42e-06 $layer=LI1_cond $X=2.865 $Y=0.85
+ $X2=2.865 $Y2=2.27
r71 53 57 6.89266 $w=5.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.865 $Y=0.51
+ $X2=2.865 $Y2=0.85
r72 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.045 $Y=0.51
+ $X2=3.045 $Y2=0.51
r73 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.005 $Y=7.63
+ $X2=3.005 $Y2=7.63
r74 47 49 16.218 $w=5.88e-07 $l=8e-07 $layer=LI1_cond $X=2.825 $Y=6.83 $X2=2.825
+ $Y2=7.63
r75 44 47 21.2861 $w=5.88e-07 $l=1.05e-06 $layer=LI1_cond $X=2.825 $Y=5.78
+ $X2=2.825 $Y2=6.83
r76 41 50 0.627685 $w=3.7e-07 $l=1.635e-06 $layer=MET1_cond $X=1.37 $Y=7.7
+ $X2=3.005 $Y2=7.7
r77 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.37 $Y=7.63
+ $X2=1.37 $Y2=7.63
r78 37 40 14.9003 $w=5.88e-07 $l=7.35e-07 $layer=LI1_cond $X=1.19 $Y=6.895
+ $X2=1.19 $Y2=7.63
r79 31 54 0.643042 $w=3.7e-07 $l=1.675e-06 $layer=MET1_cond $X=1.37 $Y=0.44
+ $X2=3.045 $Y2=0.44
r80 30 34 6.89266 $w=5.88e-07 $l=3.4e-07 $layer=LI1_cond $X=1.19 $Y=0.51
+ $X2=1.19 $Y2=0.85
r81 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.37 $Y=0.51
+ $X2=1.37 $Y2=0.51
r82 26 83 0.0921373 $w=3.7e-07 $l=2.4e-07 $layer=MET1_cond $X=4.08 $Y=7.7
+ $X2=4.32 $Y2=7.7
r83 26 50 0.412698 $w=3.7e-07 $l=1.075e-06 $layer=MET1_cond $X=4.08 $Y=7.7
+ $X2=3.005 $Y2=7.7
r84 25 75 0.0921373 $w=3.7e-07 $l=2.4e-07 $layer=MET1_cond $X=4.08 $Y=0.44
+ $X2=4.32 $Y2=0.44
r85 25 54 0.397342 $w=3.7e-07 $l=1.035e-06 $layer=MET1_cond $X=4.08 $Y=0.44
+ $X2=3.045 $Y2=0.44
r86 8 68 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.125
+ $Y=0.755 $X2=4.265 $Y2=0.9
r87 7 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.725
+ $Y=6.685 $X2=2.865 $Y2=6.83
r88 6 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.725
+ $Y=5.635 $X2=2.865 $Y2=5.78
r89 5 61 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.725
+ $Y=3.175 $X2=2.865 $Y2=3.32
r90 4 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.725
+ $Y=2.125 $X2=2.865 $Y2=2.27
r91 3 57 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.725
+ $Y=0.705 $X2=2.865 $Y2=0.85
r92 2 37 91 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=2 $X=0.935
+ $Y=6.685 $X2=1.075 $Y2=6.895
r93 1 34 91 $w=1.7e-07 $l=4.53156e-07 $layer=licon1_NDIFF $count=2 $X=0.935
+ $Y=1.035 $X2=1.305 $Y2=0.85
.ends

