* File: sky130_fd_sc_hvl__o21ai_1.pex.spice
* Created: Wed Sep  2 09:08:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__O21AI_1%VNB 5 7 11 25
r24 7 25 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0.058
r25 7 11 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0
r26 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r27 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__O21AI_1%VPB 4 6 14 21
r25 10 21 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=4.07
+ $X2=1.68 $Y2=4.013
r26 10 14 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=4.07
+ $X2=3.12 $Y2=4.07
r27 9 14 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=3.12 $Y2=4.07
r28 9 10 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r29 6 21 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=4.012
+ $X2=1.68 $Y2=4.013
r30 4 14 52 $w=1.7e-07 $l=3.16221e-06 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=3.12 $Y2=4.07
r31 4 9 52 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__O21AI_1%A1 3 7 9 10 15
r27 15 17 6.72742 $w=6.09e-07 $l=8.5e-08 $layer=POLY_cond $X=0.69 $Y=1.75
+ $X2=0.775 $Y2=1.75
r28 13 15 0.395731 $w=6.09e-07 $l=5e-09 $layer=POLY_cond $X=0.685 $Y=1.75
+ $X2=0.69 $Y2=1.75
r29 10 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=1.67 $X2=0.69 $Y2=1.67
r30 9 10 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.24 $Y=1.67 $X2=0.69
+ $Y2=1.67
r31 5 17 7.48396 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.775 $Y=2.085
+ $X2=0.775 $Y2=1.75
r32 5 7 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.775 $Y=2.085 $X2=0.775
+ $Y2=2.965
r33 1 13 7.48396 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.685 $Y=1.415
+ $X2=0.685 $Y2=1.75
r34 1 3 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.685 $Y=1.415 $X2=0.685
+ $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HVL__O21AI_1%A2 1 2 6 12
c27 6 0 8.58809e-20 $X=1.485 $Y=0.91
r28 9 12 142.853 $w=5e-07 $l=1.335e-06 $layer=POLY_cond $X=1.485 $Y=1.63
+ $X2=1.485 $Y2=2.965
r29 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.63 $X2=1.42 $Y2=1.63
r30 6 9 77.0442 $w=5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.485 $Y=0.91 $X2=1.485
+ $Y2=1.63
r31 2 10 11.7504 $w=2.53e-07 $l=2.6e-07 $layer=LI1_cond $X=1.68 $Y=1.632
+ $X2=1.42 $Y2=1.632
r32 1 10 9.94265 $w=2.53e-07 $l=2.2e-07 $layer=LI1_cond $X=1.2 $Y=1.632 $X2=1.42
+ $Y2=1.632
.ends

.subckt PM_SKY130_FD_SC_HVL__O21AI_1%B1 3 7 9 10 14
c29 10 0 8.58809e-20 $X=3.12 $Y=2.035
r30 14 17 19.0792 $w=6.6e-07 $l=1.95e-07 $layer=POLY_cond $X=2.345 $Y=1.89
+ $X2=2.345 $Y2=2.085
r31 14 16 41.7774 $w=6.6e-07 $l=4.75e-07 $layer=POLY_cond $X=2.345 $Y=1.89
+ $X2=2.345 $Y2=1.415
r32 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=1.89 $X2=2.49 $Y2=1.89
r33 9 10 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.962 $X2=3.12
+ $Y2=1.962
r34 9 15 5.48782 $w=3.13e-07 $l=1.5e-07 $layer=LI1_cond $X=2.64 $Y=1.962
+ $X2=2.49 $Y2=1.962
r35 7 17 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.265 $Y=2.965
+ $X2=2.265 $Y2=2.085
r36 3 16 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.265 $Y=0.91 $X2=2.265
+ $Y2=1.415
.ends

.subckt PM_SKY130_FD_SC_HVL__O21AI_1%VPWR 1 2 7 10 20 27
r25 24 27 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.335 $Y=3.63
+ $X2=3.055 $Y2=3.63
r26 23 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.055 $Y=3.59
+ $X2=3.055 $Y2=3.59
r27 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.335 $Y=3.59
+ $X2=2.335 $Y2=3.59
r28 20 23 15.4747 $w=9.48e-07 $l=1.205e-06 $layer=LI1_cond $X=2.695 $Y=2.385
+ $X2=2.695 $Y2=3.59
r29 14 17 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.205 $Y=3.63
+ $X2=0.925 $Y2=3.63
r30 13 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.925 $Y=3.59
+ $X2=0.925 $Y2=3.59
r31 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.205 $Y=3.59
+ $X2=0.205 $Y2=3.59
r32 10 13 16.0526 $w=9.48e-07 $l=1.25e-06 $layer=LI1_cond $X=0.565 $Y=2.34
+ $X2=0.565 $Y2=3.59
r33 7 24 0.251458 $w=3.7e-07 $l=6.55e-07 $layer=MET1_cond $X=1.68 $Y=3.63
+ $X2=2.335 $Y2=3.63
r34 7 17 0.289849 $w=3.7e-07 $l=7.55e-07 $layer=MET1_cond $X=1.68 $Y=3.63
+ $X2=0.925 $Y2=3.63
r35 2 23 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.515
+ $Y=2.215 $X2=2.655 $Y2=3.59
r36 2 20 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=2.515
+ $Y=2.215 $X2=2.655 $Y2=2.385
r37 1 13 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.24
+ $Y=2.215 $X2=0.385 $Y2=3.59
r38 1 10 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.24
+ $Y=2.215 $X2=0.385 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__O21AI_1%Y 1 2 9 10 13 15 16 17 18 38 40
r36 40 41 1.974 $w=5.78e-07 $l=7.5e-08 $layer=LI1_cond $X=1.855 $Y=2.035
+ $X2=1.855 $Y2=2.11
r37 18 35 11.2054 $w=4.73e-07 $l=4.45e-07 $layer=LI1_cond $X=1.802 $Y=3.145
+ $X2=1.802 $Y2=3.59
r38 17 18 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=1.802 $Y=2.775
+ $X2=1.802 $Y2=3.145
r39 16 17 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=1.802 $Y=2.405
+ $X2=1.802 $Y2=2.775
r40 16 27 1.63674 $w=4.73e-07 $l=6.5e-08 $layer=LI1_cond $X=1.802 $Y=2.405
+ $X2=1.802 $Y2=2.34
r41 15 40 0.10311 $w=5.78e-07 $l=5e-09 $layer=LI1_cond $X=1.855 $Y=2.03
+ $X2=1.855 $Y2=2.035
r42 15 38 8.47923 $w=5.78e-07 $l=9e-08 $layer=LI1_cond $X=1.855 $Y=2.03
+ $X2=1.855 $Y2=1.94
r43 15 27 5.66563 $w=4.73e-07 $l=2.25e-07 $layer=LI1_cond $X=1.802 $Y=2.115
+ $X2=1.802 $Y2=2.34
r44 15 41 0.125903 $w=4.73e-07 $l=5e-09 $layer=LI1_cond $X=1.802 $Y=2.115
+ $X2=1.802 $Y2=2.11
r45 11 13 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=2.655 $Y=1.455
+ $X2=2.655 $Y2=0.66
r46 9 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.49 $Y=1.54
+ $X2=2.655 $Y2=1.455
r47 9 10 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.49 $Y=1.54
+ $X2=2.145 $Y2=1.54
r48 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.06 $Y=1.625
+ $X2=2.145 $Y2=1.54
r49 7 38 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.06 $Y=1.625
+ $X2=2.06 $Y2=1.94
r50 2 35 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.735
+ $Y=2.215 $X2=1.875 $Y2=3.59
r51 2 27 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.735
+ $Y=2.215 $X2=1.875 $Y2=2.34
r52 1 13 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.515
+ $Y=0.535 $X2=2.655 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__O21AI_1%A_30_107# 1 2 9 11 12 15
r28 13 15 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.875 $Y=1.105
+ $X2=1.875 $Y2=0.66
r29 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.71 $Y=1.19
+ $X2=1.875 $Y2=1.105
r30 11 12 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=1.71 $Y=1.19
+ $X2=0.46 $Y2=1.19
r31 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.295 $Y=1.105
+ $X2=0.46 $Y2=1.19
r32 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.295 $Y=1.105
+ $X2=0.295 $Y2=0.66
r33 2 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.735
+ $Y=0.535 $X2=1.875 $Y2=0.66
r34 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.535 $X2=0.295 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__O21AI_1%VGND 1 4 7
r18 8 11 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.725 $Y=0.44
+ $X2=1.445 $Y2=0.44
r19 7 13 3.70112 $w=8.88e-07 $l=2.7e-07 $layer=LI1_cond $X=1.085 $Y=0.48
+ $X2=1.085 $Y2=0.75
r20 7 11 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.445 $Y=0.48
+ $X2=1.445 $Y2=0.48
r21 7 8 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.725 $Y=0.48
+ $X2=0.725 $Y2=0.48
r22 4 11 0.0902178 $w=3.7e-07 $l=2.35e-07 $layer=MET1_cond $X=1.68 $Y=0.44
+ $X2=1.445 $Y2=0.44
r23 1 13 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=0.935
+ $Y=0.535 $X2=1.075 $Y2=0.75
.ends

