* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
*.PININFO A1:I A2:I B1:I B2:I VGND:I VNB:I VPB:I VPWR:I X:O
MMPA0 VPWR A1 VPB phv m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MMPA1 sndA1 A2 VPB phv m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMPB0 VPWR B1 VPB phv m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MMPB1 sndB1 B2 VPB phv m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIPX X y VPB phv m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MMNA0 pndA A1 VNB nhv m=1 w=0.75 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMNA1 pndA A2 VNB nhv m=1 w=0.75 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMNB0 y B1 VNB nhv m=1 w=0.75 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MMNB1 y B2 VNB nhv m=1 w=0.75 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MMINX X y VNB nhv m=1 w=0.75 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_hvl__o22a_1
