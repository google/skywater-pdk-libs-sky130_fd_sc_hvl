* File: sky130_fd_sc_hvl__o22ai_1.pxi.spice
* Created: Fri Aug 28 09:38:55 2020
* 
x_PM_SKY130_FD_SC_HVL__O22AI_1%VNB N_VNB_M1006_b VNB N_VNB_c_7_p VNB
+ PM_SKY130_FD_SC_HVL__O22AI_1%VNB
x_PM_SKY130_FD_SC_HVL__O22AI_1%VPB N_VPB_M1002_b VPB N_VPB_c_31_p VPB
+ PM_SKY130_FD_SC_HVL__O22AI_1%VPB
x_PM_SKY130_FD_SC_HVL__O22AI_1%B1 N_B1_c_60_n N_B1_M1006_g N_B1_M1002_g B1
+ N_B1_c_61_n N_B1_c_62_n PM_SKY130_FD_SC_HVL__O22AI_1%B1
x_PM_SKY130_FD_SC_HVL__O22AI_1%B2 B2 N_B2_M1001_g N_B2_c_90_n N_B2_M1003_g
+ PM_SKY130_FD_SC_HVL__O22AI_1%B2
x_PM_SKY130_FD_SC_HVL__O22AI_1%A2 N_A2_M1000_g N_A2_M1004_g A2 N_A2_c_123_n
+ N_A2_c_126_n PM_SKY130_FD_SC_HVL__O22AI_1%A2
x_PM_SKY130_FD_SC_HVL__O22AI_1%A1 N_A1_M1005_g N_A1_M1007_g A1 A1 N_A1_c_157_n
+ PM_SKY130_FD_SC_HVL__O22AI_1%A1
x_PM_SKY130_FD_SC_HVL__O22AI_1%VPWR N_VPWR_M1002_s N_VPWR_M1005_d VPWR
+ N_VPWR_c_180_n N_VPWR_c_183_n N_VPWR_c_186_n PM_SKY130_FD_SC_HVL__O22AI_1%VPWR
x_PM_SKY130_FD_SC_HVL__O22AI_1%Y N_Y_M1006_d N_Y_M1003_d N_Y_c_222_n N_Y_c_217_n
+ N_Y_c_226_n N_Y_c_218_n N_Y_c_216_n Y Y Y Y N_Y_c_221_n Y
+ PM_SKY130_FD_SC_HVL__O22AI_1%Y
x_PM_SKY130_FD_SC_HVL__O22AI_1%A_36_113# N_A_36_113#_M1006_s N_A_36_113#_M1001_d
+ N_A_36_113#_M1007_d N_A_36_113#_c_262_n N_A_36_113#_c_263_n
+ N_A_36_113#_c_265_n N_A_36_113#_c_267_n N_A_36_113#_c_268_n
+ N_A_36_113#_c_269_n N_A_36_113#_c_270_n PM_SKY130_FD_SC_HVL__O22AI_1%A_36_113#
x_PM_SKY130_FD_SC_HVL__O22AI_1%VGND N_VGND_M1000_d VGND N_VGND_c_305_n
+ N_VGND_c_307_n PM_SKY130_FD_SC_HVL__O22AI_1%VGND
cc_1 N_VNB_M1006_b N_B1_c_60_n 0.0416236f $X=-0.33 $Y=-0.265 $X2=0.715 $Y2=1.425
cc_2 N_VNB_M1006_b N_B1_c_61_n 0.0153315f $X=-0.33 $Y=-0.265 $X2=0.385 $Y2=1.7
cc_3 N_VNB_M1006_b N_B1_c_62_n 0.0733945f $X=-0.33 $Y=-0.265 $X2=0.785 $Y2=1.675
cc_4 N_VNB_M1006_b N_B2_M1001_g 0.0771667f $X=-0.33 $Y=-0.265 $X2=0.785
+ $Y2=1.925
cc_5 N_VNB_M1006_b N_B2_c_90_n 0.00428125f $X=-0.33 $Y=-0.265 $X2=0.155 $Y2=1.58
cc_6 N_VNB_M1006_b N_A2_M1000_g 0.0556164f $X=-0.33 $Y=-0.265 $X2=0.715 $Y2=0.94
cc_7 N_VNB_c_7_p N_A2_M1000_g 5.66372e-19 $X=0.24 $Y=0 $X2=0.715 $Y2=0.94
cc_8 N_VNB_M1006_b A2 0.00199371f $X=-0.33 $Y=-0.265 $X2=0.155 $Y2=1.58
cc_9 N_VNB_M1006_b N_A2_c_123_n 0.0287598f $X=-0.33 $Y=-0.265 $X2=0.385 $Y2=1.7
cc_10 N_VNB_M1006_b N_A1_M1007_g 0.0465714f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_11 N_VNB_c_7_p N_A1_M1007_g 7.01222e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_12 N_VNB_M1006_b A1 0.00778592f $X=-0.33 $Y=-0.265 $X2=0.385 $Y2=1.675
cc_13 N_VNB_M1006_b N_A1_c_157_n 0.0542819f $X=-0.33 $Y=-0.265 $X2=0.715
+ $Y2=1.675
cc_14 N_VNB_M1006_b N_Y_c_216_n 0.0027787f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_15 N_VNB_M1006_b N_A_36_113#_c_262_n 0.0329145f $X=-0.33 $Y=-0.265 $X2=0.385
+ $Y2=1.7
cc_16 N_VNB_M1006_b N_A_36_113#_c_263_n 0.124375f $X=-0.33 $Y=-0.265 $X2=0.715
+ $Y2=1.675
cc_17 N_VNB_c_7_p N_A_36_113#_c_263_n 0.00498793f $X=0.24 $Y=0 $X2=0.715
+ $Y2=1.675
cc_18 N_VNB_M1006_b N_A_36_113#_c_265_n 0.0264953f $X=-0.33 $Y=-0.265 $X2=0.785
+ $Y2=1.675
cc_19 N_VNB_c_7_p N_A_36_113#_c_265_n 0.00109438f $X=0.24 $Y=0 $X2=0.785
+ $Y2=1.675
cc_20 N_VNB_M1006_b N_A_36_113#_c_267_n 0.00561831f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_21 N_VNB_M1006_b N_A_36_113#_c_268_n 0.0181814f $X=-0.33 $Y=-0.265 $X2=0.385
+ $Y2=1.7
cc_22 N_VNB_M1006_b N_A_36_113#_c_269_n 0.0043722f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_23 N_VNB_M1006_b N_A_36_113#_c_270_n 0.0159283f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_24 N_VNB_c_7_p N_A_36_113#_c_270_n 5.57033e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_25 N_VNB_M1006_b N_VGND_c_305_n 0.0545569f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_26 N_VNB_c_7_p N_VGND_c_305_n 0.0031162f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_27 N_VNB_M1006_b N_VGND_c_307_n 0.0755567f $X=-0.33 $Y=-0.265 $X2=0.385
+ $Y2=1.7
cc_28 N_VNB_c_7_p N_VGND_c_307_n 0.410192f $X=0.24 $Y=0 $X2=0.385 $Y2=1.7
cc_29 N_VPB_M1002_b N_B1_M1002_g 0.0604871f $X=-0.33 $Y=1.885 $X2=0.785
+ $Y2=2.965
cc_30 VPB N_B1_M1002_g 0.00970178f $X=0 $Y=3.955 $X2=0.785 $Y2=2.965
cc_31 N_VPB_c_31_p N_B1_M1002_g 0.0137101f $X=3.6 $Y=4.07 $X2=0.785 $Y2=2.965
cc_32 N_VPB_M1002_b N_B1_c_62_n 0.0161206f $X=-0.33 $Y=1.885 $X2=0.785 $Y2=1.675
cc_33 N_VPB_M1002_b N_B2_M1001_g 0.0505536f $X=-0.33 $Y=1.885 $X2=0.785
+ $Y2=1.925
cc_34 VPB N_B2_M1001_g 0.00970178f $X=0 $Y=3.955 $X2=0.785 $Y2=1.925
cc_35 N_VPB_c_31_p N_B2_M1001_g 0.018494f $X=3.6 $Y=4.07 $X2=0.785 $Y2=1.925
cc_36 N_VPB_M1002_b A2 0.00302372f $X=-0.33 $Y=1.885 $X2=0.155 $Y2=1.58
cc_37 N_VPB_M1002_b N_A2_c_123_n 0.0235459f $X=-0.33 $Y=1.885 $X2=0.385 $Y2=1.7
cc_38 N_VPB_M1002_b N_A2_c_126_n 0.0336119f $X=-0.33 $Y=1.885 $X2=0.715
+ $Y2=1.675
cc_39 VPB N_A2_c_126_n 0.00970178f $X=0 $Y=3.955 $X2=0.715 $Y2=1.675
cc_40 N_VPB_c_31_p N_A2_c_126_n 0.0161677f $X=3.6 $Y=4.07 $X2=0.715 $Y2=1.675
cc_41 N_VPB_M1002_b N_A1_M1005_g 0.0411028f $X=-0.33 $Y=1.885 $X2=0.715 $Y2=0.94
cc_42 VPB N_A1_M1005_g 0.00970178f $X=0 $Y=3.955 $X2=0.715 $Y2=0.94
cc_43 N_VPB_c_31_p N_A1_M1005_g 0.0137101f $X=3.6 $Y=4.07 $X2=0.715 $Y2=0.94
cc_44 N_VPB_M1002_b A1 0.0173206f $X=-0.33 $Y=1.885 $X2=0.385 $Y2=1.675
cc_45 N_VPB_M1002_b N_A1_c_157_n 0.0244107f $X=-0.33 $Y=1.885 $X2=0.715
+ $Y2=1.675
cc_46 N_VPB_M1002_b N_VPWR_c_180_n 0.0660851f $X=-0.33 $Y=1.885 $X2=0.385
+ $Y2=1.675
cc_47 VPB N_VPWR_c_180_n 0.00487913f $X=0 $Y=3.955 $X2=0.385 $Y2=1.675
cc_48 N_VPB_c_31_p N_VPWR_c_180_n 0.063841f $X=3.6 $Y=4.07 $X2=0.385 $Y2=1.675
cc_49 N_VPB_M1002_b N_VPWR_c_183_n 0.0543016f $X=-0.33 $Y=1.885 $X2=0.385
+ $Y2=1.7
cc_50 VPB N_VPWR_c_183_n 0.00538585f $X=0 $Y=3.955 $X2=0.385 $Y2=1.7
cc_51 N_VPB_c_31_p N_VPWR_c_183_n 0.0659756f $X=3.6 $Y=4.07 $X2=0.385 $Y2=1.7
cc_52 N_VPB_M1002_b N_VPWR_c_186_n 0.0499498f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_186_n 0.407263f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_54 N_VPB_c_31_p N_VPWR_c_186_n 0.0175634f $X=3.6 $Y=4.07 $X2=0 $Y2=0
cc_55 N_VPB_M1002_b N_Y_c_217_n 0.00415002f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_56 N_VPB_M1002_b N_Y_c_218_n 0.00151825f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_57 VPB N_Y_c_218_n 5.14916e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_58 N_VPB_c_31_p N_Y_c_218_n 0.00887752f $X=3.6 $Y=4.07 $X2=0 $Y2=0
cc_59 N_VPB_M1002_b N_Y_c_221_n 0.00887177f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_60 N_B1_c_60_n N_B2_M1001_g 0.0169167f $X=0.715 $Y=1.425 $X2=0 $Y2=0
cc_61 N_B1_c_62_n N_B2_M1001_g 0.163505f $X=0.785 $Y=1.675 $X2=0 $Y2=0
cc_62 N_B1_c_62_n N_B2_c_90_n 0.00181283f $X=0.785 $Y=1.675 $X2=0 $Y2=0
cc_63 N_B1_M1002_g N_VPWR_c_180_n 0.10148f $X=0.785 $Y=2.965 $X2=0.24 $Y2=0
cc_64 N_B1_c_61_n N_VPWR_c_180_n 0.0168044f $X=0.385 $Y=1.7 $X2=0.24 $Y2=0
cc_65 N_B1_c_62_n N_VPWR_c_180_n 0.00757493f $X=0.785 $Y=1.675 $X2=0.24 $Y2=0
cc_66 N_B1_M1002_g N_VPWR_c_186_n 0.0023336f $X=0.785 $Y=2.965 $X2=0 $Y2=0
cc_67 N_B1_c_60_n N_Y_c_222_n 0.00471324f $X=0.715 $Y=1.425 $X2=0 $Y2=0
cc_68 N_B1_c_61_n N_Y_c_222_n 0.0224481f $X=0.385 $Y=1.7 $X2=0 $Y2=0
cc_69 N_B1_c_62_n N_Y_c_222_n 0.02559f $X=0.785 $Y=1.675 $X2=0 $Y2=0
cc_70 N_B1_M1002_g N_Y_c_217_n 0.00861473f $X=0.785 $Y=2.965 $X2=0 $Y2=0
cc_71 N_B1_M1002_g N_Y_c_226_n 0.0130082f $X=0.785 $Y=2.965 $X2=0.24 $Y2=0
cc_72 N_B1_c_60_n N_Y_c_216_n 0.0334847f $X=0.715 $Y=1.425 $X2=3.6 $Y2=0
cc_73 N_B1_c_62_n N_Y_c_216_n 0.00263447f $X=0.785 $Y=1.675 $X2=3.6 $Y2=0
cc_74 N_B1_M1002_g Y 4.18849e-19 $X=0.785 $Y=2.965 $X2=0 $Y2=0
cc_75 N_B1_M1002_g N_Y_c_221_n 8.33916e-19 $X=0.785 $Y=2.965 $X2=0 $Y2=0
cc_76 N_B1_c_60_n N_A_36_113#_c_262_n 0.0246583f $X=0.715 $Y=1.425 $X2=0 $Y2=0
cc_77 N_B1_c_61_n N_A_36_113#_c_262_n 0.0265457f $X=0.385 $Y=1.7 $X2=0 $Y2=0
cc_78 N_B1_c_62_n N_A_36_113#_c_262_n 0.00762292f $X=0.785 $Y=1.675 $X2=0 $Y2=0
cc_79 N_B1_c_60_n N_A_36_113#_c_263_n 0.0156294f $X=0.715 $Y=1.425 $X2=0 $Y2=0
cc_80 N_B1_c_60_n N_A_36_113#_c_265_n 4.26793e-19 $X=0.715 $Y=1.425 $X2=0 $Y2=0
cc_81 N_B1_c_60_n N_VGND_c_307_n 0.0173641f $X=0.715 $Y=1.425 $X2=0.24 $Y2=0
cc_82 N_B2_M1001_g N_A2_M1000_g 0.0500596f $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_83 N_B2_M1001_g A2 7.40318e-19 $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_84 N_B2_c_90_n N_A2_c_123_n 6.70176e-19 $X=1.43 $Y=1.645 $X2=0.24 $Y2=0
cc_85 N_B2_M1001_g N_A2_c_126_n 0.0358171f $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_86 N_B2_M1001_g N_VPWR_c_180_n 0.0530067f $X=1.495 $Y=0.94 $X2=0.24 $Y2=0
cc_87 N_B2_M1001_g N_VPWR_c_183_n 6.30873e-19 $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_88 N_B2_M1001_g N_VPWR_c_186_n 0.0196953f $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_89 N_B2_M1001_g N_Y_c_222_n 0.00223219f $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_90 N_B2_c_90_n N_Y_c_222_n 0.0160571f $X=1.43 $Y=1.645 $X2=0 $Y2=0
cc_91 N_B2_M1001_g N_Y_c_217_n 0.0192329f $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_92 N_B2_c_90_n N_Y_c_217_n 0.0302118f $X=1.43 $Y=1.645 $X2=0 $Y2=0
cc_93 N_B2_M1001_g N_Y_c_218_n 0.00517036f $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_94 N_B2_M1001_g N_Y_c_216_n 0.0207508f $X=1.495 $Y=0.94 $X2=3.6 $Y2=0
cc_95 N_B2_c_90_n N_Y_c_216_n 0.0149624f $X=1.43 $Y=1.645 $X2=3.6 $Y2=0
cc_96 N_B2_M1001_g Y 0.0262987f $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_97 N_B2_M1001_g Y 0.0160195f $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_98 N_B2_M1001_g N_Y_c_221_n 0.0291654f $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_99 N_B2_c_90_n N_Y_c_221_n 0.00517569f $X=1.43 $Y=1.645 $X2=0 $Y2=0
cc_100 N_B2_M1001_g N_A_36_113#_c_263_n 0.0198402f $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_101 N_B2_M1001_g N_A_36_113#_c_267_n 0.0067609f $X=1.495 $Y=0.94 $X2=0 $Y2=0
cc_102 N_B2_M1001_g N_A_36_113#_c_269_n 0.00357092f $X=1.495 $Y=0.94 $X2=1.92
+ $Y2=0
cc_103 N_B2_c_90_n N_A_36_113#_c_269_n 0.00674588f $X=1.43 $Y=1.645 $X2=1.92
+ $Y2=0
cc_104 N_B2_M1001_g N_VGND_c_307_n 0.0298849f $X=1.495 $Y=0.94 $X2=0.24 $Y2=0
cc_105 N_A2_c_126_n N_A1_M1005_g 0.0759736f $X=2.312 $Y=2.105 $X2=0 $Y2=0
cc_106 N_A2_M1000_g N_A1_M1007_g 0.0232259f $X=2.275 $Y=0.94 $X2=0 $Y2=0
cc_107 A2 A1 0.0204076f $X=2.555 $Y=1.95 $X2=0.24 $Y2=0
cc_108 N_A2_c_123_n A1 2.28443e-19 $X=2.415 $Y=1.89 $X2=0.24 $Y2=0
cc_109 N_A2_M1000_g N_A1_c_157_n 0.00729262f $X=2.275 $Y=0.94 $X2=0 $Y2=0
cc_110 A2 N_A1_c_157_n 0.00296132f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_111 N_A2_c_123_n N_A1_c_157_n 0.0759736f $X=2.415 $Y=1.89 $X2=0 $Y2=0
cc_112 A2 N_VPWR_c_183_n 0.0326434f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_113 N_A2_c_126_n N_VPWR_c_183_n 0.0757857f $X=2.312 $Y=2.105 $X2=0 $Y2=0
cc_114 N_A2_c_126_n N_VPWR_c_186_n 0.0125055f $X=2.312 $Y=2.105 $X2=0 $Y2=0
cc_115 N_A2_c_126_n N_Y_c_218_n 0.00135461f $X=2.312 $Y=2.105 $X2=0 $Y2=0
cc_116 A2 N_Y_c_221_n 0.00778746f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_117 N_A2_c_123_n N_Y_c_221_n 0.00258709f $X=2.415 $Y=1.89 $X2=0 $Y2=0
cc_118 N_A2_c_126_n N_Y_c_221_n 0.00255801f $X=2.312 $Y=2.105 $X2=0 $Y2=0
cc_119 N_A2_M1000_g N_A_36_113#_c_267_n 0.00503751f $X=2.275 $Y=0.94 $X2=0 $Y2=0
cc_120 N_A2_M1000_g N_A_36_113#_c_268_n 0.0209272f $X=2.275 $Y=0.94 $X2=0 $Y2=0
cc_121 A2 N_A_36_113#_c_268_n 0.0355461f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_122 N_A2_c_123_n N_A_36_113#_c_268_n 0.0170019f $X=2.415 $Y=1.89 $X2=0 $Y2=0
cc_123 N_A2_M1000_g N_VGND_c_305_n 0.0507364f $X=2.275 $Y=0.94 $X2=0 $Y2=0
cc_124 N_A2_c_123_n N_VGND_c_305_n 2.76268e-19 $X=2.415 $Y=1.89 $X2=0 $Y2=0
cc_125 N_A2_M1000_g N_VGND_c_307_n 0.00784072f $X=2.275 $Y=0.94 $X2=0.24 $Y2=0
cc_126 N_A1_M1005_g N_VPWR_c_183_n 0.0959711f $X=3.06 $Y=2.965 $X2=0 $Y2=0
cc_127 A1 N_VPWR_c_183_n 0.0459066f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_128 N_A1_c_157_n N_VPWR_c_183_n 5.06543e-19 $X=3.21 $Y=1.89 $X2=0 $Y2=0
cc_129 N_A1_M1005_g N_VPWR_c_186_n 0.00233214f $X=3.06 $Y=2.965 $X2=0 $Y2=0
cc_130 A1 N_A_36_113#_c_268_n 0.0494519f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_131 N_A1_c_157_n N_A_36_113#_c_268_n 0.0382053f $X=3.21 $Y=1.89 $X2=0 $Y2=0
cc_132 N_A1_M1007_g N_A_36_113#_c_270_n 0.0106824f $X=3.155 $Y=0.94 $X2=1.92
+ $Y2=0.058
cc_133 N_A1_M1007_g N_VGND_c_305_n 0.0586819f $X=3.155 $Y=0.94 $X2=0 $Y2=0
cc_134 N_A1_c_157_n N_VGND_c_305_n 0.0024204f $X=3.21 $Y=1.89 $X2=0 $Y2=0
cc_135 N_A1_M1007_g N_VGND_c_307_n 0.0104481f $X=3.155 $Y=0.94 $X2=0.24 $Y2=0
cc_136 N_VPWR_c_180_n A_207_443# 0.00109099f $X=0.395 $Y=2.365 $X2=0 $Y2=3.985
cc_137 N_VPWR_c_186_n N_Y_M1003_d 0.00335282f $X=3.5 $Y=3.59 $X2=0 $Y2=0
cc_138 N_VPWR_c_180_n N_Y_c_217_n 0.0283781f $X=0.395 $Y=2.365 $X2=0.24 $Y2=4.07
cc_139 N_VPWR_c_180_n N_Y_c_226_n 0.0136575f $X=0.395 $Y=2.365 $X2=0.24 $Y2=4.07
cc_140 N_VPWR_c_180_n N_Y_c_218_n 0.010914f $X=0.395 $Y=2.365 $X2=3.6 $Y2=4.07
cc_141 N_VPWR_c_183_n N_Y_c_218_n 0.0405196f $X=3.45 $Y=2.385 $X2=3.6 $Y2=4.07
cc_142 N_VPWR_c_186_n N_Y_c_218_n 0.0276416f $X=3.5 $Y=3.59 $X2=3.6 $Y2=4.07
cc_143 N_VPWR_c_180_n Y 0.0646602f $X=0.395 $Y=2.365 $X2=1.92 $Y2=4.013
cc_144 N_VPWR_c_186_n Y 0.0179532f $X=3.5 $Y=3.59 $X2=1.92 $Y2=4.07
cc_145 N_VPWR_c_180_n N_Y_c_221_n 0.0122206f $X=0.395 $Y=2.365 $X2=0 $Y2=0
cc_146 N_VPWR_c_183_n A_520_443# 0.00109099f $X=3.45 $Y=2.385 $X2=0 $Y2=3.985
cc_147 N_VPWR_c_183_n N_A_36_113#_c_268_n 0.00546208f $X=3.45 $Y=2.385 $X2=1.92
+ $Y2=4.013
cc_148 N_Y_c_216_n N_A_36_113#_c_262_n 0.0429133f $X=1.105 $Y=0.7 $X2=0 $Y2=0
cc_149 N_Y_c_216_n N_A_36_113#_c_263_n 0.0332907f $X=1.105 $Y=0.7 $X2=0 $Y2=0
cc_150 N_Y_c_216_n N_A_36_113#_c_267_n 0.0124065f $X=1.105 $Y=0.7 $X2=0 $Y2=0
cc_151 N_Y_c_221_n N_A_36_113#_c_268_n 0.00270146f $X=1.785 $Y=2.435 $X2=0 $Y2=0
cc_152 N_Y_c_221_n N_A_36_113#_c_269_n 0.007017f $X=1.785 $Y=2.435 $X2=1.92
+ $Y2=0
cc_153 N_Y_c_216_n N_VGND_c_307_n 0.0369324f $X=1.105 $Y=0.7 $X2=0.24 $Y2=0
cc_154 N_A_36_113#_c_263_n N_VGND_c_305_n 0.00489946f $X=1.8 $Y=0.35 $X2=0 $Y2=0
cc_155 N_A_36_113#_c_267_n N_VGND_c_305_n 0.0371633f $X=1.885 $Y=0.69 $X2=0
+ $Y2=0
cc_156 N_A_36_113#_c_268_n N_VGND_c_305_n 0.077064f $X=3.42 $Y=1.54 $X2=0 $Y2=0
cc_157 N_A_36_113#_c_270_n N_VGND_c_305_n 0.0330149f $X=3.545 $Y=0.69 $X2=0
+ $Y2=0
cc_158 N_A_36_113#_M1001_d N_VGND_c_307_n 0.00442064f $X=1.745 $Y=0.565 $X2=0.24
+ $Y2=0
cc_159 N_A_36_113#_M1007_d N_VGND_c_307_n 0.00141794f $X=3.405 $Y=0.565 $X2=0.24
+ $Y2=0
cc_160 N_A_36_113#_c_262_n N_VGND_c_307_n 0.0359456f $X=0.325 $Y=0.69 $X2=0.24
+ $Y2=0
cc_161 N_A_36_113#_c_263_n N_VGND_c_307_n 0.0619502f $X=1.8 $Y=0.35 $X2=0.24
+ $Y2=0
cc_162 N_A_36_113#_c_265_n N_VGND_c_307_n 0.011429f $X=0.49 $Y=0.35 $X2=0.24
+ $Y2=0
cc_163 N_A_36_113#_c_267_n N_VGND_c_307_n 0.0215781f $X=1.885 $Y=0.69 $X2=0.24
+ $Y2=0
cc_164 N_A_36_113#_c_270_n N_VGND_c_307_n 0.0248336f $X=3.545 $Y=0.69 $X2=0.24
+ $Y2=0
