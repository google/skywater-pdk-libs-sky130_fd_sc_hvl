* File: sky130_fd_sc_hvl__dfsbp_1.spice
* Created: Wed Sep  2 09:05:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__dfsbp_1.pex.spice"
.subckt sky130_fd_sc_hvl__dfsbp_1  VNB VPB CLK D SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1023 N_VGND_M1023_d N_CLK_M1023_g N_A_30_112#_M1023_s N_VNB_M1023_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1005 N_A_339_112#_M1005_d N_A_30_112#_M1005_g N_VGND_M1023_d N_VNB_M1023_b NHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1001 N_A_605_109#_M1001_d N_D_M1001_g N_VGND_M1001_s N_VNB_M1023_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1014 N_A_761_109#_M1014_d N_A_30_112#_M1014_g N_A_605_109#_M1001_d
+ N_VNB_M1023_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0
+ M=1 R=0.84 SA=250001 SB=250002 A=0.21 P=1.84 MULT=1
MM1007 A_917_109# N_A_339_112#_M1007_g N_A_761_109#_M1014_d N_VNB_M1023_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1008 N_VGND_M1008_d N_A_959_83#_M1008_g A_917_109# N_VNB_M1023_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1025 A_1325_107# N_A_761_109#_M1025_g N_A_959_83#_M1025_s N_VNB_M1023_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1027 N_VGND_M1027_d N_SET_B_M1027_g A_1325_107# N_VNB_M1023_b NHV L=0.5 W=0.42
+ AD=0.0879308 AS=0.0441 PD=0.807692 PS=0.63 NRD=25.7754 NRS=13.566 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1029 N_A_1642_107#_M1029_d N_A_761_109#_M1029_g N_VGND_M1027_d N_VNB_M1023_b
+ NHV L=0.5 W=0.75 AD=0.19875 AS=0.157019 PD=2.03 PS=1.44231 NRD=0 NRS=0 M=1
+ R=1.5 SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1028 N_A_1874_543#_M1028_d N_A_30_112#_M1028_g N_A_1755_153#_M1028_s
+ N_VNB_M1023_b NHV L=0.5 W=0.42 AD=0.145097 AS=0.1197 PD=1.04821 PS=1.41
+ NRD=78.831 NRS=0 M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1010 N_A_1642_107#_M1010_d N_A_339_112#_M1010_g N_A_1874_543#_M1028_d
+ N_VNB_M1023_b NHV L=0.5 W=0.75 AD=0.375 AS=0.259103 PD=2.5 PS=1.87179
+ NRD=13.6686 NRS=44.1408 M=1 R=1.5 SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1019 A_2427_107# N_A_2156_417#_M1019_g N_A_1755_153#_M1019_s N_VNB_M1023_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1020 N_VGND_M1020_d N_SET_B_M1020_g A_2427_107# N_VNB_M1023_b NHV L=0.5 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250001
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1003 N_VGND_M1003_d N_A_1874_543#_M1003_g N_A_2156_417#_M1003_s N_VNB_M1023_b
+ NHV L=0.5 W=0.42 AD=0.0879308 AS=0.1197 PD=0.807692 PS=1.41 NRD=41.895 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1016 N_Q_N_M1016_d N_A_1874_543#_M1016_g N_VGND_M1003_d N_VNB_M1023_b NHV
+ L=0.5 W=0.75 AD=0.21375 AS=0.157019 PD=2.07 PS=1.44231 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1013 N_VGND_M1013_d N_A_1874_543#_M1013_g N_A_3129_479#_M1013_s N_VNB_M1023_b
+ NHV L=0.5 W=0.42 AD=0.0879308 AS=0.1197 PD=0.807692 PS=1.41 NRD=25.7754 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1002 N_Q_M1002_d N_A_3129_479#_M1002_g N_VGND_M1013_d N_VNB_M1023_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.157019 PD=2.07 PS=1.44231 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1017 N_VPWR_M1017_d N_CLK_M1017_g N_A_30_112#_M1017_s N_VPB_M1017_b PHV L=0.5
+ W=0.75 AD=0.105 AS=0.21375 PD=1.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1030 N_A_339_112#_M1030_d N_A_30_112#_M1030_g N_VPWR_M1017_d N_VPB_M1017_b PHV
+ L=0.5 W=0.75 AD=0.21375 AS=0.105 PD=2.07 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1022 N_A_605_109#_M1022_d N_D_M1022_g N_VPWR_M1022_s N_VPB_M1017_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1575 PD=0.7 PS=1.59 NRD=0 NRS=40.9122 M=1 R=0.84
+ SA=250000 SB=250009 A=0.21 P=1.84 MULT=1
MM1012 N_A_761_109#_M1012_d N_A_339_112#_M1012_g N_A_605_109#_M1022_d
+ N_VPB_M1017_b PHV L=0.5 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0
+ M=1 R=0.84 SA=250001 SB=250008 A=0.21 P=1.84 MULT=1
MM1031 A_976_543# N_A_30_112#_M1031_g N_A_761_109#_M1012_d N_VPB_M1017_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250002 SB=250007 A=0.21 P=1.84 MULT=1
MM1009 N_VPWR_M1009_d N_A_959_83#_M1009_g A_976_543# N_VPB_M1017_b PHV L=0.5
+ W=0.42 AD=0.1323 AS=0.0441 PD=1.05 PS=0.63 NRD=52.2958 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250007 A=0.21 P=1.84 MULT=1
MM1006 N_A_959_83#_M1006_d N_A_761_109#_M1006_g N_VPWR_M1009_d N_VPB_M1017_b PHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.1323 PD=0.7 PS=1.05 NRD=0 NRS=106.864 M=1 R=0.84
+ SA=250004 SB=250005 A=0.21 P=1.84 MULT=1
MM1032 N_VPWR_M1032_d N_SET_B_M1032_g N_A_959_83#_M1006_d N_VPB_M1017_b PHV
+ L=0.5 W=0.42 AD=0.124876 AS=0.0588 PD=0.981972 PS=0.7 NRD=172.798 NRS=0 M=1
+ R=0.84 SA=250004 SB=250005 A=0.21 P=1.84 MULT=1
MM1033 A_1732_543# N_A_761_109#_M1033_g N_VPWR_M1032_d N_VPB_M1017_b PHV L=0.5
+ W=1 AD=0.105 AS=0.297324 PD=1.21 PS=2.33803 NRD=9.5309 NRS=0 M=1 R=2 SA=250002
+ SB=250002 A=0.5 P=3 MULT=1
MM1000 N_A_1874_543#_M1000_d N_A_30_112#_M1000_g A_1732_543# N_VPB_M1017_b PHV
+ L=0.5 W=1 AD=0.233239 AS=0.105 PD=1.96479 PS=1.21 NRD=0 NRS=9.5309 M=1 R=2
+ SA=250003 SB=250001 A=0.5 P=3 MULT=1
MM1021 A_2053_543# N_A_339_112#_M1021_g N_A_1874_543#_M1000_d N_VPB_M1017_b PHV
+ L=0.5 W=0.42 AD=0.10815 AS=0.0979606 PD=0.935 PS=0.825211 NRD=92.0811
+ NRS=52.2958 M=1 R=0.84 SA=250007 SB=250002 A=0.21 P=1.84 MULT=1
MM1011 N_VPWR_M1011_d N_A_2156_417#_M1011_g A_2053_543# N_VPB_M1017_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.10815 PD=0.7 PS=0.935 NRD=0 NRS=92.0811 M=1 R=0.84
+ SA=250008 SB=250001 A=0.21 P=1.84 MULT=1
MM1004 N_A_1874_543#_M1004_d N_SET_B_M1004_g N_VPWR_M1011_d N_VPB_M1017_b PHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250009 SB=250000 A=0.21 P=1.84 MULT=1
MM1026 N_VPWR_M1026_d N_A_1874_543#_M1026_g N_A_2156_417#_M1026_s N_VPB_M1017_b
+ PHV L=0.5 W=0.42 AD=0.103622 AS=0.1197 PD=0.829062 PS=1.41 NRD=52.2958 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1018 N_Q_N_M1018_d N_A_1874_543#_M1018_g N_VPWR_M1026_d N_VPB_M1017_b PHV
+ L=0.5 W=1.5 AD=0.4275 AS=0.370078 PD=3.57 PS=2.96094 NRD=0 NRS=0 M=1 R=3
+ SA=250000 SB=250000 A=0.75 P=4 MULT=1
MM1024 N_VPWR_M1024_d N_A_1874_543#_M1024_g N_A_3129_479#_M1024_s N_VPB_M1017_b
+ PHV L=0.5 W=0.75 AD=0.1575 AS=0.21375 PD=1.19571 PS=2.07 NRD=29.2803 NRS=0 M=1
+ R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1015 N_Q_M1015_d N_A_3129_479#_M1015_g N_VPWR_M1024_d N_VPB_M1017_b PHV L=0.5
+ W=1 AD=0.285 AS=0.21 PD=2.57 PS=1.59429 NRD=0 NRS=0 M=1 R=2 SA=250001
+ SB=250000 A=0.5 P=3 MULT=1
DX34_noxref N_VNB_M1023_b N_VPB_M1017_b NWDIODE A=45.137 P=43.04
*
.include "sky130_fd_sc_hvl__dfsbp_1.pxi.spice"
*
.ends
*
*
