* File: sky130_fd_sc_hvl__lsbufhv2hv_hl_1.pxi.spice
* Created: Fri Aug 28 09:36:36 2020
* 
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%VNB N_VNB_M0_noxref_b VNB VNB N_VNB_c_7_p
+ VNB PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%VNB
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%VPB N_VPB_X4_noxref_D1 N_VPB_X6_noxref_D1
+ VPB N_VPB_c_25_n N_VPB_c_26_n N_VPB_c_27_n
+ PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%VPB
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%LOWHVPWR N_LOWHVPWR_M1003_d
+ N_LOWHVPWR_M1003_b N_LOWHVPWR_c_48_n N_LOWHVPWR_c_49_n LOWHVPWR
+ N_LOWHVPWR_c_52_n PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%LOWHVPWR
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%A_662_81# N_A_662_81#_M1_noxref_d
+ N_A_662_81#_M1001_d N_A_662_81#_M0_noxref_g N_A_662_81#_M1003_g
+ N_A_662_81#_c_79_n N_A_662_81#_c_80_n N_A_662_81#_c_82_n N_A_662_81#_c_95_n
+ N_A_662_81#_c_83_n N_A_662_81#_c_84_n N_A_662_81#_c_85_n
+ PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%A_662_81#
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%A A A A N_A_M1_noxref_g N_A_c_126_n
+ N_A_M1001_g PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%A
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%X N_X_M0_noxref_s N_X_M1003_s X X X X X X
+ X N_X_c_141_n PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%X
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%VGND N_VGND_M0_noxref_d VGND VGND
+ N_VGND_c_162_n PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%VGND
cc_1 N_VNB_M0_noxref_b N_VPB_c_25_n 0.0021751f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_2 N_VNB_M0_noxref_b N_VPB_c_26_n 0.0021751f $X=-0.33 $Y=-0.265 $X2=8.4
+ $Y2=4.07
cc_3 N_VNB_M0_noxref_b N_VPB_c_27_n 0.0830934f $X=-0.33 $Y=-0.265 $X2=8.4
+ $Y2=4.07
cc_4 N_VNB_M0_noxref_b LOWHVPWR 0.211657f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_5 N_VNB_M0_noxref_b N_A_662_81#_c_79_n 0.0211189f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_6 N_VNB_M0_noxref_b N_A_662_81#_c_80_n 0.0479081f $X=-0.33 $Y=-0.265 $X2=8.4
+ $Y2=4.07
cc_7 N_VNB_c_7_p N_A_662_81#_c_80_n 5.81195e-19 $X=0.24 $Y=0 $X2=8.4 $Y2=4.07
cc_8 N_VNB_M0_noxref_b N_A_662_81#_c_82_n 0.0140542f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_9 N_VNB_M0_noxref_b N_A_662_81#_c_83_n 0.0588473f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_10 N_VNB_M0_noxref_b N_A_662_81#_c_84_n 0.00770964f $X=-0.33 $Y=-0.265
+ $X2=8.4 $Y2=4.07
cc_11 N_VNB_M0_noxref_b N_A_662_81#_c_85_n 0.0476113f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_c_7_p N_A_662_81#_c_85_n 0.00119158f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_13 N_VNB_M0_noxref_b N_A_M1_noxref_g 0.130438f $X=-0.33 $Y=-0.265 $X2=7.425
+ $Y2=1.885
cc_14 N_VNB_c_7_p N_A_M1_noxref_g 0.00137776f $X=0.24 $Y=0 $X2=7.425 $Y2=1.885
cc_15 N_VNB_M0_noxref_b N_X_c_141_n 0.0673249f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_16 N_VNB_c_7_p N_X_c_141_n 0.00111241f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_17 N_VNB_M0_noxref_b VGND 0.437967f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_18 N_VNB_c_7_p VGND 0.924781f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_19 N_VNB_M0_noxref_b VGND 0.545305f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_20 VNB VGND 0.925009f $X=0 $Y=8.025 $X2=0 $Y2=0
cc_21 N_VNB_M0_noxref_b N_VGND_c_162_n 0.0503123f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_22 N_VNB_c_7_p N_VGND_c_162_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_23 N_VNB_M0_noxref_b VPWR 0.098711f $X=-0.33 $Y=-0.265 $X2=0 $Y2=3.985
cc_24 N_VNB_M0_noxref_b VPWR 0.224313f $X=-0.33 $Y=-0.265 $X2=7.755 $Y2=3.985
cc_25 N_VPB_c_27_n N_LOWHVPWR_M1003_b 0.0270352f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_26 N_VPB_c_27_n N_LOWHVPWR_c_48_n 0.0319699f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_27 N_VPB_c_27_n N_LOWHVPWR_c_49_n 0.00818046f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_28 N_VPB_X4_noxref_D1 LOWHVPWR 0.050189f $X=-0.33 $Y=1.885 $X2=0.24 $Y2=0
cc_29 N_VPB_X6_noxref_D1 LOWHVPWR 0.0721485f $X=7.425 $Y=1.885 $X2=0.24 $Y2=0
cc_30 N_VPB_c_27_n N_LOWHVPWR_c_52_n 0.044651f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_31 N_VPB_c_27_n N_A_662_81#_M1003_g 0.00472565f $X=8.4 $Y=4.07 $X2=0
+ $Y2=8.025
cc_32 N_VPB_c_27_n N_X_c_141_n 0.0201335f $X=8.4 $Y=4.07 $X2=8.4 $Y2=0
cc_33 N_VPB_X4_noxref_D1 VPWR 0.0336658f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_34 N_VPB_X6_noxref_D1 VPWR 0.0422033f $X=7.425 $Y=1.885 $X2=0 $Y2=0
cc_35 N_VPB_c_25_n VPWR 0.00613319f $X=0.24 $Y=4.07 $X2=0 $Y2=0
cc_36 N_VPB_c_26_n VPWR 0.00931478f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_37 N_VPB_c_27_n VPWR 0.914101f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_38 N_VPB_X4_noxref_D1 VPWR 0.0565882f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_39 N_VPB_X6_noxref_D1 VPWR 0.078157f $X=7.425 $Y=1.885 $X2=0 $Y2=0
cc_40 N_VPB_c_25_n VPWR 0.00613319f $X=0.24 $Y=4.07 $X2=0 $Y2=0
cc_41 N_VPB_c_26_n VPWR 0.00931478f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_42 N_VPB_c_27_n VPWR 0.910625f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_43 LOWHVPWR N_A_662_81#_M1001_d 0.00215632f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_44 N_LOWHVPWR_M1003_b N_A_662_81#_M1003_g 0.0931955f $X=2.8 $Y=1.885 $X2=0
+ $Y2=8.025
cc_45 N_LOWHVPWR_c_49_n N_A_662_81#_M1003_g 0.00639755f $X=3.875 $Y=4.265 $X2=0
+ $Y2=8.025
cc_46 LOWHVPWR N_A_662_81#_M1003_g 0.00840344f $X=0.07 $Y=3.02 $X2=0 $Y2=8.025
cc_47 N_LOWHVPWR_c_52_n N_A_662_81#_M1003_g 0.0895392f $X=4.055 $Y=2.65 $X2=0
+ $Y2=8.025
cc_48 N_LOWHVPWR_M1003_b N_A_662_81#_c_82_n 0.0590451f $X=2.8 $Y=1.885 $X2=0
+ $Y2=0
cc_49 LOWHVPWR N_A_662_81#_c_82_n 0.0426117f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_50 N_LOWHVPWR_c_52_n N_A_662_81#_c_95_n 0.0132268f $X=4.055 $Y=2.65 $X2=0
+ $Y2=0
cc_51 N_LOWHVPWR_M1003_b N_A_662_81#_c_83_n 0.00472629f $X=2.8 $Y=1.885 $X2=0.24
+ $Y2=8.14
cc_52 N_LOWHVPWR_M1003_b N_A_M1_noxref_g 0.0998977f $X=2.8 $Y=1.885 $X2=0 $Y2=0
cc_53 LOWHVPWR N_A_M1_noxref_g 0.0214753f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_54 N_LOWHVPWR_c_52_n N_A_M1_noxref_g 0.0171228f $X=4.055 $Y=2.65 $X2=0 $Y2=0
cc_55 LOWHVPWR N_A_c_126_n 0.0167112f $X=0.07 $Y=3.02 $X2=0 $Y2=8.025
cc_56 N_LOWHVPWR_c_52_n N_A_c_126_n 0.0339226f $X=4.055 $Y=2.65 $X2=0 $Y2=8.025
cc_57 LOWHVPWR N_X_M1003_s 8.77815e-19 $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_58 N_LOWHVPWR_M1003_b N_X_c_141_n 0.0876553f $X=2.8 $Y=1.885 $X2=8.4 $Y2=0
cc_59 N_LOWHVPWR_c_49_n N_X_c_141_n 0.0162127f $X=3.875 $Y=4.265 $X2=8.4 $Y2=0
cc_60 LOWHVPWR N_X_c_141_n 0.053365f $X=0.07 $Y=3.02 $X2=8.4 $Y2=0
cc_61 N_LOWHVPWR_c_52_n N_X_c_141_n 0.0750012f $X=4.055 $Y=2.65 $X2=8.4 $Y2=0
cc_62 N_LOWHVPWR_M1003_d VPWR 2.12955e-19 $X=3.915 $Y=2.525 $X2=0 $Y2=0
cc_63 N_LOWHVPWR_M1003_b VPWR 0.0276466f $X=2.8 $Y=1.885 $X2=0 $Y2=0
cc_64 LOWHVPWR VPWR 0.909182f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_65 N_LOWHVPWR_c_52_n VPWR 0.0575297f $X=4.055 $Y=2.65 $X2=0 $Y2=0
cc_66 N_LOWHVPWR_M1003_b VPWR 0.0345944f $X=2.8 $Y=1.885 $X2=0 $Y2=0
cc_67 N_LOWHVPWR_c_48_n VPWR 0.0991109f $X=4.89 $Y=4.38 $X2=0 $Y2=0
cc_68 N_LOWHVPWR_c_49_n VPWR 0.117504f $X=3.875 $Y=4.265 $X2=0 $Y2=0
cc_69 N_A_662_81#_c_79_n N_A_M1_noxref_g 0.0418619f $X=4.865 $Y=1.52 $X2=0 $Y2=0
cc_70 N_A_662_81#_c_80_n N_A_M1_noxref_g 0.0193356f $X=4.95 $Y=0.745 $X2=0 $Y2=0
cc_71 N_A_662_81#_c_82_n N_A_M1_noxref_g 0.0357848f $X=4.95 $Y=2.65 $X2=0 $Y2=0
cc_72 N_A_662_81#_c_95_n N_A_M1_noxref_g 0.00239611f $X=3.73 $Y=1.56 $X2=0 $Y2=0
cc_73 N_A_662_81#_c_83_n N_A_M1_noxref_g 0.0524552f $X=3.73 $Y=1.56 $X2=0 $Y2=0
cc_74 N_A_662_81#_c_85_n N_A_M1_noxref_g 0.014314f $X=3.612 $Y=1.395 $X2=0 $Y2=0
cc_75 N_A_662_81#_c_79_n N_A_c_126_n 0.0249855f $X=4.865 $Y=1.52 $X2=0 $Y2=8.025
cc_76 N_A_662_81#_c_82_n N_A_c_126_n 0.0690189f $X=4.95 $Y=2.65 $X2=0 $Y2=8.025
cc_77 N_A_662_81#_c_95_n N_A_c_126_n 0.00968782f $X=3.73 $Y=1.56 $X2=0 $Y2=8.025
cc_78 N_A_662_81#_c_83_n N_A_c_126_n 0.00385482f $X=3.73 $Y=1.56 $X2=0 $Y2=8.025
cc_79 N_A_662_81#_M1003_g N_X_c_141_n 0.0314398f $X=3.665 $Y=3.275 $X2=8.4 $Y2=0
cc_80 N_A_662_81#_c_95_n N_X_c_141_n 0.0494349f $X=3.73 $Y=1.56 $X2=8.4 $Y2=0
cc_81 N_A_662_81#_c_83_n N_X_c_141_n 0.0245808f $X=3.73 $Y=1.56 $X2=8.4 $Y2=0
cc_82 N_A_662_81#_c_85_n N_X_c_141_n 0.0280292f $X=3.612 $Y=1.395 $X2=8.4 $Y2=0
cc_83 N_A_662_81#_M1_noxref_d VGND 0.00221032f $X=4.81 $Y=0.535 $X2=0 $Y2=0
cc_84 N_A_662_81#_c_80_n VGND 0.028425f $X=4.95 $Y=0.745 $X2=0 $Y2=0
cc_85 N_A_662_81#_c_85_n VGND 0.0119319f $X=3.612 $Y=1.395 $X2=0 $Y2=0
cc_86 N_A_662_81#_c_79_n N_VGND_c_162_n 0.0501274f $X=4.865 $Y=1.52 $X2=-0.33
+ $Y2=-0.265
cc_87 N_A_662_81#_c_80_n N_VGND_c_162_n 0.0257644f $X=4.95 $Y=0.745 $X2=-0.33
+ $Y2=-0.265
cc_88 N_A_662_81#_c_95_n N_VGND_c_162_n 0.0253119f $X=3.73 $Y=1.56 $X2=-0.33
+ $Y2=-0.265
cc_89 N_A_662_81#_c_83_n N_VGND_c_162_n 0.00281087f $X=3.73 $Y=1.56 $X2=-0.33
+ $Y2=-0.265
cc_90 N_A_662_81#_c_85_n N_VGND_c_162_n 0.0490642f $X=3.612 $Y=1.395 $X2=-0.33
+ $Y2=-0.265
cc_91 N_A_662_81#_M1003_g VPWR 0.00273887f $X=3.665 $Y=3.275 $X2=0 $Y2=0
cc_92 N_A_662_81#_c_82_n VPWR 0.00859591f $X=4.95 $Y=2.65 $X2=0 $Y2=0
cc_93 N_A_M1_noxref_g VGND 0.0202943f $X=4.56 $Y=0.745 $X2=0 $Y2=0
cc_94 N_A_M1_noxref_g N_VGND_c_162_n 0.0450534f $X=4.56 $Y=0.745 $X2=-0.33
+ $Y2=-0.265
cc_95 N_A_M1_noxref_g VPWR 0.0102904f $X=4.56 $Y=0.745 $X2=0 $Y2=0
cc_96 N_X_c_141_n VGND 0.0404606f $X=3.17 $Y=0.68 $X2=0 $Y2=0
cc_97 N_X_c_141_n N_VGND_c_162_n 0.0600788f $X=3.17 $Y=0.68 $X2=-0.33 $Y2=-0.265
cc_98 N_X_M1003_s VPWR 2.45755e-19 $X=3.13 $Y=2.525 $X2=0 $Y2=0
cc_99 N_X_c_141_n VPWR 0.0437272f $X=3.17 $Y=0.68 $X2=0 $Y2=0
cc_100 N_X_c_141_n VPWR 9.68375e-19 $X=3.17 $Y=0.68 $X2=0 $Y2=0
