* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__probe_p_8 A VGND VNB VPB VPWR X
M1000 X a_45_443# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=1.68e+12p pd=1.424e+07u as=2.9175e+12p ps=2.189e+07u
M1001 X a_45_443# VGND VNB nhv w=750000u l=500000u
+  ad=8.4e+11p pd=8.24e+06u as=1.45875e+12p ps=1.289e+07u
M1002 VGND a_45_443# X VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_45_443# A VGND VNB nhv w=750000u l=500000u
+  ad=4.2375e+11p pd=4.13e+06u as=0p ps=0u
M1004 X a_45_443# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_45_443# X VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_45_443# VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=8.475e+11p ps=7.13e+06u
M1007 VPWR A a_45_443# VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A a_45_443# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_45_443# VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_45_443# X VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_45_443# X VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_45_443# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_45_443# VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_45_443# X VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A a_45_443# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_45_443# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_45_443# X VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_45_443# X VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_45_443# A VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_45_443# X VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_45_443# VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
