* File: sky130_fd_sc_hvl__conb_1.pex.spice
* Created: Wed Sep  2 09:04:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__CONB_1%VNB 5 7 11 25
r18 7 25 5.20833e-05 $w=2.4e-06 $l=1e-09 $layer=MET1_cond $X=1.2 $Y=0.057
+ $X2=1.2 $Y2=0.058
r19 7 11 0.00296875 $w=2.4e-06 $l=5.7e-08 $layer=MET1_cond $X=1.2 $Y=0.057
+ $X2=1.2 $Y2=0
r20 5 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r21 5 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__CONB_1%VPB 4 6 14 21
r21 10 21 0.00296875 $w=2.4e-06 $l=5.7e-08 $layer=MET1_cond $X=1.2 $Y=4.07
+ $X2=1.2 $Y2=4.013
r22 10 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=4.07
+ $X2=2.16 $Y2=4.07
r23 9 14 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=2.16 $Y2=4.07
r24 9 10 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r25 6 21 5.20833e-05 $w=2.4e-06 $l=1e-09 $layer=MET1_cond $X=1.2 $Y=4.012
+ $X2=1.2 $Y2=4.013
r26 4 14 72.8 $w=1.7e-07 $l=2.20209e-06 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=2.16 $Y2=4.07
r27 4 9 72.8 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__CONB_1%HI 2 4 6 10 11 12 13 20
c37 2 0 1.59574e-19 $X=0.84 $Y=1.82
r38 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=2.775 $X2=1.2
+ $Y2=3.145
r39 11 12 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=2.405 $X2=1.2
+ $Y2=2.775
r40 11 22 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=1.2 $Y=2.405 $X2=1.2
+ $Y2=2.185
r41 10 22 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.2 $Y=2.06 $X2=1.2
+ $Y2=2.185
r42 10 30 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=1.2 $Y=2.06 $X2=0.74
+ $Y2=2.06
r43 7 20 30.7442 $w=6.7e-07 $l=3.85e-07 $layer=POLY_cond $X=0.455 $Y=0.735
+ $X2=0.84 $Y2=0.735
r44 6 9 14.3948 $w=5.73e-07 $l=5.05e-07 $layer=LI1_cond $X=0.577 $Y=0.565
+ $X2=0.577 $Y2=1.07
r45 6 7 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.455
+ $Y=0.565 $X2=0.455 $Y2=0.565
r46 4 30 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.74 $Y=1.935
+ $X2=0.74 $Y2=2.06
r47 4 9 39.8745 $w=2.48e-07 $l=8.65e-07 $layer=LI1_cond $X=0.74 $Y=1.935
+ $X2=0.74 $Y2=1.07
r48 1 20 9.23499 $w=5.1e-07 $l=3.35e-07 $layer=POLY_cond $X=0.84 $Y=1.07
+ $X2=0.84 $Y2=0.735
r49 1 2 78.6808 $w=5.1e-07 $l=7.5e-07 $layer=POLY_cond $X=0.84 $Y=1.07 $X2=0.84
+ $Y2=1.82
.ends

.subckt PM_SKY130_FD_SC_HVL__CONB_1%VPWR 1 2 3 7 9
r25 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.59
+ $X2=0.72 $Y2=3.59
r26 7 13 6.36417 $w=5.08e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=3.48
+ $X2=0.72 $Y2=3.48
r27 6 9 30.7442 $w=6.7e-07 $l=3.85e-07 $layer=POLY_cond $X=0.455 $Y=3.51
+ $X2=0.84 $Y2=3.51
r28 6 7 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.455 $Y=3.34
+ $X2=0.455 $Y2=3.34
r29 3 14 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.63 $X2=0.72
+ $Y2=3.63
r30 2 9 9.23499 $w=5.1e-07 $l=3.35e-07 $layer=POLY_cond $X=0.84 $Y=3.175
+ $X2=0.84 $Y2=3.51
r31 1 2 137.429 $w=5.1e-07 $l=1.31e-06 $layer=POLY_cond $X=0.84 $Y=1.865
+ $X2=0.84 $Y2=3.175
.ends

.subckt PM_SKY130_FD_SC_HVL__CONB_1%VGND 2 5 10 11 16 17
r25 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.04 $Y=0.48
+ $X2=2.04 $Y2=0.48
r26 11 16 3.22006 $w=3.38e-07 $l=9.5e-08 $layer=LI1_cond $X=1.945 $Y=0.455
+ $X2=2.04 $Y2=0.455
r27 10 11 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.945
+ $Y=0.565 $X2=1.945 $Y2=0.565
r28 7 10 30.7442 $w=6.7e-07 $l=3.85e-07 $layer=POLY_cond $X=1.56 $Y=0.735
+ $X2=1.945 $Y2=0.735
r29 5 17 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=1.2 $Y=0.44 $X2=2.04
+ $Y2=0.44
r30 1 7 9.23499 $w=5.1e-07 $l=3.35e-07 $layer=POLY_cond $X=1.56 $Y=1.07 $X2=1.56
+ $Y2=0.735
r31 1 2 78.6808 $w=5.1e-07 $l=7.5e-07 $layer=POLY_cond $X=1.56 $Y=1.07 $X2=1.56
+ $Y2=1.82
.ends

.subckt PM_SKY130_FD_SC_HVL__CONB_1%LO 1 2 5 6 9 10 11 12 13
c40 13 0 1.59574e-19 $X=1.68 $Y=2.035
r41 29 35 0.73951 $w=2.65e-07 $l=1.33e-07 $layer=LI1_cond $X=1.662 $Y=1.765
+ $X2=1.662 $Y2=1.632
r42 13 29 11.7419 $w=2.63e-07 $l=2.7e-07 $layer=LI1_cond $X=1.662 $Y=2.035
+ $X2=1.662 $Y2=1.765
r43 12 35 0.782791 $w=2.63e-07 $l=1.8e-08 $layer=LI1_cond $X=1.68 $Y=1.632
+ $X2=1.662 $Y2=1.632
r44 11 35 20.0916 $w=2.63e-07 $l=4.62e-07 $layer=LI1_cond $X=1.2 $Y=1.632
+ $X2=1.662 $Y2=1.632
r45 10 11 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.2 $Y=1.295
+ $X2=1.2 $Y2=1.5
r46 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=0.925 $X2=1.2
+ $Y2=1.295
r47 7 13 49.5768 $w=2.63e-07 $l=1.14e-06 $layer=LI1_cond $X=1.662 $Y=3.175
+ $X2=1.662 $Y2=2.035
r48 6 19 30.7442 $w=6.7e-07 $l=3.85e-07 $layer=POLY_cond $X=1.945 $Y=3.51
+ $X2=1.56 $Y2=3.51
r49 5 7 6.96725 $w=5.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.82 $Y=3.34 $X2=1.82
+ $Y2=3.175
r50 5 6 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.945 $Y=3.34
+ $X2=1.945 $Y2=3.34
r51 2 19 9.23499 $w=5.1e-07 $l=3.35e-07 $layer=POLY_cond $X=1.56 $Y=3.175
+ $X2=1.56 $Y2=3.51
r52 1 2 137.429 $w=5.1e-07 $l=1.31e-06 $layer=POLY_cond $X=1.56 $Y=1.865
+ $X2=1.56 $Y2=3.175
.ends

