* File: sky130_fd_sc_hvl__schmittbuf_1.pxi.spice
* Created: Wed Sep  2 09:09:49 2020
* 
x_PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%VNB N_VNB_M1001_b VNB N_VNB_c_4_p VNB
+ PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%VNB
x_PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%VPB N_VPB_M1006_b VPB N_VPB_c_35_p VPB
+ PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%VPB
x_PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_117_181# N_A_117_181#_M1007_s
+ N_A_117_181#_M1005_s N_A_117_181#_c_73_n N_A_117_181#_M1006_g
+ N_A_117_181#_c_74_n N_A_117_181#_M1000_g N_A_117_181#_M1004_g
+ N_A_117_181#_M1001_g N_A_117_181#_c_112_p N_A_117_181#_c_77_n
+ N_A_117_181#_c_78_n N_A_117_181#_c_79_n N_A_117_181#_c_90_n
+ N_A_117_181#_c_91_n N_A_117_181#_c_80_n N_A_117_181#_c_81_n
+ PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_117_181#
x_PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A N_A_M1007_g N_A_M1005_g N_A_c_160_n
+ N_A_M1003_g N_A_M1002_g A A A PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A
x_PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_78_463# N_A_78_463#_X8_noxref_D1
+ N_A_78_463#_M1006_s N_A_78_463#_c_204_n N_A_78_463#_c_199_n
+ N_A_78_463#_c_200_n N_A_78_463#_c_202_n N_A_78_463#_c_205_n
+ PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_78_463#
x_PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_64_207# N_A_64_207#_M1001_s
+ N_A_64_207#_X9_noxref_D0 N_A_64_207#_c_232_n N_A_64_207#_c_233_n
+ N_A_64_207#_c_236_n N_A_64_207#_c_230_n N_A_64_207#_c_231_n
+ N_A_64_207#_c_240_n PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_64_207#
x_PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_231_463# N_A_231_463#_M1006_d
+ N_A_231_463#_M1005_d N_A_231_463#_c_262_n N_A_231_463#_c_263_n
+ N_A_231_463#_c_265_n N_A_231_463#_c_267_n
+ PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_231_463#
x_PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%VPWR N_VPWR_M1002_d VPWR N_VPWR_c_287_n
+ N_VPWR_c_290_n PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%VPWR
x_PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%X N_X_M1000_d N_X_M1004_d X X X X X X X
+ N_X_c_314_n PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%X
x_PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_217_207# N_A_217_207#_M1001_d
+ N_A_217_207#_M1007_d N_A_217_207#_c_328_n N_A_217_207#_c_329_n
+ N_A_217_207#_c_330_n PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_217_207#
x_PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%VGND N_VGND_M1003_d VGND N_VGND_c_354_n
+ N_VGND_c_356_n PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%VGND
cc_1 N_VNB_M1001_b N_A_117_181#_c_73_n 0.0776594f $X=-0.33 $Y=-0.265 $X2=0.905
+ $Y2=1.985
cc_2 N_VNB_M1001_b N_A_117_181#_c_74_n 0.0298979f $X=-0.33 $Y=-0.265 $X2=4.615
+ $Y2=1.725
cc_3 N_VNB_M1001_b N_A_117_181#_M1000_g 0.0928973f $X=-0.33 $Y=-0.265 $X2=4.615
+ $Y2=0.91
cc_4 N_VNB_c_4_p N_A_117_181#_M1000_g 0.00112492f $X=0.24 $Y=0 $X2=4.615
+ $Y2=0.91
cc_5 N_VNB_M1001_b N_A_117_181#_c_77_n 0.0333783f $X=-0.33 $Y=-0.265 $X2=1.47
+ $Y2=1.82
cc_6 N_VNB_M1001_b N_A_117_181#_c_78_n 0.00889381f $X=-0.33 $Y=-0.265 $X2=1.745
+ $Y2=1.985
cc_7 N_VNB_M1001_b N_A_117_181#_c_79_n 0.00193849f $X=-0.33 $Y=-0.265 $X2=4.605
+ $Y2=1.89
cc_8 N_VNB_M1001_b N_A_117_181#_c_80_n 0.0192231f $X=-0.33 $Y=-0.265 $X2=3.855
+ $Y2=1.78
cc_9 N_VNB_M1001_b N_A_117_181#_c_81_n 0.0108238f $X=-0.33 $Y=-0.265 $X2=4.21
+ $Y2=1.78
cc_10 N_VNB_M1001_b N_A_M1007_g 0.0425834f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_11 N_VNB_M1001_b N_A_c_160_n 0.0508346f $X=-0.33 $Y=-0.265 $X2=0.905 $Y2=2.69
cc_12 N_VNB_M1001_b N_A_M1003_g 0.0486113f $X=-0.33 $Y=-0.265 $X2=4.615
+ $Y2=1.725
cc_13 N_VNB_M1001_b A 0.00288218f $X=-0.33 $Y=-0.265 $X2=0.87 $Y2=1.245
cc_14 N_VNB_M1001_b N_A_78_463#_c_199_n 0.00748908f $X=-0.33 $Y=-0.265 $X2=4.615
+ $Y2=0.91
cc_15 N_VNB_M1001_b N_A_78_463#_c_200_n 0.0137608f $X=-0.33 $Y=-0.265 $X2=4.615
+ $Y2=0.91
cc_16 N_VNB_c_4_p N_A_78_463#_c_200_n 3.587e-19 $X=0.24 $Y=0 $X2=4.615 $Y2=0.91
cc_17 N_VNB_M1001_b N_A_78_463#_c_202_n 0.045508f $X=-0.33 $Y=-0.265 $X2=4.615
+ $Y2=2.055
cc_18 N_VNB_c_4_p N_A_78_463#_c_202_n 0.00244368f $X=0.24 $Y=0 $X2=4.615
+ $Y2=2.055
cc_19 N_VNB_M1001_b N_A_64_207#_c_230_n 0.0122625f $X=-0.33 $Y=-0.265 $X2=4.615
+ $Y2=1.725
cc_20 N_VNB_M1001_b N_A_64_207#_c_231_n 0.0329411f $X=-0.33 $Y=-0.265 $X2=4.615
+ $Y2=0.91
cc_21 N_VNB_M1001_b N_X_c_314_n 0.0648184f $X=-0.33 $Y=-0.265 $X2=1.155
+ $Y2=1.815
cc_22 N_VNB_c_4_p N_X_c_314_n 7.67181e-19 $X=0.24 $Y=0 $X2=1.155 $Y2=1.815
cc_23 N_VNB_M1001_b N_A_217_207#_c_328_n 0.0153652f $X=-0.33 $Y=-0.265 $X2=0.905
+ $Y2=1.985
cc_24 N_VNB_M1001_b N_A_217_207#_c_329_n 0.00721573f $X=-0.33 $Y=-0.265
+ $X2=0.905 $Y2=2.69
cc_25 N_VNB_M1001_b N_A_217_207#_c_330_n 0.0051476f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_26 N_VNB_M1001_b N_VGND_c_354_n 0.0906178f $X=-0.33 $Y=-0.265 $X2=0.905
+ $Y2=1.985
cc_27 N_VNB_c_4_p N_VGND_c_354_n 0.0042154f $X=0.24 $Y=0 $X2=0.905 $Y2=1.985
cc_28 N_VNB_M1001_b N_VGND_c_356_n 0.121252f $X=-0.33 $Y=-0.265 $X2=4.615
+ $Y2=1.725
cc_29 N_VNB_c_4_p N_VGND_c_356_n 0.564953f $X=0.24 $Y=0 $X2=4.615 $Y2=1.725
cc_30 N_VPB_M1006_b N_A_117_181#_c_73_n 0.0078896f $X=-0.33 $Y=1.885 $X2=0.905
+ $Y2=1.985
cc_31 N_VPB_M1006_b N_A_117_181#_M1006_g 0.0663052f $X=-0.33 $Y=1.885 $X2=0.905
+ $Y2=2.69
cc_32 N_VPB_M1006_b N_A_117_181#_c_74_n 0.0305058f $X=-0.33 $Y=1.885 $X2=4.615
+ $Y2=1.725
cc_33 N_VPB_M1006_b N_A_117_181#_M1004_g 0.0509878f $X=-0.33 $Y=1.885 $X2=4.615
+ $Y2=2.965
cc_34 VPB N_A_117_181#_M1004_g 0.00970178f $X=0 $Y=3.955 $X2=4.615 $Y2=2.965
cc_35 N_VPB_c_35_p N_A_117_181#_M1004_g 0.0172225f $X=5.04 $Y=4.07 $X2=4.615
+ $Y2=2.965
cc_36 N_VPB_M1006_b N_A_117_181#_c_77_n 0.0198216f $X=-0.33 $Y=1.885 $X2=1.47
+ $Y2=1.82
cc_37 N_VPB_M1006_b N_A_117_181#_c_78_n 0.00229781f $X=-0.33 $Y=1.885 $X2=1.745
+ $Y2=1.985
cc_38 N_VPB_M1006_b N_A_117_181#_c_90_n 0.00958261f $X=-0.33 $Y=1.885 $X2=1.845
+ $Y2=2.46
cc_39 N_VPB_M1006_b N_A_117_181#_c_91_n 0.00779824f $X=-0.33 $Y=1.885 $X2=1.832
+ $Y2=2.33
cc_40 N_VPB_M1006_b N_A_117_181#_c_81_n 0.00391011f $X=-0.33 $Y=1.885 $X2=4.21
+ $Y2=1.78
cc_41 N_VPB_M1006_b N_A_M1005_g 0.0418906f $X=-0.33 $Y=1.885 $X2=0.905 $Y2=1.985
cc_42 N_VPB_M1006_b N_A_c_160_n 0.0353943f $X=-0.33 $Y=1.885 $X2=0.905 $Y2=2.69
cc_43 N_VPB_M1006_b N_A_M1002_g 0.0514285f $X=-0.33 $Y=1.885 $X2=4.615 $Y2=2.055
cc_44 N_VPB_M1006_b A 0.00806722f $X=-0.33 $Y=1.885 $X2=0.87 $Y2=1.245
cc_45 N_VPB_M1006_b N_A_78_463#_c_204_n 0.00277455f $X=-0.33 $Y=1.885 $X2=0.905
+ $Y2=2.69
cc_46 N_VPB_M1006_b N_A_78_463#_c_205_n 0.00544011f $X=-0.33 $Y=1.885 $X2=0.87
+ $Y2=1.245
cc_47 N_VPB_M1006_b N_A_64_207#_c_232_n 0.0783095f $X=-0.33 $Y=1.885 $X2=0.905
+ $Y2=2.69
cc_48 N_VPB_M1006_b N_A_64_207#_c_233_n 0.0105695f $X=-0.33 $Y=1.885 $X2=0.905
+ $Y2=2.69
cc_49 VPB N_A_64_207#_c_233_n 0.00130475f $X=0 $Y=3.955 $X2=0.905 $Y2=2.69
cc_50 N_VPB_c_35_p N_A_64_207#_c_233_n 0.0170967f $X=5.04 $Y=4.07 $X2=0.905
+ $Y2=2.69
cc_51 N_VPB_M1006_b N_A_64_207#_c_236_n 0.00427244f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_52 VPB N_A_64_207#_c_236_n 4.57356e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_53 N_VPB_c_35_p N_A_64_207#_c_236_n 0.00616416f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_54 N_VPB_M1006_b N_A_64_207#_c_230_n 0.0129021f $X=-0.33 $Y=1.885 $X2=4.615
+ $Y2=1.725
cc_55 N_VPB_M1006_b N_A_64_207#_c_240_n 0.00808015f $X=-0.33 $Y=1.885 $X2=0.835
+ $Y2=1.245
cc_56 VPB N_A_64_207#_c_240_n 8.70177e-19 $X=0 $Y=3.955 $X2=0.835 $Y2=1.245
cc_57 N_VPB_c_35_p N_A_64_207#_c_240_n 0.0138665f $X=5.04 $Y=4.07 $X2=0.835
+ $Y2=1.245
cc_58 N_VPB_M1006_b N_A_231_463#_c_262_n 0.0168314f $X=-0.33 $Y=1.885 $X2=0.905
+ $Y2=2.69
cc_59 N_VPB_M1006_b N_A_231_463#_c_263_n 0.0365505f $X=-0.33 $Y=1.885 $X2=4.615
+ $Y2=1.725
cc_60 N_VPB_c_35_p N_A_231_463#_c_263_n 0.0183157f $X=5.04 $Y=4.07 $X2=4.615
+ $Y2=1.725
cc_61 N_VPB_M1006_b N_A_231_463#_c_265_n 0.0115049f $X=-0.33 $Y=1.885 $X2=4.615
+ $Y2=0.91
cc_62 N_VPB_c_35_p N_A_231_463#_c_265_n 0.00385317f $X=5.04 $Y=4.07 $X2=4.615
+ $Y2=0.91
cc_63 N_VPB_M1006_b N_A_231_463#_c_267_n 0.00199424f $X=-0.33 $Y=1.885 $X2=4.615
+ $Y2=2.055
cc_64 N_VPB_M1006_b N_VPWR_c_287_n 0.0210333f $X=-0.33 $Y=1.885 $X2=4.615
+ $Y2=0.91
cc_65 VPB N_VPWR_c_287_n 0.00465345f $X=0 $Y=3.955 $X2=4.615 $Y2=0.91
cc_66 N_VPB_c_35_p N_VPWR_c_287_n 0.0690836f $X=5.04 $Y=4.07 $X2=4.615 $Y2=0.91
cc_67 N_VPB_M1006_b N_VPWR_c_290_n 0.0696609f $X=-0.33 $Y=1.885 $X2=4.615
+ $Y2=2.055
cc_68 VPB N_VPWR_c_290_n 0.563914f $X=0 $Y=3.955 $X2=4.615 $Y2=2.055
cc_69 N_VPB_c_35_p N_VPWR_c_290_n 0.0247309f $X=5.04 $Y=4.07 $X2=4.615 $Y2=2.055
cc_70 N_VPB_M1006_b N_X_c_314_n 0.0684789f $X=-0.33 $Y=1.885 $X2=1.155 $Y2=1.815
cc_71 VPB N_X_c_314_n 9.65216e-19 $X=0 $Y=3.955 $X2=1.155 $Y2=1.815
cc_72 N_VPB_c_35_p N_X_c_314_n 0.0139605f $X=5.04 $Y=4.07 $X2=1.155 $Y2=1.815
cc_73 N_A_117_181#_c_77_n N_A_M1007_g 0.00378861f $X=1.47 $Y=1.82 $X2=0 $Y2=0
cc_74 N_A_117_181#_c_78_n N_A_M1007_g 0.0136782f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_75 N_A_117_181#_c_80_n N_A_M1007_g 0.0268696f $X=3.855 $Y=1.78 $X2=0 $Y2=0
cc_76 N_A_117_181#_c_90_n N_A_M1005_g 0.0211944f $X=1.845 $Y=2.46 $X2=0 $Y2=0
cc_77 N_A_117_181#_c_77_n N_A_c_160_n 0.00853467f $X=1.47 $Y=1.82 $X2=0 $Y2=0
cc_78 N_A_117_181#_c_78_n N_A_c_160_n 0.00508868f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A_117_181#_c_90_n N_A_c_160_n 0.00114415f $X=1.845 $Y=2.46 $X2=0 $Y2=0
cc_80 N_A_117_181#_c_91_n N_A_c_160_n 0.0113114f $X=1.832 $Y=2.33 $X2=0 $Y2=0
cc_81 N_A_117_181#_c_80_n N_A_c_160_n 0.00326629f $X=3.855 $Y=1.78 $X2=0 $Y2=0
cc_82 N_A_117_181#_c_81_n N_A_c_160_n 0.00107435f $X=4.21 $Y=1.78 $X2=0 $Y2=0
cc_83 N_A_117_181#_c_80_n N_A_M1003_g 0.0402166f $X=3.855 $Y=1.78 $X2=0.24 $Y2=0
cc_84 N_A_117_181#_c_81_n N_A_M1003_g 0.00493054f $X=4.21 $Y=1.78 $X2=0.24 $Y2=0
cc_85 N_A_117_181#_c_78_n A 0.0110113f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A_117_181#_c_91_n A 0.0125231f $X=1.832 $Y=2.33 $X2=0 $Y2=0
cc_87 N_A_117_181#_c_80_n A 0.0935709f $X=3.855 $Y=1.78 $X2=0 $Y2=0
cc_88 N_A_117_181#_c_81_n A 0.0081712f $X=4.21 $Y=1.78 $X2=0 $Y2=0
cc_89 N_A_117_181#_M1006_g N_A_78_463#_c_204_n 0.0208075f $X=0.905 $Y=2.69 $X2=0
+ $Y2=0
cc_90 N_A_117_181#_c_73_n N_A_78_463#_c_199_n 0.057566f $X=0.905 $Y=1.985 $X2=0
+ $Y2=0
cc_91 N_A_117_181#_M1006_g N_A_78_463#_c_199_n 0.0129103f $X=0.905 $Y=2.69 $X2=0
+ $Y2=0
cc_92 N_A_117_181#_c_112_p N_A_78_463#_c_199_n 0.0249855f $X=1.6 $Y=1.82 $X2=0
+ $Y2=0
cc_93 N_A_117_181#_c_73_n N_A_78_463#_c_202_n 0.00913541f $X=0.905 $Y=1.985
+ $X2=0 $Y2=0
cc_94 N_A_117_181#_c_73_n N_A_78_463#_c_205_n 0.00190494f $X=0.905 $Y=1.985
+ $X2=0 $Y2=0
cc_95 N_A_117_181#_M1006_g N_A_78_463#_c_205_n 0.024107f $X=0.905 $Y=2.69 $X2=0
+ $Y2=0
cc_96 N_A_117_181#_c_73_n N_A_64_207#_c_232_n 0.00399134f $X=0.905 $Y=1.985
+ $X2=0 $Y2=0
cc_97 N_A_117_181#_M1006_g N_A_64_207#_c_232_n 0.00540047f $X=0.905 $Y=2.69
+ $X2=0 $Y2=0
cc_98 N_A_117_181#_M1006_g N_A_64_207#_c_233_n 0.00253462f $X=0.905 $Y=2.69
+ $X2=0 $Y2=0
cc_99 N_A_117_181#_c_73_n N_A_64_207#_c_230_n 0.00478364f $X=0.905 $Y=1.985
+ $X2=0.24 $Y2=0
cc_100 N_A_117_181#_c_73_n N_A_64_207#_c_231_n 0.00984309f $X=0.905 $Y=1.985
+ $X2=0 $Y2=0
cc_101 N_A_117_181#_M1006_g N_A_64_207#_c_240_n 0.0123235f $X=0.905 $Y=2.69
+ $X2=0 $Y2=0
cc_102 N_A_117_181#_M1006_g N_A_231_463#_c_262_n 0.00827946f $X=0.905 $Y=2.69
+ $X2=0 $Y2=0
cc_103 N_A_117_181#_c_112_p N_A_231_463#_c_262_n 0.0139183f $X=1.6 $Y=1.82 $X2=0
+ $Y2=0
cc_104 N_A_117_181#_c_77_n N_A_231_463#_c_262_n 0.00557092f $X=1.47 $Y=1.82
+ $X2=0 $Y2=0
cc_105 N_A_117_181#_c_91_n N_A_231_463#_c_262_n 0.0573119f $X=1.832 $Y=2.33
+ $X2=0 $Y2=0
cc_106 N_A_117_181#_c_90_n N_A_231_463#_c_263_n 0.0252252f $X=1.845 $Y=2.46
+ $X2=0.24 $Y2=0
cc_107 N_A_117_181#_c_90_n N_A_231_463#_c_267_n 0.0251896f $X=1.845 $Y=2.46
+ $X2=0 $Y2=0
cc_108 N_A_117_181#_c_91_n N_A_231_463#_c_267_n 2.50571e-19 $X=1.832 $Y=2.33
+ $X2=0 $Y2=0
cc_109 N_A_117_181#_c_74_n N_VPWR_c_287_n 0.0057493f $X=4.615 $Y=1.725 $X2=0
+ $Y2=0
cc_110 N_A_117_181#_M1004_g N_VPWR_c_287_n 0.0580959f $X=4.615 $Y=2.965 $X2=0
+ $Y2=0
cc_111 N_A_117_181#_c_80_n N_VPWR_c_287_n 0.0172059f $X=3.855 $Y=1.78 $X2=0
+ $Y2=0
cc_112 N_A_117_181#_c_81_n N_VPWR_c_287_n 0.0416819f $X=4.21 $Y=1.78 $X2=0 $Y2=0
cc_113 N_A_117_181#_M1006_g N_VPWR_c_290_n 0.00631521f $X=0.905 $Y=2.69 $X2=0
+ $Y2=0
cc_114 N_A_117_181#_M1004_g N_VPWR_c_290_n 0.0184324f $X=4.615 $Y=2.965 $X2=0
+ $Y2=0
cc_115 N_A_117_181#_c_74_n N_X_c_314_n 0.0115334f $X=4.615 $Y=1.725 $X2=0 $Y2=0
cc_116 N_A_117_181#_M1000_g N_X_c_314_n 0.0378537f $X=4.615 $Y=0.91 $X2=0 $Y2=0
cc_117 N_A_117_181#_M1004_g N_X_c_314_n 0.0405885f $X=4.615 $Y=2.965 $X2=0 $Y2=0
cc_118 N_A_117_181#_c_79_n N_X_c_314_n 0.032524f $X=4.605 $Y=1.89 $X2=0 $Y2=0
cc_119 N_A_117_181#_c_81_n N_X_c_314_n 0.00420812f $X=4.21 $Y=1.78 $X2=0 $Y2=0
cc_120 N_A_117_181#_c_80_n N_A_217_207#_M1007_d 0.00176773f $X=3.855 $Y=1.78
+ $X2=0 $Y2=0
cc_121 N_A_117_181#_M1007_s N_A_217_207#_c_328_n 0.00230047f $X=1.65 $Y=1.125
+ $X2=0 $Y2=0
cc_122 N_A_117_181#_c_73_n N_A_217_207#_c_328_n 2.48632e-19 $X=0.905 $Y=1.985
+ $X2=0 $Y2=0
cc_123 N_A_117_181#_c_112_p N_A_217_207#_c_328_n 0.00689064f $X=1.6 $Y=1.82
+ $X2=0 $Y2=0
cc_124 N_A_117_181#_c_77_n N_A_217_207#_c_328_n 0.00382318f $X=1.47 $Y=1.82
+ $X2=0 $Y2=0
cc_125 N_A_117_181#_c_78_n N_A_217_207#_c_328_n 0.0228236f $X=1.745 $Y=1.985
+ $X2=0 $Y2=0
cc_126 N_A_117_181#_c_80_n N_A_217_207#_c_328_n 0.0167561f $X=3.855 $Y=1.78
+ $X2=0 $Y2=0
cc_127 N_A_117_181#_c_73_n N_A_217_207#_c_329_n 0.0162495f $X=0.905 $Y=1.985
+ $X2=0 $Y2=0
cc_128 N_A_117_181#_c_112_p N_A_217_207#_c_329_n 0.0178469f $X=1.6 $Y=1.82 $X2=0
+ $Y2=0
cc_129 N_A_117_181#_c_78_n N_A_217_207#_c_329_n 0.006863f $X=1.745 $Y=1.985
+ $X2=0 $Y2=0
cc_130 N_A_117_181#_c_78_n N_A_217_207#_c_330_n 6.85235e-19 $X=1.745 $Y=1.985
+ $X2=0 $Y2=0
cc_131 N_A_117_181#_c_80_n N_A_217_207#_c_330_n 0.0162949f $X=3.855 $Y=1.78
+ $X2=0 $Y2=0
cc_132 N_A_117_181#_c_80_n N_VGND_M1003_d 0.00245157f $X=3.855 $Y=1.78 $X2=0
+ $Y2=0
cc_133 N_A_117_181#_c_74_n N_VGND_c_354_n 0.00132781f $X=4.615 $Y=1.725 $X2=0
+ $Y2=0
cc_134 N_A_117_181#_M1000_g N_VGND_c_354_n 0.0518393f $X=4.615 $Y=0.91 $X2=0
+ $Y2=0
cc_135 N_A_117_181#_c_79_n N_VGND_c_354_n 0.0181508f $X=4.605 $Y=1.89 $X2=0
+ $Y2=0
cc_136 N_A_117_181#_c_80_n N_VGND_c_354_n 0.0723462f $X=3.855 $Y=1.78 $X2=0
+ $Y2=0
cc_137 N_A_117_181#_c_73_n N_VGND_c_356_n 0.00356325f $X=0.905 $Y=1.985 $X2=0.24
+ $Y2=0
cc_138 N_A_117_181#_M1000_g N_VGND_c_356_n 0.0150791f $X=4.615 $Y=0.91 $X2=0.24
+ $Y2=0
cc_139 N_A_M1007_g N_A_78_463#_c_202_n 6.32475e-19 $X=2.165 $Y=1.335 $X2=0 $Y2=0
cc_140 N_A_M1005_g N_A_231_463#_c_262_n 0.00485524f $X=2.235 $Y=2.69 $X2=0 $Y2=0
cc_141 N_A_M1005_g N_A_231_463#_c_263_n 0.0222914f $X=2.235 $Y=2.69 $X2=0.24
+ $Y2=0
cc_142 N_A_M1005_g N_A_231_463#_c_267_n 0.0292059f $X=2.235 $Y=2.69 $X2=0 $Y2=0
cc_143 N_A_c_160_n N_A_231_463#_c_267_n 7.63737e-19 $X=2.945 $Y=1.725 $X2=0
+ $Y2=0
cc_144 N_A_M1002_g N_A_231_463#_c_267_n 0.0263501f $X=3.015 $Y=2.69 $X2=0 $Y2=0
cc_145 A N_A_231_463#_c_267_n 0.0226763f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_146 N_A_M1002_g N_VPWR_c_287_n 0.0355526f $X=3.015 $Y=2.69 $X2=0 $Y2=0
cc_147 A N_VPWR_c_287_n 0.00397758f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_148 N_A_M1002_g N_VPWR_c_290_n 0.0102412f $X=3.015 $Y=2.69 $X2=0 $Y2=0
cc_149 N_A_M1007_g N_A_217_207#_c_328_n 0.0268758f $X=2.165 $Y=1.335 $X2=0 $Y2=0
cc_150 N_A_M1007_g N_A_217_207#_c_329_n 0.00364144f $X=2.165 $Y=1.335 $X2=0
+ $Y2=0
cc_151 N_A_M1007_g N_A_217_207#_c_330_n 0.0115658f $X=2.165 $Y=1.335 $X2=0 $Y2=0
cc_152 N_A_M1003_g N_A_217_207#_c_330_n 0.0117354f $X=2.945 $Y=1.335 $X2=0 $Y2=0
cc_153 N_A_M1003_g N_VGND_c_354_n 0.0189566f $X=2.945 $Y=1.335 $X2=0 $Y2=0
cc_154 N_A_M1003_g N_VGND_c_356_n 0.0112668f $X=2.945 $Y=1.335 $X2=0.24 $Y2=0
cc_155 N_A_78_463#_c_204_n N_A_64_207#_c_232_n 0.0559351f $X=0.515 $Y=2.46 $X2=0
+ $Y2=0
cc_156 N_A_78_463#_c_199_n N_A_64_207#_c_232_n 0.00655667f $X=0.79 $Y=2.165
+ $X2=0 $Y2=0
cc_157 N_A_78_463#_c_205_n N_A_64_207#_c_232_n 0.0133946f $X=0.79 $Y=2.25 $X2=0
+ $Y2=0
cc_158 N_A_78_463#_c_204_n N_A_64_207#_c_233_n 0.0074717f $X=0.515 $Y=2.46 $X2=0
+ $Y2=0
cc_159 N_A_78_463#_c_199_n N_A_64_207#_c_230_n 0.0127878f $X=0.79 $Y=2.165
+ $X2=0.24 $Y2=0
cc_160 N_A_78_463#_c_205_n N_A_64_207#_c_230_n 0.00696349f $X=0.79 $Y=2.25
+ $X2=0.24 $Y2=0
cc_161 N_A_78_463#_c_199_n N_A_64_207#_c_231_n 0.0373159f $X=0.79 $Y=2.165 $X2=0
+ $Y2=0
cc_162 N_A_78_463#_c_204_n N_A_231_463#_c_262_n 0.0111595f $X=0.515 $Y=2.46
+ $X2=0 $Y2=0
cc_163 N_A_78_463#_c_205_n N_A_231_463#_c_262_n 0.00140122f $X=0.79 $Y=2.25
+ $X2=0 $Y2=0
cc_164 N_A_78_463#_c_204_n N_VPWR_c_290_n 0.00699215f $X=0.515 $Y=2.46 $X2=0
+ $Y2=0
cc_165 N_A_78_463#_c_202_n N_A_217_207#_c_328_n 0.0424266f $X=1.845 $Y=0.68
+ $X2=0 $Y2=0
cc_166 N_A_78_463#_c_199_n N_A_217_207#_c_329_n 0.0290289f $X=0.79 $Y=2.165
+ $X2=0 $Y2=0
cc_167 N_A_78_463#_c_202_n N_A_217_207#_c_329_n 0.0242676f $X=1.845 $Y=0.68
+ $X2=0 $Y2=0
cc_168 N_A_78_463#_X8_noxref_D1 N_VGND_c_356_n 0.00782386f $X=1.72 $Y=0.535
+ $X2=0.24 $Y2=0
cc_169 N_A_78_463#_c_200_n N_VGND_c_356_n 0.0109822f $X=0.875 $Y=0.682 $X2=0.24
+ $Y2=0
cc_170 N_A_78_463#_c_202_n N_VGND_c_356_n 0.0478825f $X=1.845 $Y=0.68 $X2=0.24
+ $Y2=0
cc_171 N_A_64_207#_X9_noxref_D0 N_VPWR_c_290_n 0.0274476f $X=0.78 $Y=3.425 $X2=0
+ $Y2=0
cc_172 N_A_64_207#_c_232_n N_VPWR_c_290_n 0.0121791f $X=0.17 $Y=3.485 $X2=0
+ $Y2=0
cc_173 N_A_64_207#_c_233_n N_VPWR_c_290_n 0.0214088f $X=0.74 $Y=3.57 $X2=0 $Y2=0
cc_174 N_A_64_207#_c_236_n N_VPWR_c_290_n 0.0090597f $X=0.255 $Y=3.57 $X2=0
+ $Y2=0
cc_175 N_A_64_207#_c_240_n N_VPWR_c_290_n 0.0306796f $X=0.905 $Y=3.57 $X2=0
+ $Y2=0
cc_176 N_A_64_207#_c_231_n N_VGND_c_356_n 0.0107361f $X=0.445 $Y=1.255 $X2=0.24
+ $Y2=0
cc_177 N_A_231_463#_c_263_n N_VPWR_c_287_n 0.00815017f $X=2.46 $Y=3.32 $X2=0.24
+ $Y2=4.07
cc_178 N_A_231_463#_c_267_n N_VPWR_c_287_n 0.0337481f $X=2.625 $Y=2.45 $X2=0.24
+ $Y2=4.07
cc_179 N_A_231_463#_c_263_n N_VPWR_c_290_n 0.0563871f $X=2.46 $Y=3.32 $X2=5.04
+ $Y2=4.07
cc_180 N_A_231_463#_c_265_n N_VPWR_c_290_n 0.0116935f $X=1.46 $Y=3.32 $X2=5.04
+ $Y2=4.07
cc_181 N_VPWR_c_287_n N_X_c_314_n 0.0681753f $X=3.31 $Y=3.56 $X2=2.64 $Y2=4.07
cc_182 N_VPWR_c_290_n N_X_c_314_n 0.0419719f $X=4.39 $Y=3.56 $X2=2.64 $Y2=4.07
cc_183 N_X_c_314_n N_VGND_c_354_n 0.0463675f $X=5.005 $Y=0.68 $X2=0 $Y2=0
cc_184 N_X_c_314_n N_VGND_c_356_n 0.0324928f $X=5.005 $Y=0.68 $X2=0.24 $Y2=0
cc_185 N_A_217_207#_c_330_n N_VGND_c_354_n 0.0125386f $X=2.555 $Y=1.06 $X2=0
+ $Y2=0
cc_186 N_A_217_207#_c_328_n N_VGND_c_356_n 0.0190504f $X=2.39 $Y=1.06 $X2=0.24
+ $Y2=0
cc_187 N_A_217_207#_c_329_n N_VGND_c_356_n 0.00177956f $X=1.225 $Y=1.06 $X2=0.24
+ $Y2=0
cc_188 N_A_217_207#_c_330_n N_VGND_c_356_n 0.0147915f $X=2.555 $Y=1.06 $X2=0.24
+ $Y2=0
