* File: sky130_fd_sc_hvl__dlclkp_1.pex.spice
* Created: Wed Sep  2 09:05:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__DLCLKP_1%VNB 5 7 17 24
c81 5 0 6.67964e-20 $X=-0.33 $Y=-0.265
r82 11 24 2.46376 $w=2.3e-07 $l=3.84e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r83 7 17 3.0797 $w=2.3e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=9.84
+ $Y2=0
r84 7 24 0.61594 $w=2.3e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.08
+ $Y2=0
r85 5 17 0.885714 $w=1.7e-07 $l=1.785e-06 $layer=mcon $count=10 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r86 5 11 0.885714 $w=1.7e-07 $l=1.785e-06 $layer=mcon $count=10 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__DLCLKP_1%VPB 4 6 14 15 21
r94 14 15 0.885714 $w=1.7e-07 $l=1.785e-06 $layer=mcon $count=10 $X=9.84 $Y=4.07
+ $X2=9.84 $Y2=4.07
r95 10 21 2.46376 $w=2.3e-07 $l=3.84e-06 $layer=MET1_cond $X=0.24 $Y=4.07
+ $X2=4.08 $Y2=4.07
r96 9 14 626.31 $w=1.68e-07 $l=9.6e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=9.84
+ $Y2=4.07
r97 9 10 0.885714 $w=1.7e-07 $l=1.785e-06 $layer=mcon $count=10 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r98 6 15 3.0797 $w=2.3e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=4.07 $X2=9.84
+ $Y2=4.07
r99 6 21 0.61594 $w=2.3e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=4.07 $X2=4.08
+ $Y2=4.07
r100 4 14 17.3333 $w=1.7e-07 $l=9.88241e-06 $layer=licon1_NTAP_notbjt $count=10
+ $X=0 $Y=3.985 $X2=9.84 $Y2=4.07
r101 4 9 17.3333 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=10
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__DLCLKP_1%GATE 1 2 6 10 12
r16 9 12 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=0.695 $Y=1.55
+ $X2=0.695 $Y2=2.6
r17 9 10 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.775
+ $Y=1.55 $X2=0.775 $Y2=1.55
r18 6 9 58.3182 $w=5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.695 $Y=1.005
+ $X2=0.695 $Y2=1.55
r19 1 2 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.775 $Y=1.665
+ $X2=0.775 $Y2=2.035
r20 1 10 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.775 $Y=1.665
+ $X2=0.775 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_HVL__DLCLKP_1%A_231_71# 1 2 9 12 14 17 19 22 25 28 32 37
+ 38 40 41 43 44 45 47 51 55
c114 19 0 4.52609e-21 $X=2.64 $Y=0.45
c115 12 0 1.75473e-19 $X=4.885 $Y=2.495
r116 41 57 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.84 $Y=3.13
+ $X2=4.84 $Y2=2.965
r117 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.01
+ $Y=3.13 $X2=5.01 $Y2=3.13
r118 38 40 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=4.07 $Y=3.11
+ $X2=5.01 $Y2=3.11
r119 35 38 6.81649 $w=2.1e-07 $l=1.48492e-07 $layer=LI1_cond $X=3.965 $Y=3.005
+ $X2=4.07 $Y2=3.11
r120 35 37 30.368 $w=2.08e-07 $l=5.75e-07 $layer=LI1_cond $X=3.965 $Y=3.005
+ $X2=3.965 $Y2=2.43
r121 34 45 3.98977 $w=2.3e-07 $l=9.44722e-08 $layer=LI1_cond $X=3.965 $Y=1.295
+ $X2=3.945 $Y2=1.21
r122 34 37 59.9437 $w=2.08e-07 $l=1.135e-06 $layer=LI1_cond $X=3.965 $Y=1.295
+ $X2=3.965 $Y2=2.43
r123 30 45 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.945 $Y=1.125
+ $X2=3.945 $Y2=1.21
r124 30 32 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.945 $Y=1.125
+ $X2=3.945 $Y2=0.87
r125 29 44 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.97 $Y=1.21
+ $X2=2.805 $Y2=1.21
r126 28 45 2.45049 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.82 $Y=1.21
+ $X2=3.945 $Y2=1.21
r127 28 29 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=3.82 $Y=1.21
+ $X2=2.97 $Y2=1.21
r128 26 51 128.407 $w=5e-07 $l=1.2e-06 $layer=POLY_cond $X=2.775 $Y=1.46
+ $X2=2.775 $Y2=2.66
r129 26 47 63.1335 $w=5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.775 $Y=1.46
+ $X2=2.775 $Y2=0.87
r130 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.805
+ $Y=1.46 $X2=2.805 $Y2=1.46
r131 23 44 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.805 $Y=1.295
+ $X2=2.805 $Y2=1.21
r132 23 25 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=1.295
+ $X2=2.805 $Y2=1.46
r133 22 44 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.725 $Y=1.125
+ $X2=2.805 $Y2=1.21
r134 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.725 $Y=0.535
+ $X2=2.725 $Y2=1.125
r135 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.64 $Y=0.45
+ $X2=2.725 $Y2=0.535
r136 19 43 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.64 $Y=0.45
+ $X2=1.865 $Y2=0.45
r137 17 55 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=0.52
+ $X2=1.49 $Y2=0.685
r138 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.66
+ $Y=0.52 $X2=1.66 $Y2=0.52
r139 14 43 7.98337 $w=3.03e-07 $l=1.52e-07 $layer=LI1_cond $X=1.713 $Y=0.517
+ $X2=1.865 $Y2=0.517
r140 14 16 2.00261 $w=3.03e-07 $l=5.3e-08 $layer=LI1_cond $X=1.713 $Y=0.517
+ $X2=1.66 $Y2=0.517
r141 12 57 50.2928 $w=5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.885 $Y=2.495
+ $X2=4.885 $Y2=2.965
r142 9 55 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.445 $Y=1.005
+ $X2=1.445 $Y2=0.685
r143 2 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.805
+ $Y=2.285 $X2=3.945 $Y2=2.43
r144 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.805
+ $Y=0.66 $X2=3.945 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_HVL__DLCLKP_1%A_239_419# 1 2 9 13 15 18 21 25 26 29 30
+ 31 34 35 37 39 42 44 45 48
c122 45 0 2.11044e-19 $X=5.14 $Y=1.78
c123 37 0 1.1081e-19 $X=5.43 $Y=3.385
c124 13 0 2.1354e-20 $X=4.885 $Y=1.005
r125 46 48 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.22 $Y=2.51
+ $X2=5.43 $Y2=2.51
r126 45 54 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.97 $Y=1.78
+ $X2=4.97 $Y2=1.615
r127 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.14
+ $Y=1.78 $X2=5.14 $Y2=1.78
r128 39 41 10.2694 $w=2.48e-07 $l=2.1e-07 $layer=LI1_cond $X=2.345 $Y=0.87
+ $X2=2.345 $Y2=1.08
r129 36 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=2.595
+ $X2=5.43 $Y2=2.51
r130 36 37 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=5.43 $Y=2.595
+ $X2=5.43 $Y2=3.385
r131 35 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.22 $Y=2.425
+ $X2=5.22 $Y2=2.51
r132 34 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.22 $Y=1.945
+ $X2=5.22 $Y2=1.78
r133 34 35 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=5.22 $Y=1.945
+ $X2=5.22 $Y2=2.425
r134 30 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.345 $Y=3.47
+ $X2=5.43 $Y2=3.385
r135 30 31 107.973 $w=1.68e-07 $l=1.655e-06 $layer=LI1_cond $X=5.345 $Y=3.47
+ $X2=3.69 $Y2=3.47
r136 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.605 $Y=3.385
+ $X2=3.69 $Y2=3.47
r137 28 29 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=3.605 $Y=2.315
+ $X2=3.605 $Y2=3.385
r138 27 42 2.06925 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.495 $Y=2.23
+ $X2=2.385 $Y2=2.23
r139 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.52 $Y=2.23
+ $X2=3.605 $Y2=2.315
r140 26 27 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=3.52 $Y=2.23
+ $X2=2.495 $Y2=2.23
r141 23 25 38.5021 $w=2.18e-07 $l=7.35e-07 $layer=LI1_cond $X=2.385 $Y=3.165
+ $X2=2.385 $Y2=2.43
r142 22 42 4.36305 $w=2.07e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=2.315
+ $X2=2.385 $Y2=2.23
r143 22 25 6.02413 $w=2.18e-07 $l=1.15e-07 $layer=LI1_cond $X=2.385 $Y=2.315
+ $X2=2.385 $Y2=2.43
r144 21 42 4.36305 $w=2.07e-07 $l=9.12688e-08 $layer=LI1_cond $X=2.372 $Y=2.145
+ $X2=2.385 $Y2=2.23
r145 21 41 60.5734 $w=1.93e-07 $l=1.065e-06 $layer=LI1_cond $X=2.372 $Y=2.145
+ $X2=2.372 $Y2=1.08
r146 18 51 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.53 $Y=3.3
+ $X2=1.53 $Y2=3.135
r147 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.7 $Y=3.3
+ $X2=1.7 $Y2=3.3
r148 15 23 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=2.275 $Y=3.275
+ $X2=2.385 $Y2=3.165
r149 15 17 30.1207 $w=2.18e-07 $l=5.75e-07 $layer=LI1_cond $X=2.275 $Y=3.275
+ $X2=1.7 $Y2=3.275
r150 13 54 65.2736 $w=5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.885 $Y=1.005
+ $X2=4.885 $Y2=1.615
r151 9 51 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.445 $Y=2.6
+ $X2=1.445 $Y2=3.135
r152 2 25 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.26
+ $Y=2.285 $X2=2.385 $Y2=2.43
r153 1 39 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.26
+ $Y=0.66 $X2=2.385 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_HVL__DLCLKP_1%A_1069_133# 1 2 9 14 19 20 22 23 26 30 32
+ 34 37 44 48
c78 23 0 1.53715e-19 $X=5.845 $Y=1.98
c79 9 0 1.06584e-19 $X=5.595 $Y=1.005
r80 38 48 111.286 $w=5e-07 $l=1.04e-06 $layer=POLY_cond $X=7.705 $Y=1.55
+ $X2=7.705 $Y2=2.59
r81 38 44 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.705 $Y=1.55
+ $X2=7.705 $Y2=1.065
r82 37 40 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.62 $Y=1.55
+ $X2=7.62 $Y2=1.72
r83 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.62
+ $Y=1.55 $X2=7.62 $Y2=1.55
r84 34 35 11.0976 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.795 $Y=1.72
+ $X2=6.795 $Y2=1.98
r85 33 34 2.2115 $w=2.1e-07 $l=1.35e-07 $layer=LI1_cond $X=6.93 $Y=1.72
+ $X2=6.795 $Y2=1.72
r86 32 40 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=7.455 $Y=1.72
+ $X2=7.62 $Y2=1.72
r87 32 33 27.7273 $w=2.08e-07 $l=5.25e-07 $layer=LI1_cond $X=7.455 $Y=1.72
+ $X2=6.93 $Y2=1.72
r88 28 35 4.48172 $w=2.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.795 $Y=2.085
+ $X2=6.795 $Y2=1.98
r89 28 30 17.5001 $w=2.68e-07 $l=4.1e-07 $layer=LI1_cond $X=6.795 $Y=2.085
+ $X2=6.795 $Y2=2.495
r90 24 34 4.48172 $w=2.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.795 $Y=1.615
+ $X2=6.795 $Y2=1.72
r91 24 26 26.0367 $w=2.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.795 $Y=1.615
+ $X2=6.795 $Y2=1.005
r92 22 35 2.2115 $w=2.1e-07 $l=1.35e-07 $layer=LI1_cond $X=6.66 $Y=1.98
+ $X2=6.795 $Y2=1.98
r93 22 23 43.0433 $w=2.08e-07 $l=8.15e-07 $layer=LI1_cond $X=6.66 $Y=1.98
+ $X2=5.845 $Y2=1.98
r94 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.68
+ $Y=1.62 $X2=5.68 $Y2=1.62
r95 17 23 7.26367 $w=2.1e-07 $l=2.11069e-07 $layer=LI1_cond $X=5.68 $Y=1.875
+ $X2=5.845 $Y2=1.98
r96 17 19 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.68 $Y=1.875
+ $X2=5.68 $Y2=1.62
r97 15 20 93.5508 $w=3.3e-07 $l=5.35e-07 $layer=POLY_cond $X=5.68 $Y=2.155
+ $X2=5.68 $Y2=1.62
r98 14 15 42.5715 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.595 $Y=2.495
+ $X2=5.595 $Y2=2.155
r99 11 20 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=5.68 $Y=1.345
+ $X2=5.68 $Y2=1.62
r100 9 11 42.5715 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.595 $Y=1.005
+ $X2=5.595 $Y2=1.345
r101 2 30 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.625
+ $Y=2.285 $X2=6.765 $Y2=2.495
r102 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.625
+ $Y=0.795 $X2=6.765 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HVL__DLCLKP_1%A_303_311# 1 2 3 4 14 15 16 17 18 19 22 26
+ 31 34 41 48 50 52 53 56 64 69 71 74
c139 71 0 1.1081e-19 $X=6.375 $Y=1.005
c140 52 0 1.24125e-19 $X=4.495 $Y=2.495
c141 48 0 2.1354e-20 $X=4.517 $Y=0.395
c142 34 0 1.06584e-19 $X=6.125 $Y=1.28
r143 69 71 34.2419 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.375 $Y=0.685
+ $X2=6.375 $Y2=1.005
r144 65 69 52.6077 $w=3.39e-07 $l=3.7e-07 $layer=POLY_cond $X=6.745 $Y=0.495
+ $X2=6.375 $Y2=0.495
r145 64 65 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.745
+ $Y=0.52 $X2=6.745 $Y2=0.52
r146 61 64 12.4391 $w=3.13e-07 $l=3.4e-07 $layer=LI1_cond $X=6.405 $Y=0.512
+ $X2=6.745 $Y2=0.512
r147 59 74 107.541 $w=5e-07 $l=1.005e-06 $layer=POLY_cond $X=6.375 $Y=1.49
+ $X2=6.375 $Y2=2.495
r148 59 71 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.375 $Y=1.49
+ $X2=6.375 $Y2=1.005
r149 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.29
+ $Y=1.49 $X2=6.29 $Y2=1.49
r150 52 53 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=4.517 $Y=2.495
+ $X2=4.517 $Y2=2.33
r151 45 48 10.5778 $w=2.78e-07 $l=2.57e-07 $layer=LI1_cond $X=4.26 $Y=0.395
+ $X2=4.517 $Y2=0.395
r152 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.26
+ $Y=0.41 $X2=4.26 $Y2=0.41
r153 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.02
+ $Y=1.72 $X2=2.02 $Y2=1.72
r154 38 41 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.835 $Y=1.72
+ $X2=2.02 $Y2=1.72
r155 36 61 4.34843 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=6.405 $Y=0.67
+ $X2=6.405 $Y2=0.512
r156 36 56 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=6.405 $Y=0.67
+ $X2=6.405 $Y2=1.195
r157 35 50 2.40986 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=4.66 $Y=1.28
+ $X2=4.517 $Y2=1.28
r158 34 58 6.63049 $w=3.63e-07 $l=2.1e-07 $layer=LI1_cond $X=6.307 $Y=1.28
+ $X2=6.307 $Y2=1.49
r159 34 56 5.9984 $w=3.63e-07 $l=8.5e-08 $layer=LI1_cond $X=6.307 $Y=1.28
+ $X2=6.307 $Y2=1.195
r160 34 35 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=6.125 $Y=1.28
+ $X2=4.66 $Y2=1.28
r161 32 50 4.02809 $w=2.27e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.46 $Y=1.365
+ $X2=4.517 $Y2=1.28
r162 32 53 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=4.46 $Y=1.365
+ $X2=4.46 $Y2=2.33
r163 29 50 4.02809 $w=2.27e-07 $l=8.5e-08 $layer=LI1_cond $X=4.517 $Y=1.195
+ $X2=4.517 $Y2=1.28
r164 29 31 7.68295 $w=2.83e-07 $l=1.9e-07 $layer=LI1_cond $X=4.517 $Y=1.195
+ $X2=4.517 $Y2=1.005
r165 28 48 0.630043 $w=2.85e-07 $l=1.4e-07 $layer=LI1_cond $X=4.517 $Y=0.535
+ $X2=4.517 $Y2=0.395
r166 28 31 19.0052 $w=2.83e-07 $l=4.7e-07 $layer=LI1_cond $X=4.517 $Y=0.535
+ $X2=4.517 $Y2=1.005
r167 24 38 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=1.885
+ $X2=1.835 $Y2=1.72
r168 24 26 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.835 $Y=1.885
+ $X2=1.835 $Y2=2.37
r169 20 38 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=1.555
+ $X2=1.835 $Y2=1.72
r170 20 22 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=1.835 $Y=1.555
+ $X2=1.835 $Y2=1.005
r171 19 42 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.035 $Y=1.72
+ $X2=2.02 $Y2=1.72
r172 18 46 38.9663 $w=3.64e-07 $l=1.68953e-07 $layer=POLY_cond $X=4.425 $Y=0.38
+ $X2=4.26 $Y2=0.372
r173 17 69 50.756 $w=3.39e-07 $l=3.02076e-07 $layer=POLY_cond $X=6.125 $Y=0.38
+ $X2=6.375 $Y2=0.495
r174 17 18 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=6.125 $Y=0.38
+ $X2=4.425 $Y2=0.38
r175 15 46 38.9663 $w=3.64e-07 $l=2.19499e-07 $layer=POLY_cond $X=4.095 $Y=0.245
+ $X2=4.26 $Y2=0.372
r176 15 16 979.383 $w=1.5e-07 $l=1.91e-06 $layer=POLY_cond $X=4.095 $Y=0.245
+ $X2=2.185 $Y2=0.245
r177 14 19 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.11 $Y=1.555
+ $X2=2.035 $Y2=1.72
r178 13 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.11 $Y=0.32
+ $X2=2.185 $Y2=0.245
r179 13 14 633.266 $w=1.5e-07 $l=1.235e-06 $layer=POLY_cond $X=2.11 $Y=0.32
+ $X2=2.11 $Y2=1.555
r180 4 52 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=2.285 $X2=4.495 $Y2=2.495
r181 3 26 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=2.225 $X2=1.835 $Y2=2.37
r182 2 31 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=4.37
+ $Y=0.795 $X2=4.495 $Y2=1.005
r183 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.795 $X2=1.835 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HVL__DLCLKP_1%CLK 1 3 4 7 8 9 10 13 14 20 25 26 27 30 34
+ 37 44 48
c102 37 0 4.52609e-21 $X=3.555 $Y=0.87
c103 10 0 1.82094e-19 $X=8.235 $Y=3.38
c104 1 0 8.39567e-20 $X=3.555 $Y=2.21
r105 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.525
+ $Y=1.55 $X2=3.525 $Y2=1.55
r106 37 40 72.764 $w=5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.555 $Y=0.87
+ $X2=3.555 $Y2=1.55
r107 34 41 1.75894 $w=5.08e-07 $l=7.5e-08 $layer=LI1_cond $X=3.6 $Y=1.72
+ $X2=3.525 $Y2=1.72
r108 31 48 74.9041 $w=5e-07 $l=7e-07 $layer=POLY_cond $X=8.485 $Y=1.89 $X2=8.485
+ $Y2=2.59
r109 31 44 88.2799 $w=5e-07 $l=8.25e-07 $layer=POLY_cond $X=8.485 $Y=1.89
+ $X2=8.485 $Y2=1.065
r110 30 33 5.41921 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=8.515 $Y=1.89
+ $X2=8.515 $Y2=2.025
r111 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.515
+ $Y=1.89 $X2=8.515 $Y2=1.89
r112 27 33 50.7075 $w=2.48e-07 $l=1.1e-06 $layer=LI1_cond $X=8.475 $Y=3.125
+ $X2=8.475 $Y2=2.025
r113 25 27 6.36223 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=8.417 $Y=3.29
+ $X2=8.417 $Y2=3.125
r114 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.4
+ $Y=3.29 $X2=8.4 $Y2=3.29
r115 21 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.4 $Y=3.305
+ $X2=8.4 $Y2=3.29
r116 20 26 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=8.4 $Y=3.095
+ $X2=8.4 $Y2=3.29
r117 18 48 27.2865 $w=5e-07 $l=2.55e-07 $layer=POLY_cond $X=8.485 $Y=2.845
+ $X2=8.485 $Y2=2.59
r118 18 20 32.941 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.485 $Y=2.845
+ $X2=8.485 $Y2=3.095
r119 14 16 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=5.46 $Y=3.38 $X2=5.46
+ $Y2=3.58
r120 12 40 54.573 $w=5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.555 $Y=2.06
+ $X2=3.555 $Y2=1.55
r121 12 13 6.88608 $w=5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.555 $Y=2.06
+ $X2=3.555 $Y2=2.135
r122 11 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.535 $Y=3.38
+ $X2=5.46 $Y2=3.38
r123 10 21 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.235 $Y=3.38
+ $X2=8.4 $Y2=3.305
r124 10 11 1384.47 $w=1.5e-07 $l=2.7e-06 $layer=POLY_cond $X=8.235 $Y=3.38
+ $X2=5.535 $Y2=3.38
r125 8 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.385 $Y=3.58
+ $X2=5.46 $Y2=3.58
r126 8 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=5.385 $Y=3.58
+ $X2=4.295 $Y2=3.58
r127 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.22 $Y=3.505
+ $X2=4.295 $Y2=3.58
r128 6 7 664.032 $w=1.5e-07 $l=1.295e-06 $layer=POLY_cond $X=4.22 $Y=2.21
+ $X2=4.22 $Y2=3.505
r129 5 13 23.237 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.805 $Y=2.135
+ $X2=3.555 $Y2=2.135
r130 4 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.145 $Y=2.135
+ $X2=4.22 $Y2=2.21
r131 4 5 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.145 $Y=2.135
+ $X2=3.805 $Y2=2.135
r132 1 13 6.88608 $w=5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.555 $Y=2.21
+ $X2=3.555 $Y2=2.135
r133 1 3 43.38 $w=5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.555 $Y=2.21 $X2=3.555
+ $Y2=2.66
.ends

.subckt PM_SKY130_FD_SC_HVL__DLCLKP_1%A_1438_171# 1 2 9 12 14 19 22 26 28 29 30
+ 33
r59 29 34 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.28 $Y=1.56
+ $X2=9.28 $Y2=1.725
r60 29 33 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.28 $Y=1.56
+ $X2=9.28 $Y2=1.395
r61 28 30 19.9963 $w=3.38e-07 $l=5.05e-07 $layer=LI1_cond $X=9.45 $Y=1.555
+ $X2=8.945 $Y2=1.555
r62 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.45
+ $Y=1.56 $X2=9.45 $Y2=1.56
r63 25 26 2.36881 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=8.18 $Y=1.47
+ $X2=8.067 $Y2=1.47
r64 25 30 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=8.18 $Y=1.47
+ $X2=8.945 $Y2=1.47
r65 20 26 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=8.067 $Y=1.555
+ $X2=8.067 $Y2=1.47
r66 20 22 41.2318 $w=2.23e-07 $l=8.05e-07 $layer=LI1_cond $X=8.067 $Y=1.555
+ $X2=8.067 $Y2=2.36
r67 19 26 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=8.067 $Y=1.385
+ $X2=8.067 $Y2=1.47
r68 18 19 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=8.067 $Y=1.215
+ $X2=8.067 $Y2=1.385
r69 14 18 7.1387 $w=3.3e-07 $l=2.13787e-07 $layer=LI1_cond $X=7.955 $Y=1.05
+ $X2=8.067 $Y2=1.215
r70 14 16 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=7.955 $Y=1.05
+ $X2=7.315 $Y2=1.05
r71 12 34 132.687 $w=5e-07 $l=1.24e-06 $layer=POLY_cond $X=9.325 $Y=2.965
+ $X2=9.325 $Y2=1.725
r72 9 33 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.325 $Y=0.91 $X2=9.325
+ $Y2=1.395
r73 2 22 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.955
+ $Y=2.215 $X2=8.095 $Y2=2.36
r74 1 16 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=7.19
+ $Y=0.855 $X2=7.315 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_HVL__DLCLKP_1%VPWR 1 2 3 4 5 18 22 24 26 28 32 36 40 42
+ 44 45 46 48 67 71 72 78 80 81 89
c110 80 0 1.82094e-19 $X=9.36 $Y=3.56
c111 72 0 8.39567e-20 $X=3.165 $Y=3.63
c112 26 0 1.75473e-19 $X=5.985 $Y=2.495
r113 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.56
+ $X2=9.36 $Y2=3.56
r114 77 80 13.2375 $w=3.68e-07 $l=4.25e-07 $layer=LI1_cond $X=8.935 $Y=3.63
+ $X2=9.36 $Y2=3.63
r115 77 78 7.556 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.935 $Y=3.63
+ $X2=8.77 $Y2=3.63
r116 75 76 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.8 $Y=3.56 $X2=5.8
+ $Y2=3.56
r117 70 89 0.353193 $w=3.7e-07 $l=9.2e-07 $layer=MET1_cond $X=3.16 $Y=3.63
+ $X2=4.08 $Y2=3.63
r118 69 72 0.155736 $w=3.68e-07 $l=5e-09 $layer=LI1_cond $X=3.16 $Y=3.63
+ $X2=3.165 $Y2=3.63
r119 69 71 16.4502 $w=3.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.16 $Y=3.63
+ $X2=2.665 $Y2=3.63
r120 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.16 $Y=3.56
+ $X2=3.16 $Y2=3.56
r121 65 67 3.52417 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=0.945 $Y=3.63
+ $X2=1.025 $Y2=3.63
r122 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.945 $Y=3.685
+ $X2=0.945 $Y2=3.685
r123 63 81 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.64 $Y=3.63
+ $X2=9.36 $Y2=3.63
r124 62 78 7.20909 $w=1.98e-07 $l=1.3e-07 $layer=LI1_cond $X=8.64 $Y=3.715
+ $X2=8.77 $Y2=3.715
r125 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.64 $Y=3.7
+ $X2=8.64 $Y2=3.7
r126 59 63 0.399262 $w=3.7e-07 $l=1.04e-06 $layer=MET1_cond $X=7.6 $Y=3.63
+ $X2=8.64 $Y2=3.63
r127 59 76 0.69103 $w=3.7e-07 $l=1.8e-06 $layer=MET1_cond $X=7.6 $Y=3.63 $X2=5.8
+ $Y2=3.63
r128 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.6 $Y=3.56 $X2=7.6
+ $Y2=3.56
r129 56 70 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.44 $Y=3.63
+ $X2=3.16 $Y2=3.63
r130 56 66 0.573939 $w=3.7e-07 $l=1.495e-06 $layer=MET1_cond $X=2.44 $Y=3.63
+ $X2=0.945 $Y2=3.63
r131 55 71 9.97306 $w=2.58e-07 $l=2.25e-07 $layer=LI1_cond $X=2.44 $Y=3.685
+ $X2=2.665 $Y2=3.685
r132 55 67 62.7195 $w=2.58e-07 $l=1.415e-06 $layer=LI1_cond $X=2.44 $Y=3.685
+ $X2=1.025 $Y2=3.685
r133 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.44 $Y=3.685
+ $X2=2.44 $Y2=3.685
r134 51 66 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=0.585 $Y=3.63
+ $X2=0.945 $Y2=3.63
r135 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.585 $Y=3.56
+ $X2=0.585 $Y2=3.56
r136 48 65 3.27045 $w=3.68e-07 $l=1.05e-07 $layer=LI1_cond $X=0.84 $Y=3.63
+ $X2=0.945 $Y2=3.63
r137 48 50 7.94251 $w=3.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.84 $Y=3.63
+ $X2=0.585 $Y2=3.63
r138 46 76 0.291768 $w=3.7e-07 $l=7.6e-07 $layer=MET1_cond $X=5.04 $Y=3.63
+ $X2=5.8 $Y2=3.63
r139 46 89 0.368549 $w=3.7e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.63
+ $X2=4.08 $Y2=3.63
r140 45 62 31.8864 $w=1.98e-07 $l=5.75e-07 $layer=LI1_cond $X=8.065 $Y=3.715
+ $X2=8.64 $Y2=3.715
r141 44 58 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.88 $Y=3.63
+ $X2=7.6 $Y2=3.63
r142 44 45 8.17894 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=7.88 $Y=3.63
+ $X2=8.065 $Y2=3.63
r143 41 58 3.73765 $w=3.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.48 $Y=3.63
+ $X2=7.6 $Y2=3.63
r144 41 42 4.69202 $w=3.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.48 $Y=3.63
+ $X2=7.315 $Y2=3.63
r145 40 50 4.51633 $w=3.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.44 $Y=3.63
+ $X2=0.585 $Y2=3.63
r146 36 39 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=8.935 $Y=2.36
+ $X2=8.935 $Y2=3.23
r147 34 77 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=8.935 $Y=3.445
+ $X2=8.935 $Y2=3.63
r148 34 39 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=8.935 $Y=3.445
+ $X2=8.935 $Y2=3.23
r149 30 42 1.75761 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=7.315 $Y=3.445
+ $X2=7.315 $Y2=3.63
r150 30 32 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=7.315 $Y=3.445
+ $X2=7.315 $Y2=2.36
r151 29 75 3.28189 $w=3.7e-07 $l=2.33e-07 $layer=LI1_cond $X=6.15 $Y=3.63
+ $X2=5.917 $Y2=3.63
r152 28 42 4.69202 $w=3.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.15 $Y=3.63
+ $X2=7.315 $Y2=3.63
r153 28 29 31.1471 $w=3.68e-07 $l=1e-06 $layer=LI1_cond $X=7.15 $Y=3.63 $X2=6.15
+ $Y2=3.63
r154 24 75 3.56359 $w=3.3e-07 $l=2.16345e-07 $layer=LI1_cond $X=5.985 $Y=3.445
+ $X2=5.917 $Y2=3.63
r155 24 26 33.1764 $w=3.28e-07 $l=9.5e-07 $layer=LI1_cond $X=5.985 $Y=3.445
+ $X2=5.985 $Y2=2.495
r156 20 72 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=3.165 $Y=3.445
+ $X2=3.165 $Y2=3.63
r157 20 22 30.5572 $w=3.28e-07 $l=8.75e-07 $layer=LI1_cond $X=3.165 $Y=3.445
+ $X2=3.165 $Y2=2.57
r158 16 40 6.84548 $w=3.7e-07 $l=2.5446e-07 $layer=LI1_cond $X=0.275 $Y=3.445
+ $X2=0.44 $Y2=3.63
r159 16 18 37.5417 $w=3.28e-07 $l=1.075e-06 $layer=LI1_cond $X=0.275 $Y=3.445
+ $X2=0.275 $Y2=2.37
r160 5 39 300 $w=1.7e-07 $l=1.11051e-06 $layer=licon1_PDIFF $count=2 $X=8.735
+ $Y=2.215 $X2=8.935 $Y2=3.23
r161 5 36 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=8.735
+ $Y=2.215 $X2=8.935 $Y2=2.36
r162 4 32 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=7.19
+ $Y=2.215 $X2=7.315 $Y2=2.36
r163 3 26 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.845
+ $Y=2.285 $X2=5.985 $Y2=2.495
r164 2 22 300 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=2 $X=3.025
+ $Y=2.285 $X2=3.165 $Y2=2.57
r165 1 18 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.225 $X2=0.305 $Y2=2.37
.ends

.subckt PM_SKY130_FD_SC_HVL__DLCLKP_1%GCLK 1 2 9 11 12 13 22 38
r21 29 31 38.2043 $w=3.63e-07 $l=1.21e-06 $layer=LI1_cond $X=9.812 $Y=2.36
+ $X2=9.812 $Y2=3.57
r22 26 38 1.3261 $w=3.63e-07 $l=4.2e-08 $layer=LI1_cond $X=9.812 $Y=2.077
+ $X2=9.812 $Y2=2.035
r23 22 34 3.41465 $w=2.68e-07 $l=8e-08 $layer=LI1_cond $X=9.86 $Y=1.295 $X2=9.86
+ $Y2=1.215
r24 13 38 0.694623 $w=3.63e-07 $l=2.2e-08 $layer=LI1_cond $X=9.812 $Y=2.013
+ $X2=9.812 $Y2=2.035
r25 13 36 4.52998 $w=3.63e-07 $l=1.18e-07 $layer=LI1_cond $X=9.812 $Y=2.013
+ $X2=9.812 $Y2=1.895
r26 13 29 8.27233 $w=3.63e-07 $l=2.62e-07 $layer=LI1_cond $X=9.812 $Y=2.098
+ $X2=9.812 $Y2=2.36
r27 13 26 0.663049 $w=3.63e-07 $l=2.1e-08 $layer=LI1_cond $X=9.812 $Y=2.098
+ $X2=9.812 $Y2=2.077
r28 12 36 9.81711 $w=2.68e-07 $l=2.3e-07 $layer=LI1_cond $X=9.86 $Y=1.665
+ $X2=9.86 $Y2=1.895
r29 11 34 0.898996 $w=3.63e-07 $l=3e-09 $layer=LI1_cond $X=9.812 $Y=1.212
+ $X2=9.812 $Y2=1.215
r30 11 12 15.7074 $w=2.68e-07 $l=3.68e-07 $layer=LI1_cond $X=9.86 $Y=1.297
+ $X2=9.86 $Y2=1.665
r31 11 22 0.0853661 $w=2.68e-07 $l=2e-09 $layer=LI1_cond $X=9.86 $Y=1.297
+ $X2=9.86 $Y2=1.295
r32 7 11 5.65171 $w=3.63e-07 $l=1.79e-07 $layer=LI1_cond $X=9.812 $Y=1.033
+ $X2=9.812 $Y2=1.212
r33 7 9 11.1455 $w=3.63e-07 $l=3.53e-07 $layer=LI1_cond $X=9.812 $Y=1.033
+ $X2=9.812 $Y2=0.68
r34 2 31 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=9.575
+ $Y=2.215 $X2=9.715 $Y2=3.57
r35 2 29 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=9.575
+ $Y=2.215 $X2=9.715 $Y2=2.36
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.575
+ $Y=0.535 $X2=9.715 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__DLCLKP_1%VGND 1 2 3 4 15 17 19 23 27 28 31 34 39 47
+ 57 58 65
r94 57 58 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=9.345 $Y=0.51
+ $X2=9.345 $Y2=0.51
r95 55 57 12.7703 $w=3.68e-07 $l=4.1e-07 $layer=LI1_cond $X=8.935 $Y=0.44
+ $X2=9.345 $Y2=0.44
r96 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.035 $Y=0.51
+ $X2=6.035 $Y2=0.51
r97 51 65 0.107494 $w=3.7e-07 $l=2.8e-07 $layer=MET1_cond $X=3.8 $Y=0.44
+ $X2=4.08 $Y2=0.44
r98 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.8 $Y=0.44 $X2=3.8
+ $Y2=0.44
r99 48 51 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=3.44 $Y=0.44
+ $X2=3.8 $Y2=0.44
r100 47 50 9.42489 $w=4.66e-07 $l=4.34741e-07 $layer=LI1_cond $X=3.44 $Y=0.605
+ $X2=3.8 $Y2=0.44
r101 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.44 $Y=0.51
+ $X2=3.44 $Y2=0.51
r102 45 47 7.19957 $w=4.66e-07 $l=2.75e-07 $layer=LI1_cond $X=3.165 $Y=0.605
+ $X2=3.44 $Y2=0.605
r103 42 58 0.829236 $w=3.7e-07 $l=2.16e-06 $layer=MET1_cond $X=7.185 $Y=0.44
+ $X2=9.345 $Y2=0.44
r104 42 54 0.441491 $w=3.7e-07 $l=1.15e-06 $layer=MET1_cond $X=7.185 $Y=0.44
+ $X2=6.035 $Y2=0.44
r105 41 42 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.185 $Y=0.44
+ $X2=7.185 $Y2=0.44
r106 39 55 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.77 $Y=0.44
+ $X2=8.935 $Y2=0.44
r107 39 41 49.3682 $w=3.68e-07 $l=1.585e-06 $layer=LI1_cond $X=8.77 $Y=0.44
+ $X2=7.185 $Y2=0.44
r108 34 53 3.22716 $w=3.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=0.44
+ $X2=5.985 $Y2=0.44
r109 34 36 26.9422 $w=3.68e-07 $l=8.65e-07 $layer=LI1_cond $X=5.82 $Y=0.44
+ $X2=4.955 $Y2=0.44
r110 32 48 1.08261 $w=3.7e-07 $l=2.82e-06 $layer=MET1_cond $X=0.62 $Y=0.44
+ $X2=3.44 $Y2=0.44
r111 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.62 $Y=0.51
+ $X2=0.62 $Y2=0.51
r112 28 54 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=4.955 $Y=0.44
+ $X2=6.035 $Y2=0.44
r113 28 65 0.335917 $w=3.7e-07 $l=8.75e-07 $layer=MET1_cond $X=4.955 $Y=0.44
+ $X2=4.08 $Y2=0.44
r114 28 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.955 $Y=0.44
+ $X2=4.955 $Y2=0.44
r115 27 31 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=0.47 $Y=0.495
+ $X2=0.62 $Y2=0.495
r116 23 25 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=8.935 $Y=0.68
+ $X2=8.935 $Y2=1.09
r117 21 55 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=8.935 $Y=0.625
+ $X2=8.935 $Y2=0.44
r118 21 23 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=8.935 $Y=0.625
+ $X2=8.935 $Y2=0.68
r119 17 53 3.61833 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=5.985 $Y=0.625
+ $X2=5.985 $Y2=0.44
r120 17 19 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.985 $Y=0.625
+ $X2=5.985 $Y2=0.94
r121 13 27 6.94204 $w=2.6e-07 $l=2.20624e-07 $layer=LI1_cond $X=0.305 $Y=0.625
+ $X2=0.47 $Y2=0.495
r122 13 15 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.305 $Y=0.625
+ $X2=0.305 $Y2=1.005
r123 4 25 182 $w=1.7e-07 $l=3.19726e-07 $layer=licon1_NDIFF $count=1 $X=8.735
+ $Y=0.855 $X2=8.935 $Y2=1.09
r124 4 23 182 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_NDIFF $count=1 $X=8.735
+ $Y=0.855 $X2=8.935 $Y2=0.68
r125 3 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.845
+ $Y=0.795 $X2=5.985 $Y2=0.94
r126 2 45 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.66 $X2=3.165 $Y2=0.87
r127 1 15 182 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.795 $X2=0.305 $Y2=1.005
.ends

