# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  24.96000 BY  8.140000 ;
  SYMMETRY X Y R90 ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 21.070000 5.975000 21.400000 6.455000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.750000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.315000 5.545000 14.985000 5.875000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  2.180000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.645000 1.280000 1.920000 ;
        RECT 1.060000 1.920000 2.840000 2.140000 ;
        RECT 1.060000 2.140000 1.280000 5.115000 ;
        RECT 2.620000 0.645000 2.840000 1.920000 ;
        RECT 2.620000 2.140000 2.840000 5.115000 ;
    END
  END X
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 17.785000 4.435000 21.400000 4.605000 ;
        RECT 17.785000 4.605000 18.035000 5.465000 ;
        RECT 17.795000 3.905000 20.420000 4.235000 ;
        RECT 17.815000 2.335000 18.065000 3.535000 ;
        RECT 17.815000 3.535000 20.420000 3.705000 ;
        RECT 18.765000 4.605000 18.935000 5.465000 ;
        RECT 18.795000 2.675000 18.965000 3.535000 ;
        RECT 19.665000 3.705000 20.420000 3.905000 ;
        RECT 19.665000 4.235000 20.420000 4.435000 ;
        RECT 19.665000 4.605000 20.420000 5.805000 ;
        RECT 19.695000 2.675000 19.945000 3.020000 ;
        RECT 19.695000 3.020000 20.420000 3.535000 ;
        RECT 20.170000 5.805000 20.420000 5.935000 ;
        RECT 21.070000 4.605000 21.400000 5.805000 ;
    END
    PORT
      LAYER mcon ;
        RECT 19.800000 3.070000 19.970000 3.240000 ;
        RECT 20.160000 3.070000 20.330000 3.240000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 24.890000 3.305000 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  1.060000 6.195000  1.280000 6.850000 ;
        RECT  1.060000 6.850000  1.810000 7.180000 ;
        RECT  1.060000 7.180000  1.280000 7.570000 ;
        RECT  1.060000 7.570000 14.885000 7.800000 ;
        RECT  2.360000 6.195000  2.585000 7.205000 ;
        RECT  2.360000 7.205000  2.580000 7.570000 ;
        RECT  4.750000 6.195000  4.970000 7.570000 ;
        RECT  7.110000 6.195000  7.330000 7.570000 ;
        RECT  9.470000 6.195000  9.690000 7.570000 ;
        RECT 11.830000 6.195000 12.050000 7.570000 ;
        RECT 13.335000 6.195000 13.555000 7.570000 ;
        RECT 14.665000 6.195000 14.885000 7.570000 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.835000 0.255000 2.425000 0.485000 ;
        RECT 1.835000 0.485000 2.065000 1.655000 ;
    END
    PORT
      LAYER li1 ;
        RECT 17.780000 0.395000 19.950000 0.625000 ;
        RECT 17.780000 0.625000 18.110000 1.175000 ;
        RECT 18.710000 0.625000 19.040000 1.225000 ;
        RECT 19.620000 0.625000 19.950000 1.225000 ;
    END
    PORT
      LAYER li1 ;
        RECT 17.780000 6.915000 18.110000 7.515000 ;
        RECT 17.780000 7.515000 21.375000 7.745000 ;
        RECT 18.690000 6.915000 19.020000 7.515000 ;
        RECT 19.620000 6.625000 19.950000 7.515000 ;
        RECT 20.185000 6.625000 20.435000 7.515000 ;
        RECT 21.125000 6.625000 21.375000 7.515000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.035000 0.255000 3.625000 0.485000 ;
        RECT 3.395000 0.485000 3.625000 1.655000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.545000 0.255000 5.135000 0.485000 ;
        RECT 4.725000 0.485000 4.955000 1.655000 ;
    END
    PORT
      LAYER mcon ;
        RECT  1.115000 7.600000  1.285000 7.770000 ;
        RECT  1.595000 7.600000  1.765000 7.770000 ;
        RECT  1.865000 0.285000  2.035000 0.455000 ;
        RECT  2.075000 7.600000  2.245000 7.770000 ;
        RECT  2.225000 0.285000  2.395000 0.455000 ;
        RECT  2.555000 7.600000  2.725000 7.770000 ;
        RECT  3.035000 7.600000  3.205000 7.770000 ;
        RECT  3.065000 0.285000  3.235000 0.455000 ;
        RECT  3.425000 0.285000  3.595000 0.455000 ;
        RECT  3.515000 7.600000  3.685000 7.770000 ;
        RECT  3.995000 7.600000  4.165000 7.770000 ;
        RECT  4.475000 7.600000  4.645000 7.770000 ;
        RECT  4.575000 0.285000  4.745000 0.455000 ;
        RECT  4.935000 0.285000  5.105000 0.455000 ;
        RECT  4.955000 7.600000  5.125000 7.770000 ;
        RECT  5.435000 7.600000  5.605000 7.770000 ;
        RECT  5.915000 7.600000  6.085000 7.770000 ;
        RECT  6.395000 7.600000  6.565000 7.770000 ;
        RECT  6.875000 7.600000  7.045000 7.770000 ;
        RECT  7.355000 7.600000  7.525000 7.770000 ;
        RECT  7.835000 7.600000  8.005000 7.770000 ;
        RECT  8.315000 7.600000  8.485000 7.770000 ;
        RECT  8.795000 7.600000  8.965000 7.770000 ;
        RECT  9.275000 7.600000  9.445000 7.770000 ;
        RECT  9.755000 7.600000  9.925000 7.770000 ;
        RECT 10.235000 7.600000 10.405000 7.770000 ;
        RECT 10.715000 7.600000 10.885000 7.770000 ;
        RECT 11.195000 7.600000 11.365000 7.770000 ;
        RECT 11.675000 7.600000 11.845000 7.770000 ;
        RECT 12.155000 7.600000 12.325000 7.770000 ;
        RECT 12.635000 7.600000 12.805000 7.770000 ;
        RECT 13.115000 7.600000 13.285000 7.770000 ;
        RECT 13.590000 7.600000 13.760000 7.770000 ;
        RECT 14.075000 7.600000 14.245000 7.770000 ;
        RECT 14.555000 7.600000 14.725000 7.770000 ;
        RECT 17.820000 0.425000 17.990000 0.595000 ;
        RECT 17.820000 7.545000 17.990000 7.715000 ;
        RECT 18.300000 0.425000 18.470000 0.595000 ;
        RECT 18.300000 7.545000 18.470000 7.715000 ;
        RECT 18.780000 0.425000 18.950000 0.595000 ;
        RECT 18.780000 7.545000 18.950000 7.715000 ;
        RECT 19.260000 0.425000 19.430000 0.595000 ;
        RECT 19.260000 7.545000 19.430000 7.715000 ;
        RECT 19.740000 0.425000 19.910000 0.595000 ;
        RECT 19.740000 7.545000 19.910000 7.715000 ;
        RECT 20.220000 7.545000 20.390000 7.715000 ;
        RECT 20.700000 7.545000 20.870000 7.715000 ;
        RECT 21.180000 7.545000 21.350000 7.715000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 24.960000 0.625000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 24.960000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 24.960000 0.085000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000000 8.055000 24.960000 8.225000 ;
    END
    PORT
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.155000  8.055000  0.325000 8.225000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  0.635000  8.055000  0.805000 8.225000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.115000  8.055000  1.285000 8.225000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  1.595000  8.055000  1.765000 8.225000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.075000  8.055000  2.245000 8.225000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  2.555000  8.055000  2.725000 8.225000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.035000  8.055000  3.205000 8.225000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.515000  8.055000  3.685000 8.225000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  3.995000  8.055000  4.165000 8.225000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.475000  8.055000  4.645000 8.225000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  4.955000  8.055000  5.125000 8.225000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.435000  8.055000  5.605000 8.225000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  5.915000  8.055000  6.085000 8.225000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.395000  8.055000  6.565000 8.225000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  6.875000  8.055000  7.045000 8.225000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.355000  8.055000  7.525000 8.225000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  7.835000  8.055000  8.005000 8.225000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.315000  8.055000  8.485000 8.225000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  8.795000  8.055000  8.965000 8.225000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.275000  8.055000  9.445000 8.225000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT  9.755000  8.055000  9.925000 8.225000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.235000  8.055000 10.405000 8.225000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 10.715000  8.055000 10.885000 8.225000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.195000  8.055000 11.365000 8.225000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 11.675000  8.055000 11.845000 8.225000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.155000  8.055000 12.325000 8.225000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 12.635000  8.055000 12.805000 8.225000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.115000  8.055000 13.285000 8.225000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 13.595000  8.055000 13.765000 8.225000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.075000  8.055000 14.245000 8.225000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 14.555000  8.055000 14.725000 8.225000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.035000  8.055000 15.205000 8.225000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
        RECT 15.515000  8.055000 15.685000 8.225000 ;
        RECT 15.995000 -0.085000 16.165000 0.085000 ;
        RECT 15.995000  8.055000 16.165000 8.225000 ;
        RECT 16.475000 -0.085000 16.645000 0.085000 ;
        RECT 16.475000  8.055000 16.645000 8.225000 ;
        RECT 16.955000 -0.085000 17.125000 0.085000 ;
        RECT 16.955000  8.055000 17.125000 8.225000 ;
        RECT 17.435000 -0.085000 17.605000 0.085000 ;
        RECT 17.435000  8.055000 17.605000 8.225000 ;
        RECT 17.915000 -0.085000 18.085000 0.085000 ;
        RECT 17.915000  8.055000 18.085000 8.225000 ;
        RECT 18.395000 -0.085000 18.565000 0.085000 ;
        RECT 18.395000  8.055000 18.565000 8.225000 ;
        RECT 18.875000 -0.085000 19.045000 0.085000 ;
        RECT 18.875000  8.055000 19.045000 8.225000 ;
        RECT 19.355000 -0.085000 19.525000 0.085000 ;
        RECT 19.355000  8.055000 19.525000 8.225000 ;
        RECT 19.835000 -0.085000 20.005000 0.085000 ;
        RECT 19.835000  8.055000 20.005000 8.225000 ;
        RECT 20.315000 -0.085000 20.485000 0.085000 ;
        RECT 20.315000  8.055000 20.485000 8.225000 ;
        RECT 20.795000 -0.085000 20.965000 0.085000 ;
        RECT 20.795000  8.055000 20.965000 8.225000 ;
        RECT 21.275000 -0.085000 21.445000 0.085000 ;
        RECT 21.275000  8.055000 21.445000 8.225000 ;
        RECT 21.755000 -0.085000 21.925000 0.085000 ;
        RECT 21.755000  8.055000 21.925000 8.225000 ;
        RECT 22.235000 -0.085000 22.405000 0.085000 ;
        RECT 22.235000  8.055000 22.405000 8.225000 ;
        RECT 22.715000 -0.085000 22.885000 0.085000 ;
        RECT 22.715000  8.055000 22.885000 8.225000 ;
        RECT 23.195000 -0.085000 23.365000 0.085000 ;
        RECT 23.195000  8.055000 23.365000 8.225000 ;
        RECT 23.675000 -0.085000 23.845000 0.085000 ;
        RECT 23.675000  8.055000 23.845000 8.225000 ;
        RECT 24.155000 -0.085000 24.325000 0.085000 ;
        RECT 24.155000  8.055000 24.325000 8.225000 ;
        RECT 24.635000 -0.085000 24.805000 0.085000 ;
        RECT 24.635000  8.055000 24.805000 8.225000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 24.960000 0.115000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 24.960000 8.255000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 0.685000 4.155000 ;
        RECT 0.360000 4.155000 0.530000 5.180000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.135000 3.985000 9.925000 4.155000 ;
    END
    PORT
      LAYER mcon ;
        RECT 0.155000 3.985000 0.325000 4.155000 ;
        RECT 0.515000 3.985000 0.685000 4.155000 ;
        RECT 9.265000 3.985000 9.435000 4.155000 ;
        RECT 9.625000 3.985000 9.795000 4.155000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 24.960000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.655000 4.395000 2.245000 4.625000 ;
        RECT 1.835000 2.405000 2.065000 4.395000 ;
        RECT 1.835000 4.625000 2.065000 5.115000 ;
    END
    PORT
      LAYER li1 ;
        RECT 10.025000 3.515000 10.615000 3.745000 ;
        RECT 10.210000 2.015000 10.430000 3.515000 ;
        RECT 10.210000 3.745000 10.430000 5.035000 ;
        RECT 10.210000 5.035000 13.550000 5.255000 ;
        RECT 11.585000 3.515000 12.175000 3.745000 ;
        RECT 11.770000 2.015000 11.990000 3.515000 ;
        RECT 11.770000 3.745000 11.990000 5.035000 ;
        RECT 13.145000 3.515000 13.735000 3.745000 ;
        RECT 13.330000 2.015000 13.550000 3.515000 ;
        RECT 13.330000 3.745000 13.550000 5.035000 ;
    END
    PORT
      LAYER li1 ;
        RECT 14.295000 4.395000 14.885000 4.625000 ;
        RECT 14.655000 4.265000 14.885000 4.395000 ;
        RECT 14.655000 4.625000 14.885000 5.055000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.215000 4.395000 3.805000 4.625000 ;
        RECT 3.395000 2.405000 3.625000 4.395000 ;
        RECT 3.395000 4.625000 3.625000 5.115000 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.725000 2.405000 4.955000 3.515000 ;
        RECT 4.725000 3.515000 5.310000 3.755000 ;
    END
    PORT
      LAYER mcon ;
        RECT  1.685000 4.425000  1.855000 4.595000 ;
        RECT  2.045000 4.425000  2.215000 4.595000 ;
        RECT  3.245000 4.425000  3.415000 4.595000 ;
        RECT  3.605000 4.425000  3.775000 4.595000 ;
        RECT  4.750000 3.545000  4.920000 3.715000 ;
        RECT  5.110000 3.545000  5.280000 3.715000 ;
        RECT 10.055000 3.545000 10.225000 3.715000 ;
        RECT 10.415000 3.545000 10.585000 3.715000 ;
        RECT 11.615000 3.545000 11.785000 3.715000 ;
        RECT 11.975000 3.545000 12.145000 3.715000 ;
        RECT 13.175000 3.545000 13.345000 3.715000 ;
        RECT 13.535000 3.545000 13.705000 3.715000 ;
        RECT 14.325000 4.425000 14.495000 4.595000 ;
        RECT 14.685000 4.425000 14.855000 4.595000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 24.960000 3.815000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 24.960000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  1.840000 5.755000  6.520000 5.975000 ;
      RECT  1.840000 5.975000  2.060000 6.525000 ;
      RECT  3.010000 1.865000  4.170000 1.920000 ;
      RECT  3.010000 1.920000  5.730000 2.140000 ;
      RECT  3.010000 2.140000  4.170000 2.195000 ;
      RECT  3.570000 5.975000  3.790000 7.205000 ;
      RECT  3.950000 0.645000  4.170000 1.865000 ;
      RECT  3.950000 2.195000  4.170000 3.755000 ;
      RECT  5.510000 0.645000  5.730000 1.920000 ;
      RECT  5.510000 2.140000  5.730000 3.755000 ;
      RECT  5.930000 5.975000  6.150000 7.205000 ;
      RECT  6.300000 2.185000  6.995000 2.515000 ;
      RECT  6.300000 2.515000  6.520000 5.755000 ;
      RECT  7.075000 2.835000  7.435000 3.065000 ;
      RECT  7.075000 3.065000  7.305000 4.345000 ;
      RECT  7.205000 2.425000  7.805000 2.655000 ;
      RECT  7.205000 2.655000  7.435000 2.835000 ;
      RECT  7.345000 4.905000  8.080000 5.235000 ;
      RECT  7.575000 1.585000 12.770000 1.805000 ;
      RECT  7.575000 1.805000  7.805000 2.425000 ;
      RECT  7.860000 2.835000  8.080000 4.905000 ;
      RECT  7.860000 5.235000  8.080000 5.755000 ;
      RECT  7.860000 5.755000 12.775000 5.975000 ;
      RECT  8.290000 5.975000  8.510000 7.205000 ;
      RECT 10.650000 5.975000 10.870000 7.205000 ;
      RECT 10.990000 1.805000 11.210000 4.725000 ;
      RECT 12.550000 1.805000 12.770000 4.725000 ;
      RECT 12.555000 5.975000 12.775000 6.525000 ;
      RECT 13.090000 5.425000 14.105000 5.755000 ;
      RECT 13.885000 4.265000 14.105000 5.425000 ;
      RECT 13.885000 5.755000 14.105000 6.865000 ;
      RECT 13.965000 1.345000 18.530000 1.395000 ;
      RECT 13.965000 1.395000 19.940000 1.565000 ;
      RECT 13.965000 1.565000 14.295000 2.285000 ;
      RECT 17.160000 1.735000 19.465000 2.165000 ;
      RECT 17.160000 2.165000 17.380000 5.635000 ;
      RECT 17.160000 5.635000 19.465000 5.805000 ;
      RECT 17.160000 5.805000 18.020000 5.855000 ;
      RECT 17.790000 5.855000 18.020000 6.575000 ;
      RECT 17.790000 6.575000 19.450000 6.745000 ;
      RECT 18.235000 4.775000 18.565000 5.635000 ;
      RECT 18.265000 2.335000 19.940000 2.505000 ;
      RECT 18.265000 2.505000 18.595000 3.365000 ;
      RECT 18.265000 5.975000 19.940000 6.185000 ;
      RECT 18.265000 6.185000 20.900000 6.405000 ;
      RECT 18.280000 0.795000 18.530000 1.345000 ;
      RECT 18.290000 6.745000 18.460000 7.345000 ;
      RECT 19.135000 4.775000 19.465000 5.635000 ;
      RECT 19.165000 2.505000 19.495000 3.365000 ;
      RECT 19.200000 6.745000 19.450000 7.345000 ;
      RECT 19.270000 0.795000 19.440000 1.395000 ;
      RECT 19.710000 1.565000 19.940000 2.335000 ;
      RECT 20.615000 4.775000 20.900000 6.185000 ;
      RECT 20.615000 6.405000 20.900000 6.625000 ;
      RECT 20.615000 6.625000 20.945000 7.345000 ;
  END
END sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3
