* File: sky130_fd_sc_hvl__a21o_1.pex.spice
* Created: Fri Aug 28 09:32:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__A21O_1%VNB 5 7 11 25
r26 7 25 2.89352e-05 $w=4.32e-06 $l=1e-09 $layer=MET1_cond $X=2.16 $Y=0.057
+ $X2=2.16 $Y2=0.058
r27 7 11 0.00164931 $w=4.32e-06 $l=5.7e-08 $layer=MET1_cond $X=2.16 $Y=0.057
+ $X2=2.16 $Y2=0
r28 5 11 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r29 5 11 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__A21O_1%VPB 4 6 14 21
r42 10 21 0.00164931 $w=4.32e-06 $l=5.7e-08 $layer=MET1_cond $X=2.16 $Y=4.07
+ $X2=2.16 $Y2=4.013
r43 10 14 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=4.07
+ $X2=4.08 $Y2=4.07
r44 9 14 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=4.08 $Y2=4.07
r45 9 10 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r46 6 21 2.89352e-05 $w=4.32e-06 $l=1e-09 $layer=MET1_cond $X=2.16 $Y=4.012
+ $X2=2.16 $Y2=4.013
r47 4 14 40.4444 $w=1.7e-07 $l=4.12228e-06 $layer=licon1_NTAP_notbjt $count=4
+ $X=0 $Y=3.985 $X2=4.08 $Y2=4.07
r48 4 9 40.4444 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=4
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__A21O_1%A_83_283# 1 2 9 13 15 19 23 27 30 32 33 37
+ 38
r62 33 41 19.0324 $w=6e-07 $l=1.95e-07 $layer=POLY_cond $X=0.715 $Y=1.89
+ $X2=0.715 $Y2=2.085
r63 33 40 44.0004 $w=6e-07 $l=4.75e-07 $layer=POLY_cond $X=0.715 $Y=1.89
+ $X2=0.715 $Y2=1.415
r64 32 35 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.73 $Y=1.89
+ $X2=0.73 $Y2=2.015
r65 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.73
+ $Y=1.89 $X2=0.73 $Y2=1.89
r66 30 38 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.54 $Y=1.93
+ $X2=2.54 $Y2=1.325
r67 25 38 6.49277 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.555 $Y=1.2
+ $X2=2.555 $Y2=1.325
r68 25 27 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=2.555 $Y=1.2
+ $X2=2.555 $Y2=0.66
r69 24 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.87 $Y=2.015
+ $X2=1.745 $Y2=2.015
r70 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.455 $Y=2.015
+ $X2=2.54 $Y2=1.93
r71 23 24 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.455 $Y=2.015
+ $X2=1.87 $Y2=2.015
r72 19 21 57.6222 $w=2.48e-07 $l=1.25e-06 $layer=LI1_cond $X=1.745 $Y=2.34
+ $X2=1.745 $Y2=3.59
r73 17 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.745 $Y=2.1
+ $X2=1.745 $Y2=2.015
r74 17 19 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=1.745 $Y=2.1
+ $X2=1.745 $Y2=2.34
r75 16 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.015
+ $X2=0.73 $Y2=2.015
r76 15 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.62 $Y=2.015
+ $X2=1.745 $Y2=2.015
r77 15 16 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.62 $Y=2.015
+ $X2=0.895 $Y2=2.015
r78 13 40 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.765 $Y=0.91
+ $X2=0.765 $Y2=1.415
r79 9 41 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.665 $Y=2.965
+ $X2=0.665 $Y2=2.085
r80 2 21 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=1.56
+ $Y=2.215 $X2=1.705 $Y2=3.59
r81 2 19 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.56
+ $Y=2.215 $X2=1.705 $Y2=2.34
r82 1 27 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.375
+ $Y=0.535 $X2=2.515 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__A21O_1%B1 3 7 9 10 11 16
r34 16 19 29.0039 $w=5.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.11 $Y=1.63
+ $X2=2.11 $Y2=1.915
r35 16 18 21.9375 $w=5.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.11 $Y=1.63
+ $X2=2.11 $Y2=1.415
r36 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.03
+ $Y=1.63 $X2=2.03 $Y2=1.63
r37 11 17 6.115 $w=2.43e-07 $l=1.3e-07 $layer=LI1_cond $X=2.16 $Y=1.627 $X2=2.03
+ $Y2=1.627
r38 10 17 16.4635 $w=2.43e-07 $l=3.5e-07 $layer=LI1_cond $X=1.68 $Y=1.627
+ $X2=2.03 $Y2=1.627
r39 9 10 22.5785 $w=2.43e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.627 $X2=1.68
+ $Y2=1.627
r40 7 18 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.125 $Y=0.91 $X2=2.125
+ $Y2=1.415
r41 3 19 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.095 $Y=2.965
+ $X2=2.095 $Y2=1.915
.ends

.subckt PM_SKY130_FD_SC_HVL__A21O_1%A1 3 7 9 10 14
r34 14 17 24.9659 $w=5.3e-07 $l=2.45e-07 $layer=POLY_cond $X=2.89 $Y=1.67
+ $X2=2.89 $Y2=1.915
r35 14 16 25.9754 $w=5.3e-07 $l=2.55e-07 $layer=POLY_cond $X=2.89 $Y=1.67
+ $X2=2.89 $Y2=1.415
r36 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.97
+ $Y=1.67 $X2=2.97 $Y2=1.67
r37 9 10 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.67 $X2=3.6
+ $Y2=1.67
r38 9 15 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.12 $Y=1.67 $X2=2.97
+ $Y2=1.67
r39 7 16 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.905 $Y=0.91 $X2=2.905
+ $Y2=1.415
r40 3 17 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.875 $Y=2.965
+ $X2=2.875 $Y2=1.915
.ends

.subckt PM_SKY130_FD_SC_HVL__A21O_1%A2 3 7 9 15
r24 13 15 29.9457 $w=6.7e-07 $l=3.75e-07 $layer=POLY_cond $X=3.655 $Y=1.75
+ $X2=4.03 $Y2=1.75
r25 11 13 3.19421 $w=6.7e-07 $l=4e-08 $layer=POLY_cond $X=3.615 $Y=1.75
+ $X2=3.655 $Y2=1.75
r26 9 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.03
+ $Y=1.67 $X2=4.03 $Y2=1.67
r27 5 13 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.655 $Y=2.085
+ $X2=3.655 $Y2=1.75
r28 5 7 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.655 $Y=2.085 $X2=3.655
+ $Y2=2.965
r29 1 11 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.615 $Y=1.415
+ $X2=3.615 $Y2=1.75
r30 1 3 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.615 $Y=1.415 $X2=3.615
+ $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HVL__A21O_1%X 1 2 7 8 9 10 11 12 13 24 46
r16 46 47 1.94566 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=0.285 $Y=1.295
+ $X2=0.285 $Y2=1.325
r17 13 42 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=0.235 $Y=3.145
+ $X2=0.235 $Y2=3.57
r18 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=2.775
+ $X2=0.235 $Y2=3.145
r19 11 12 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=0.235 $Y=2.36
+ $X2=0.235 $Y2=2.775
r20 10 11 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=0.235 $Y=2.035
+ $X2=0.235 $Y2=2.36
r21 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.665
+ $X2=0.235 $Y2=2.035
r22 8 46 0.921954 $w=3.48e-07 $l=2.8e-08 $layer=LI1_cond $X=0.285 $Y=1.267
+ $X2=0.285 $Y2=1.295
r23 8 22 3.85245 $w=3.48e-07 $l=1.17e-07 $layer=LI1_cond $X=0.285 $Y=1.267
+ $X2=0.285 $Y2=1.15
r24 8 9 14.4286 $w=2.48e-07 $l=3.13e-07 $layer=LI1_cond $X=0.235 $Y=1.352
+ $X2=0.235 $Y2=1.665
r25 8 47 1.24464 $w=2.48e-07 $l=2.7e-08 $layer=LI1_cond $X=0.235 $Y=1.352
+ $X2=0.235 $Y2=1.325
r26 7 22 7.40856 $w=3.48e-07 $l=2.25e-07 $layer=LI1_cond $X=0.285 $Y=0.925
+ $X2=0.285 $Y2=1.15
r27 7 24 8.72564 $w=3.48e-07 $l=2.65e-07 $layer=LI1_cond $X=0.285 $Y=0.925
+ $X2=0.285 $Y2=0.66
r28 2 42 300 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.215 $X2=0.275 $Y2=3.57
r29 2 11 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.215 $X2=0.275 $Y2=2.36
r30 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.23
+ $Y=0.535 $X2=0.375 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__A21O_1%VPWR 1 2 7 10 20 27
r34 24 27 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.945 $Y=3.63
+ $X2=3.665 $Y2=3.63
r35 23 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.665 $Y=3.59
+ $X2=3.665 $Y2=3.59
r36 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.945 $Y=3.59
+ $X2=2.945 $Y2=3.59
r37 20 23 11.2368 $w=9.48e-07 $l=8.75e-07 $layer=LI1_cond $X=3.305 $Y=2.715
+ $X2=3.305 $Y2=3.59
r38 14 17 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.63 $Y=3.63
+ $X2=1.35 $Y2=3.63
r39 13 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.35 $Y=3.59
+ $X2=1.35 $Y2=3.59
r40 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.63 $Y=3.59
+ $X2=0.63 $Y2=3.59
r41 10 13 16.6056 $w=8.98e-07 $l=1.225e-06 $layer=LI1_cond $X=0.99 $Y=2.365
+ $X2=0.99 $Y2=3.59
r42 7 24 0.301366 $w=3.7e-07 $l=7.85e-07 $layer=MET1_cond $X=2.16 $Y=3.63
+ $X2=2.945 $Y2=3.63
r43 7 17 0.310963 $w=3.7e-07 $l=8.1e-07 $layer=MET1_cond $X=2.16 $Y=3.63
+ $X2=1.35 $Y2=3.63
r44 2 23 400 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=1 $X=3.125
+ $Y=2.215 $X2=3.265 $Y2=3.59
r45 2 20 400 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_PDIFF $count=1 $X=3.125
+ $Y=2.215 $X2=3.265 $Y2=2.715
r46 1 13 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=0.915
+ $Y=2.215 $X2=1.055 $Y2=3.59
r47 1 10 300 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=2 $X=0.915
+ $Y=2.215 $X2=1.055 $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_HVL__A21O_1%A_469_443# 1 2 7 9 11 13 15
r29 15 17 37.3392 $w=2.48e-07 $l=8.1e-07 $layer=LI1_cond $X=4.085 $Y=2.76
+ $X2=4.085 $Y2=3.57
r30 13 22 3.08894 $w=2.5e-07 $l=1.28e-07 $layer=LI1_cond $X=4.085 $Y=2.45
+ $X2=4.085 $Y2=2.322
r31 13 15 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=4.085 $Y=2.45
+ $X2=4.085 $Y2=2.76
r32 12 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=2.365
+ $X2=2.485 $Y2=2.365
r33 11 22 4.05423 $w=1.7e-07 $l=1.44914e-07 $layer=LI1_cond $X=3.96 $Y=2.365
+ $X2=4.085 $Y2=2.322
r34 11 12 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=3.96 $Y=2.365
+ $X2=2.65 $Y2=2.365
r35 7 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=2.45 $X2=2.485
+ $Y2=2.365
r36 7 9 39.8117 $w=3.28e-07 $l=1.14e-06 $layer=LI1_cond $X=2.485 $Y=2.45
+ $X2=2.485 $Y2=3.59
r37 2 22 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=2.215 $X2=4.045 $Y2=2.36
r38 2 17 400 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=2.215 $X2=4.045 $Y2=3.57
r39 2 15 400 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=2.215 $X2=4.045 $Y2=2.76
r40 1 20 300 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=2 $X=2.345
+ $Y=2.215 $X2=2.485 $Y2=2.365
r41 1 9 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.345
+ $Y=2.215 $X2=2.485 $Y2=3.59
.ends

.subckt PM_SKY130_FD_SC_HVL__A21O_1%VGND 1 2 7 10 25 26
r29 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.055 $Y=0.48
+ $X2=4.055 $Y2=0.48
r30 23 25 0.635417 $w=9.58e-07 $l=5e-08 $layer=LI1_cond $X=4.005 $Y=0.845
+ $X2=4.055 $Y2=0.845
r31 20 26 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=2.975 $Y=0.44
+ $X2=4.055 $Y2=0.44
r32 19 23 13.0896 $w=9.58e-07 $l=1.03e-06 $layer=LI1_cond $X=2.975 $Y=0.845
+ $X2=4.005 $Y2=0.845
r33 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.975 $Y=0.48
+ $X2=2.975 $Y2=0.48
r34 10 16 1.36398 $w=1.608e-06 $l=1.8e-07 $layer=LI1_cond $X=1.445 $Y=0.48
+ $X2=1.445 $Y2=0.66
r35 10 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.725 $Y=0.48
+ $X2=0.725 $Y2=0.48
r36 7 20 0.312883 $w=3.7e-07 $l=8.15e-07 $layer=MET1_cond $X=2.16 $Y=0.44
+ $X2=2.975 $Y2=0.44
r37 7 11 0.550904 $w=3.7e-07 $l=1.435e-06 $layer=MET1_cond $X=2.16 $Y=0.44
+ $X2=0.725 $Y2=0.44
r38 7 10 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.165 $Y=0.48
+ $X2=2.165 $Y2=0.48
r39 2 23 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.865
+ $Y=0.535 $X2=4.005 $Y2=0.66
r40 1 16 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.535 $X2=1.155 $Y2=0.66
.ends

