* File: sky130_fd_sc_hvl__sdfxtp_1.spice
* Created: Wed Sep  2 09:10:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__sdfxtp_1.pex.spice"
.subckt sky130_fd_sc_hvl__sdfxtp_1  VNB VPB SCE D SCD CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_SCE_M1011_g N_A_30_593#_M1011_s N_VNB_M1011_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250004 A=0.21 P=1.84 MULT=1
MM1025 A_342_107# N_D_M1025_g N_VGND_M1011_d N_VNB_M1011_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84 SA=250001
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1027 N_A_484_107#_M1027_d N_A_30_593#_M1027_g A_342_107# N_VNB_M1011_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1015 A_640_107# N_SCE_M1015_g N_A_484_107#_M1027_d N_VNB_M1011_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1018 N_VGND_M1018_d N_SCD_M1018_g A_640_107# N_VNB_M1011_b NHV L=0.5 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250003
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1008 N_A_938_107#_M1008_d N_CLK_M1008_g N_VGND_M1018_d N_VNB_M1011_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250004
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1019 N_A_1204_107#_M1019_d N_A_938_107#_M1019_g N_VGND_M1019_s N_VNB_M1011_b
+ NHV L=0.5 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1028 N_A_1490_107#_M1028_d N_A_938_107#_M1028_g N_A_484_107#_M1028_s
+ N_VNB_M1011_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.1533 PD=0.7 PS=1.57 NRD=0
+ NRS=21.7056 M=1 R=0.84 SA=250000 SB=250006 A=0.21 P=1.84 MULT=1
MM1021 A_1646_107# N_A_1204_107#_M1021_g N_A_1490_107#_M1028_d N_VNB_M1011_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250001 SB=250005 A=0.21 P=1.84 MULT=1
MM1022 N_VGND_M1022_d N_A_1688_81#_M1022_g A_1646_107# N_VNB_M1011_b NHV L=0.5
+ W=0.42 AD=0.0933154 AS=0.0441 PD=0.822051 PS=0.63 NRD=31.2132 NRS=13.566 M=1
+ R=0.84 SA=250002 SB=250004 A=0.21 P=1.84 MULT=1
MM1013 N_A_1688_81#_M1013_d N_A_1490_107#_M1013_g N_VGND_M1022_d N_VNB_M1011_b
+ NHV L=0.5 W=0.75 AD=0.166635 AS=0.166635 PD=1.46795 PS=1.46795 NRD=0 NRS=0 M=1
+ R=1.5 SA=250001 SB=250002 A=0.375 P=2.5 MULT=1
MM1029 N_A_2123_543#_M1029_d N_A_1204_107#_M1029_g N_A_1688_81#_M1013_d
+ N_VNB_M1011_b NHV L=0.5 W=0.42 AD=0.0672 AS=0.0933154 PD=0.74 PS=0.822051
+ NRD=10.8528 NRS=31.2132 M=1 R=0.84 SA=250003 SB=250002 A=0.21 P=1.84 MULT=1
MM1000 A_2310_107# N_A_938_107#_M1000_g N_A_2123_543#_M1029_d N_VNB_M1011_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250004 SB=250002 A=0.21 P=1.84 MULT=1
MM1001 N_VGND_M1001_d N_A_2352_81#_M1001_g A_2310_107# N_VNB_M1011_b NHV L=0.5
+ W=0.42 AD=0.0879308 AS=0.0441 PD=0.807692 PS=0.63 NRD=25.7754 NRS=13.566 M=1
+ R=0.84 SA=250005 SB=250001 A=0.21 P=1.84 MULT=1
MM1002 N_A_2352_81#_M1002_d N_A_2123_543#_M1002_g N_VGND_M1001_d N_VNB_M1011_b
+ NHV L=0.5 W=0.75 AD=0.19875 AS=0.157019 PD=2.03 PS=1.44231 NRD=0 NRS=0 M=1
+ R=1.5 SA=250003 SB=250000 A=0.375 P=2.5 MULT=1
MM1012 N_VGND_M1012_d N_A_2352_81#_M1012_g N_Q_M1012_s N_VNB_M1011_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1003 N_VPWR_M1003_d N_SCE_M1003_g N_A_30_593#_M1003_s N_VPB_M1003_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250004 A=0.21 P=1.84 MULT=1
MM1014 A_343_593# N_SCE_M1014_g N_VPWR_M1003_d N_VPB_M1003_b PHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84 SA=250001
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1016 N_A_484_107#_M1016_d N_D_M1016_g A_343_593# N_VPB_M1003_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1006 A_641_593# N_A_30_593#_M1006_g N_A_484_107#_M1016_d N_VPB_M1003_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1007 N_VPWR_M1007_d N_SCD_M1007_g A_641_593# N_VPB_M1003_b PHV L=0.5 W=0.42
+ AD=0.0879308 AS=0.0441 PD=0.807692 PS=0.63 NRD=43.1851 NRS=22.729 M=1 R=0.84
+ SA=250003 SB=250001 A=0.21 P=1.84 MULT=1
MM1009 N_A_938_107#_M1009_d N_CLK_M1009_g N_VPWR_M1007_d N_VPB_M1003_b PHV L=0.5
+ W=0.75 AD=0.19875 AS=0.157019 PD=2.03 PS=1.44231 NRD=0 NRS=0 M=1 R=1.5
+ SA=250002 SB=250000 A=0.375 P=2.5 MULT=1
MM1020 N_A_1204_107#_M1020_d N_A_938_107#_M1020_g N_VPWR_M1020_s N_VPB_M1003_b
+ PHV L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1030 N_A_1490_107#_M1030_d N_A_1204_107#_M1030_g N_A_484_107#_M1030_s
+ N_VPB_M1003_b PHV L=0.5 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250006 A=0.21 P=1.84 MULT=1
MM1024 A_1646_543# N_A_938_107#_M1024_g N_A_1490_107#_M1030_d N_VPB_M1003_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250001 SB=250005 A=0.21 P=1.84 MULT=1
MM1026 N_VPWR_M1026_d N_A_1688_81#_M1026_g A_1646_543# N_VPB_M1003_b PHV L=0.5
+ W=0.42 AD=0.0979606 AS=0.0441 PD=0.825211 PS=0.63 NRD=81.0413 NRS=22.729 M=1
+ R=0.84 SA=250002 SB=250004 A=0.21 P=1.84 MULT=1
MM1017 N_A_1688_81#_M1017_d N_A_1490_107#_M1017_g N_VPWR_M1026_d N_VPB_M1003_b
+ PHV L=0.5 W=1 AD=0.14 AS=0.233239 PD=1.28 PS=1.96479 NRD=0 NRS=0 M=1 R=2
+ SA=250001 SB=250002 A=0.5 P=3 MULT=1
MM1031 N_A_2123_543#_M1031_d N_A_938_107#_M1031_g N_A_1688_81#_M1017_d
+ N_VPB_M1003_b PHV L=0.5 W=1 AD=0.233239 AS=0.14 PD=1.96479 PS=1.28 NRD=0 NRS=0
+ M=1 R=2 SA=250002 SB=250001 A=0.5 P=3 MULT=1
MM1023 A_2302_543# N_A_1204_107#_M1023_g N_A_2123_543#_M1031_d N_VPB_M1003_b PHV
+ L=0.5 W=0.42 AD=0.0525 AS=0.0979606 PD=0.67 PS=0.825211 NRD=31.8206
+ NRS=52.2958 M=1 R=0.84 SA=250004 SB=250002 A=0.21 P=1.84 MULT=1
MM1004 N_VPWR_M1004_d N_A_2352_81#_M1004_g A_2302_543# N_VPB_M1003_b PHV L=0.5
+ W=0.42 AD=0.0920451 AS=0.0525 PD=0.81338 PS=0.67 NRD=43.1851 NRS=31.8206 M=1
+ R=0.84 SA=250005 SB=250001 A=0.21 P=1.84 MULT=1
MM1005 N_A_2352_81#_M1005_d N_A_2123_543#_M1005_g N_VPWR_M1004_d N_VPB_M1003_b
+ PHV L=0.5 W=1 AD=0.265 AS=0.219155 PD=2.53 PS=1.93662 NRD=0 NRS=0 M=1 R=2
+ SA=250002 SB=250000 A=0.5 P=3 MULT=1
MM1010 N_VPWR_M1010_d N_A_2352_81#_M1010_g N_Q_M1010_s N_VPB_M1003_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.3975 PD=3.53 PS=3.53 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
DX32_noxref N_VNB_M1011_b N_VPB_M1003_b NWDIODE A=40.404 P=36.28
*
.include "sky130_fd_sc_hvl__sdfxtp_1.pxi.spice"
*
.ends
*
*
