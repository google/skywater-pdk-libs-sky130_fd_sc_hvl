* File: sky130_fd_sc_hvl__sdfsbp_1.pex.spice
* Created: Fri Aug 28 09:39:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%VNB 5 7 11
c135 11 0 3.94641e-20 $X=0.24 $Y=0
c136 5 0 6.84108e-20 $X=-0.33 $Y=-0.265
r137 7 11 0.000353423 $w=2.016e-05 $l=5.7e-08 $layer=MET1_cond $X=10.08 $Y=0.057
+ $X2=10.08 $Y2=0
r138 5 11 0.442857 $w=1.7e-07 $l=3.57e-06 $layer=mcon $count=21 $X=19.92 $Y=0
+ $X2=19.92 $Y2=0
r139 5 11 0.442857 $w=1.7e-07 $l=3.57e-06 $layer=mcon $count=21 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%VPB 4 6 14
r162 10 14 0.442857 $w=1.7e-07 $l=3.57e-06 $layer=mcon $count=21 $X=19.92
+ $Y=4.07 $X2=19.92 $Y2=4.07
r163 9 14 1283.94 $w=1.68e-07 $l=1.968e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=19.92 $Y2=4.07
r164 9 10 0.442857 $w=1.7e-07 $l=3.57e-06 $layer=mcon $count=21 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r165 6 10 0.000353423 $w=2.016e-05 $l=5.7e-08 $layer=MET1_cond $X=10.08 $Y=4.013
+ $X2=10.08 $Y2=4.07
r166 4 14 8.66667 $w=1.7e-07 $l=1.99625e-05 $layer=licon1_NTAP_notbjt $count=21
+ $X=0 $Y=3.985 $X2=19.92 $Y2=4.07
r167 4 9 8.66667 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=21
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%SCE 1 3 6 8 10 13 14 22 24 26 27 32 33 34
+ 39 42 45 53
r77 34 53 9.71911 $w=6.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.83
+ $X2=1.795 $Y2=1.83
r78 34 45 3.92742 $w=6.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.68 $Y=1.83
+ $X2=1.46 $Y2=1.83
r79 33 45 4.6415 $w=6.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.2 $Y=1.83 $X2=1.46
+ $Y2=1.83
r80 32 33 8.56892 $w=6.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.83 $X2=1.2
+ $Y2=1.83
r81 32 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.775
+ $Y=1.66 $X2=0.775 $Y2=1.66
r82 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.845
+ $Y=1.6 $X2=2.845 $Y2=1.6
r83 27 31 31.914 $w=5.7e-07 $l=3.4e-07 $layer=POLY_cond $X=2.945 $Y=1.26
+ $X2=2.945 $Y2=1.6
r84 27 42 18.3095 $w=5.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.945 $Y=1.26
+ $X2=2.945 $Y2=1.075
r85 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.845
+ $Y=1.26 $X2=2.845 $Y2=1.26
r86 24 30 3.0698 $w=2.75e-07 $l=1.35e-07 $layer=LI1_cond $X=2.817 $Y=1.495
+ $X2=2.817 $Y2=1.63
r87 24 26 9.84815 $w=2.73e-07 $l=2.35e-07 $layer=LI1_cond $X=2.817 $Y=1.495
+ $X2=2.817 $Y2=1.26
r88 22 30 4.25224 $w=1.7e-07 $l=1.60059e-07 $layer=LI1_cond $X=2.68 $Y=1.58
+ $X2=2.817 $Y2=1.63
r89 22 53 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.68 $Y=1.58
+ $X2=1.795 $Y2=1.58
r90 19 39 67.2608 $w=5.25e-07 $l=6.6e-07 $layer=POLY_cond $X=0.697 $Y=2.32
+ $X2=0.697 $Y2=1.66
r91 14 39 31.8979 $w=5.25e-07 $l=3.13e-07 $layer=POLY_cond $X=0.697 $Y=1.347
+ $X2=0.697 $Y2=1.66
r92 14 15 26.8714 $w=5.25e-07 $l=2.62e-07 $layer=POLY_cond $X=0.697 $Y=1.347
+ $X2=0.697 $Y2=1.085
r93 13 42 31.812 $w=5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.98 $Y=0.745 $X2=2.98
+ $Y2=1.075
r94 8 19 102.922 $w=4.15e-07 $l=7.68e-07 $layer=POLY_cond $X=1.465 $Y=2.527
+ $X2=0.697 $Y2=2.527
r95 8 10 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.465 $Y=2.735 $X2=1.465
+ $Y2=3.055
r96 6 15 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.71 $Y=0.745 $X2=0.71
+ $Y2=1.085
r97 1 19 1.60816 $w=4.15e-07 $l=1.2e-08 $layer=POLY_cond $X=0.685 $Y=2.527
+ $X2=0.697 $Y2=2.527
r98 1 3 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.685 $Y=2.735 $X2=0.685
+ $Y2=3.055
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%D 3 5 7 9 15
c40 7 0 4.65845e-20 $X=2.175 $Y=3.055
r41 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.14
+ $Y=1.93 $X2=2.14 $Y2=1.93
r42 9 15 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.14 $Y=2.035
+ $X2=2.14 $Y2=1.93
r43 5 14 4.63462 $w=4.2e-07 $l=3.5e-08 $layer=POLY_cond $X=2.175 $Y=1.9 $X2=2.14
+ $Y2=1.9
r44 5 7 101.121 $w=5e-07 $l=9.45e-07 $layer=POLY_cond $X=2.175 $Y=2.11 $X2=2.175
+ $Y2=3.055
r45 1 14 86.0714 $w=4.2e-07 $l=6.5e-07 $layer=POLY_cond $X=1.49 $Y=1.9 $X2=2.14
+ $Y2=1.9
r46 1 3 101.121 $w=5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.49 $Y=1.69 $X2=1.49
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%A_30_569# 1 2 7 9 13 16 19 21 25 30 33 34
+ 36
c77 30 0 1.09754e-19 $X=2.8 $Y=2.18
c78 21 0 5.97692e-20 $X=2.635 $Y=2.62
r79 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.8 $Y=2.18
+ $X2=2.8 $Y2=2.18
r80 28 30 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=2.76 $Y=2.535
+ $X2=2.76 $Y2=2.18
r81 26 36 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.2 $Y=1.23 $X2=2.2
+ $Y2=0.745
r82 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.135
+ $Y=1.23 $X2=2.135 $Y2=1.23
r83 23 33 1.98564 $w=2.2e-07 $l=1.78e-07 $layer=LI1_cond $X=0.485 $Y=1.205
+ $X2=0.307 $Y2=1.205
r84 23 25 86.4332 $w=2.18e-07 $l=1.65e-06 $layer=LI1_cond $X=0.485 $Y=1.205
+ $X2=2.135 $Y2=1.205
r85 22 34 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.46 $Y=2.62
+ $X2=0.295 $Y2=2.62
r86 21 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.635 $Y=2.62
+ $X2=2.76 $Y2=2.535
r87 21 22 141.898 $w=1.68e-07 $l=2.175e-06 $layer=LI1_cond $X=2.635 $Y=2.62
+ $X2=0.46 $Y2=2.62
r88 17 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.295 $Y=2.705
+ $X2=0.295 $Y2=2.62
r89 17 19 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.295 $Y=2.705
+ $X2=0.295 $Y2=3.055
r90 16 34 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.215 $Y=2.535
+ $X2=0.295 $Y2=2.62
r91 15 33 4.44913 $w=2.62e-07 $l=1.49064e-07 $layer=LI1_cond $X=0.215 $Y=1.315
+ $X2=0.307 $Y2=1.205
r92 15 16 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=0.215 $Y=1.315
+ $X2=0.215 $Y2=2.535
r93 11 33 4.44913 $w=2.62e-07 $l=1.1e-07 $layer=LI1_cond $X=0.307 $Y=1.095
+ $X2=0.307 $Y2=1.205
r94 11 13 11.3621 $w=3.53e-07 $l=3.5e-07 $layer=LI1_cond $X=0.307 $Y=1.095
+ $X2=0.307 $Y2=0.745
r95 7 31 47.5188 $w=5.48e-07 $l=5.52223e-07 $layer=POLY_cond $X=2.955 $Y=2.715
+ $X2=2.92 $Y2=2.18
r96 7 9 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.955 $Y=2.715 $X2=2.955
+ $Y2=3.055
r97 2 19 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.845 $X2=0.295 $Y2=3.055
r98 1 13 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.535 $X2=0.32 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%SCD 3 7 8 9 10 11 17
c36 7 0 1.69523e-19 $X=3.677 $Y=2.715
c37 3 0 3.3847e-20 $X=3.665 $Y=3.055
r38 17 20 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.69 $Y=0.745
+ $X2=3.69 $Y2=1.27
r39 10 11 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=1.665
+ $X2=3.587 $Y2=2.035
r40 9 10 21.3703 $w=2.03e-07 $l=3.95e-07 $layer=LI1_cond $X=3.587 $Y=1.27
+ $X2=3.587 $Y2=1.665
r41 9 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.605
+ $Y=1.27 $X2=3.605 $Y2=1.27
r42 8 9 18.6652 $w=2.03e-07 $l=3.45e-07 $layer=LI1_cond $X=3.587 $Y=0.925
+ $X2=3.587 $Y2=1.27
r43 6 20 101.121 $w=5e-07 $l=9.45e-07 $layer=POLY_cond $X=3.69 $Y=2.215 $X2=3.69
+ $Y2=1.27
r44 6 7 50.9552 $w=5.25e-07 $l=5e-07 $layer=POLY_cond $X=3.677 $Y=2.215
+ $X2=3.677 $Y2=2.715
r45 3 7 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.665 $Y=3.055 $X2=3.665
+ $Y2=2.715
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%CLK 3 7 9 10 11 16
r38 16 19 53.6738 $w=5.25e-07 $l=5.25e-07 $layer=POLY_cond $X=4.622 $Y=1.645
+ $X2=4.622 $Y2=2.17
r39 16 18 19.0243 $w=5.25e-07 $l=1.85e-07 $layer=POLY_cond $X=4.622 $Y=1.645
+ $X2=4.622 $Y2=1.46
r40 10 11 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=4.545 $Y=1.645
+ $X2=4.545 $Y2=2.035
r41 10 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.545
+ $Y=1.645 $X2=4.545 $Y2=1.645
r42 9 10 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=4.545 $Y=1.295
+ $X2=4.545 $Y2=1.645
r43 7 18 76.5092 $w=5e-07 $l=7.15e-07 $layer=POLY_cond $X=4.635 $Y=0.745
+ $X2=4.635 $Y2=1.46
r44 3 19 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=4.61 $Y=3.22 $X2=4.61
+ $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%A_1243_116# 1 2 9 12 15 16 18 19 24 27 29
+ 31 32 35 39 42 45 46 47 48 50 51 52 54 56 57 58 61 67
c175 16 0 1.11272e-19 $X=13.185 $Y=2.605
c176 12 0 3.94641e-20 $X=12.43 $Y=0.91
r177 57 70 35.5806 $w=7.3e-07 $l=1.85e-07 $layer=POLY_cond $X=12.545 $Y=1.71
+ $X2=12.545 $Y2=1.895
r178 57 69 11.1291 $w=7.3e-07 $l=8.5e-08 $layer=POLY_cond $X=12.545 $Y=1.71
+ $X2=12.545 $Y2=1.625
r179 56 58 8.46257 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=12.365 $Y=1.717
+ $X2=12.2 $Y2=1.717
r180 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.365
+ $Y=1.71 $X2=12.365 $Y2=1.71
r181 51 67 20.8158 $w=6e-07 $l=2.15e-07 $layer=POLY_cond $X=7.47 $Y=2.455
+ $X2=7.47 $Y2=2.67
r182 50 52 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.355 $Y=2.455
+ $X2=7.355 $Y2=2.29
r183 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.355
+ $Y=2.455 $X2=7.355 $Y2=2.455
r184 46 47 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=6.48 $Y=1.02
+ $X2=6.48 $Y2=2.29
r185 45 58 252.807 $w=1.68e-07 $l=3.875e-06 $layer=LI1_cond $X=8.325 $Y=1.645
+ $X2=12.2 $Y2=1.645
r186 43 61 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.095 $Y=1.315
+ $X2=8.095 $Y2=0.81
r187 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.16
+ $Y=1.315 $X2=8.16 $Y2=1.315
r188 40 45 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=8.187 $Y=1.56
+ $X2=8.325 $Y2=1.645
r189 40 42 10.2672 $w=2.73e-07 $l=2.45e-07 $layer=LI1_cond $X=8.187 $Y=1.56
+ $X2=8.187 $Y2=1.315
r190 39 54 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=8.187 $Y=1.287
+ $X2=8.187 $Y2=1.15
r191 39 42 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=8.187 $Y=1.287
+ $X2=8.187 $Y2=1.315
r192 37 54 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=8.135 $Y=0.435
+ $X2=8.135 $Y2=1.15
r193 36 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=0.35
+ $X2=7.275 $Y2=0.35
r194 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.05 $Y=0.35
+ $X2=8.135 $Y2=0.435
r195 35 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.05 $Y=0.35
+ $X2=7.36 $Y2=0.35
r196 33 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.275 $Y=0.435
+ $X2=7.275 $Y2=0.35
r197 33 52 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=7.275 $Y=0.435
+ $X2=7.275 $Y2=2.29
r198 31 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.19 $Y=0.35
+ $X2=7.275 $Y2=0.35
r199 31 32 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=7.19 $Y=0.35
+ $X2=6.565 $Y2=0.35
r200 27 47 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.52 $Y=2.415
+ $X2=6.52 $Y2=2.29
r201 27 29 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=6.52 $Y=2.415
+ $X2=6.52 $Y2=2.585
r202 22 46 9.23056 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=6.377 $Y=0.833
+ $X2=6.377 $Y2=1.02
r203 22 24 1.32147 $w=3.73e-07 $l=4.3e-08 $layer=LI1_cond $X=6.377 $Y=0.833
+ $X2=6.377 $Y2=0.79
r204 21 32 8.1532 $w=1.7e-07 $l=2.26548e-07 $layer=LI1_cond $X=6.377 $Y=0.435
+ $X2=6.565 $Y2=0.35
r205 21 24 10.9098 $w=3.73e-07 $l=3.55e-07 $layer=LI1_cond $X=6.377 $Y=0.435
+ $X2=6.377 $Y2=0.79
r206 16 19 67.3138 $w=2.9e-07 $l=4.05e-07 $layer=POLY_cond $X=13.185 $Y=2.45
+ $X2=12.78 $Y2=2.45
r207 16 18 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=13.185 $Y=2.605
+ $X2=13.185 $Y2=2.925
r208 15 19 5.42818 $w=2.6e-07 $l=1.55e-07 $layer=POLY_cond $X=12.78 $Y=2.295
+ $X2=12.78 $Y2=2.45
r209 15 70 95.5591 $w=2.6e-07 $l=4e-07 $layer=POLY_cond $X=12.78 $Y=2.295
+ $X2=12.78 $Y2=1.895
r210 12 69 76.5092 $w=5e-07 $l=7.15e-07 $layer=POLY_cond $X=12.43 $Y=0.91
+ $X2=12.43 $Y2=1.625
r211 9 67 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.52 $Y=2.99 $X2=7.52
+ $Y2=2.67
r212 2 29 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.42
+ $Y=2.44 $X2=6.56 $Y2=2.585
r213 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.215
+ $Y=0.58 $X2=6.355 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%A_972_569# 1 2 9 13 15 17 19 20 22 24 26
+ 28 29 36 41 45 49 53 54 56 59 60 61 62 64 65 66 70 71 73 74 76 81 87
c213 65 0 1.11272e-19 $X=12.18 $Y=3
c214 61 0 9.67046e-20 $X=9.915 $Y=3.255
c215 56 0 1.0149e-19 $X=9.745 $Y=2.695
r216 94 95 41.6128 $w=7.05e-07 $l=5.1e-07 $layer=POLY_cond $X=6.067 $Y=1.38
+ $X2=6.067 $Y2=1.89
r217 86 87 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.19
+ $Y=2.29 $X2=12.19 $Y2=2.29
r218 81 83 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.69 $Y=3.085
+ $X2=10.69 $Y2=3.255
r219 77 96 52.3314 $w=5.25e-07 $l=5.7e-07 $layer=POLY_cond $X=8.28 $Y=2.455
+ $X2=8.28 $Y2=1.885
r220 76 79 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=8.365 $Y=2.455
+ $X2=8.365 $Y2=2.695
r221 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.365
+ $Y=2.455 $X2=8.365 $Y2=2.455
r222 70 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.285
+ $Y=1.58 $X2=13.285 $Y2=1.58
r223 68 70 26.1701 $w=2.38e-07 $l=5.45e-07 $layer=LI1_cond $X=13.285 $Y=2.125
+ $X2=13.285 $Y2=1.58
r224 67 86 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=12.335 $Y=2.21
+ $X2=12.18 $Y2=2.21
r225 66 68 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=13.165 $Y=2.21
+ $X2=13.285 $Y2=2.125
r226 66 67 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=13.165 $Y=2.21
+ $X2=12.335 $Y2=2.21
r227 64 86 2.69138 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=12.18 $Y=2.295
+ $X2=12.18 $Y2=2.21
r228 64 65 26.2088 $w=3.08e-07 $l=7.05e-07 $layer=LI1_cond $X=12.18 $Y=2.295
+ $X2=12.18 $Y2=3
r229 63 81 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.775 $Y=3.085
+ $X2=10.69 $Y2=3.085
r230 62 65 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=12.025 $Y=3.085
+ $X2=12.18 $Y2=3
r231 62 63 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=12.025 $Y=3.085
+ $X2=10.775 $Y2=3.085
r232 60 83 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.605 $Y=3.255
+ $X2=10.69 $Y2=3.255
r233 60 61 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.605 $Y=3.255
+ $X2=9.915 $Y2=3.255
r234 59 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.83 $Y=3.17
+ $X2=9.915 $Y2=3.255
r235 58 59 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=9.83 $Y=2.78
+ $X2=9.83 $Y2=3.17
r236 57 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.53 $Y=2.695
+ $X2=8.365 $Y2=2.695
r237 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.745 $Y=2.695
+ $X2=9.83 $Y2=2.78
r238 56 57 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=9.745 $Y=2.695
+ $X2=8.53 $Y2=2.695
r239 54 94 1.09398 $w=7.05e-07 $l=1.5e-08 $layer=POLY_cond $X=6.067 $Y=1.365
+ $X2=6.067 $Y2=1.38
r240 54 93 21.5565 $w=7.05e-07 $l=2.35e-07 $layer=POLY_cond $X=6.067 $Y=1.365
+ $X2=6.067 $Y2=1.13
r241 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.9
+ $Y=1.365 $X2=5.9 $Y2=1.365
r242 51 53 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.9 $Y=1.7 $X2=5.9
+ $Y2=1.365
r243 50 74 2.57001 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.19 $Y=1.785
+ $X2=5.065 $Y2=1.785
r244 49 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.735 $Y=1.785
+ $X2=5.9 $Y2=1.7
r245 49 50 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.735 $Y=1.785
+ $X2=5.19 $Y2=1.785
r246 47 74 3.87901 $w=2.37e-07 $l=9.12688e-08 $layer=LI1_cond $X=5.052 $Y=1.87
+ $X2=5.065 $Y2=1.785
r247 47 73 47.8904 $w=2.23e-07 $l=9.35e-07 $layer=LI1_cond $X=5.052 $Y=1.87
+ $X2=5.052 $Y2=2.805
r248 43 74 3.87901 $w=2.37e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=1.7
+ $X2=5.065 $Y2=1.785
r249 43 45 44.0233 $w=2.48e-07 $l=9.55e-07 $layer=LI1_cond $X=5.065 $Y=1.7
+ $X2=5.065 $Y2=0.745
r250 41 73 6.93655 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5 $Y=2.97 $X2=5
+ $Y2=2.805
r251 38 71 20.1682 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=13.347 $Y=1.415
+ $X2=13.347 $Y2=1.58
r252 36 38 36.9208 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=13.325 $Y=1.075
+ $X2=13.325 $Y2=1.415
r253 33 87 37.7162 $w=4.35e-07 $l=2.95e-07 $layer=POLY_cond $X=12.222 $Y=2.585
+ $X2=12.222 $Y2=2.29
r254 29 30 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.315 $Y=1.38
+ $X2=7.315 $Y2=1.885
r255 26 33 27.7985 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=12.255 $Y=2.835
+ $X2=12.255 $Y2=2.585
r256 26 28 36.632 $w=5e-07 $l=3.8e-07 $layer=POLY_cond $X=12.255 $Y=2.835
+ $X2=12.255 $Y2=3.215
r257 22 77 18.0568 $w=5.25e-07 $l=2.04756e-07 $layer=POLY_cond $X=8.3 $Y=2.65
+ $X2=8.28 $Y2=2.455
r258 22 24 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=8.3 $Y=2.65 $X2=8.3
+ $Y2=2.99
r259 21 30 11.1661 $w=3.5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.565 $Y=1.885
+ $X2=7.315 $Y2=1.885
r260 20 96 12.2893 $w=3.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.01 $Y=1.885
+ $X2=8.28 $Y2=1.885
r261 20 21 73.3668 $w=3.5e-07 $l=4.45e-07 $layer=POLY_cond $X=8.01 $Y=1.885
+ $X2=7.565 $Y2=1.885
r262 17 29 26.7515 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.315 $Y=1.13
+ $X2=7.315 $Y2=1.38
r263 17 19 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.315 $Y=1.13
+ $X2=7.315 $Y2=0.81
r264 16 94 10.8648 $w=5e-07 $l=3.53e-07 $layer=POLY_cond $X=6.42 $Y=1.38
+ $X2=6.067 $Y2=1.38
r265 15 29 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.065 $Y=1.38
+ $X2=7.315 $Y2=1.38
r266 15 16 69.0188 $w=5e-07 $l=6.45e-07 $layer=POLY_cond $X=7.065 $Y=1.38
+ $X2=6.42 $Y2=1.38
r267 13 95 98.9805 $w=5e-07 $l=9.25e-07 $layer=POLY_cond $X=6.17 $Y=2.815
+ $X2=6.17 $Y2=1.89
r268 9 93 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.965 $Y=0.79 $X2=5.965
+ $Y2=1.13
r269 2 41 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.86
+ $Y=2.845 $X2=5 $Y2=2.97
r270 1 45 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.885
+ $Y=0.535 $X2=5.025 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%A_1711_94# 1 2 9 10 13 15 18 22 26 31 34
c51 18 0 9.67046e-20 $X=9.075 $Y=2.345
r52 24 26 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=10.26 $Y=2.43
+ $X2=10.26 $Y2=2.905
r53 20 22 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=9.745 $Y=1.14
+ $X2=9.745 $Y2=0.745
r54 18 31 69.0188 $w=5e-07 $l=6.45e-07 $layer=POLY_cond $X=9.01 $Y=2.345
+ $X2=9.01 $Y2=2.99
r55 18 35 90.42 $w=5e-07 $l=8.45e-07 $layer=POLY_cond $X=9.01 $Y=2.345 $X2=9.01
+ $Y2=1.5
r56 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.075
+ $Y=2.345 $X2=9.075 $Y2=2.345
r57 15 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.095 $Y=2.345
+ $X2=10.26 $Y2=2.43
r58 15 17 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=10.095 $Y=2.345
+ $X2=9.075 $Y2=2.345
r59 13 35 19.3685 $w=7.05e-07 $l=2.05e-07 $layer=POLY_cond $X=8.907 $Y=1.295
+ $X2=8.907 $Y2=1.5
r60 13 34 16.4512 $w=7.05e-07 $l=1.65e-07 $layer=POLY_cond $X=8.907 $Y=1.295
+ $X2=8.907 $Y2=1.13
r61 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.075
+ $Y=1.295 $X2=9.075 $Y2=1.295
r62 10 20 7.03987 $w=2.4e-07 $l=2.16852e-07 $layer=LI1_cond $X=9.58 $Y=1.26
+ $X2=9.745 $Y2=1.14
r63 10 12 24.2493 $w=2.38e-07 $l=5.05e-07 $layer=LI1_cond $X=9.58 $Y=1.26
+ $X2=9.075 $Y2=1.26
r64 9 34 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.805 $Y=0.81 $X2=8.805
+ $Y2=1.13
r65 2 26 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=10.12
+ $Y=2.78 $X2=10.26 $Y2=2.905
r66 1 22 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.62
+ $Y=0.535 $X2=9.745 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%A_1513_120# 1 2 7 9 12 21 23 26 28 32 36
+ 39 41 42 45 49
c105 12 0 1.54156e-19 $X=11.72 $Y=0.91
r106 42 49 124.662 $w=5e-07 $l=1.165e-06 $layer=POLY_cond $X=11.545 $Y=2.05
+ $X2=11.545 $Y2=3.215
r107 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.48
+ $Y=2.05 $X2=11.48 $Y2=2.05
r108 36 38 11.4306 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=7.705 $Y=0.81
+ $X2=7.705 $Y2=1.06
r109 32 45 106.471 $w=5e-07 $l=9.95e-07 $layer=POLY_cond $X=9.87 $Y=1.995
+ $X2=9.87 $Y2=2.99
r110 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.935
+ $Y=1.995 $X2=9.935 $Y2=1.995
r111 29 39 2.49072 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=7.995 $Y=1.995
+ $X2=7.847 $Y2=1.995
r112 29 31 126.567 $w=1.68e-07 $l=1.94e-06 $layer=LI1_cond $X=7.995 $Y=1.995
+ $X2=9.935 $Y2=1.995
r113 28 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.315 $Y=1.995
+ $X2=11.48 $Y2=1.995
r114 28 31 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=11.315 $Y=1.995
+ $X2=9.935 $Y2=1.995
r115 24 39 3.95216 $w=2.32e-07 $l=8.5e-08 $layer=LI1_cond $X=7.847 $Y=2.08
+ $X2=7.847 $Y2=1.995
r116 24 26 35.5499 $w=2.93e-07 $l=9.1e-07 $layer=LI1_cond $X=7.847 $Y=2.08
+ $X2=7.847 $Y2=2.99
r117 23 39 3.95216 $w=2.32e-07 $l=1.11781e-07 $layer=LI1_cond $X=7.785 $Y=1.91
+ $X2=7.847 $Y2=1.995
r118 23 38 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=7.785 $Y=1.91
+ $X2=7.785 $Y2=1.06
r119 21 42 16.5859 $w=5e-07 $l=1.55e-07 $layer=POLY_cond $X=11.545 $Y=1.895
+ $X2=11.545 $Y2=2.05
r120 20 21 2.37791 $w=6.75e-07 $l=3e-08 $layer=POLY_cond $X=11.632 $Y=1.865
+ $X2=11.632 $Y2=1.895
r121 15 32 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=9.87 $Y=1.445
+ $X2=9.87 $Y2=1.995
r122 12 20 102.191 $w=5e-07 $l=9.55e-07 $layer=POLY_cond $X=11.72 $Y=0.91
+ $X2=11.72 $Y2=1.865
r123 7 15 38.7844 $w=3.8e-07 $l=2.65e-07 $layer=POLY_cond $X=10.135 $Y=1.255
+ $X2=9.87 $Y2=1.255
r124 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.135 $Y=1.065
+ $X2=10.135 $Y2=0.745
r125 2 26 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.77
+ $Y=2.78 $X2=7.91 $Y2=2.99
r126 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.565
+ $Y=0.6 $X2=7.705 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%SET_B 3 5 6 7 9 10 12 16 17 18 19 20 29 35
+ 39 41
c84 3 0 1.0149e-19 $X=10.65 $Y=2.99
r85 29 32 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=10.845 $Y=0.745
+ $X2=10.845 $Y2=1.295
r86 20 41 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.27 $Y=1.295
+ $X2=12.185 $Y2=1.295
r87 20 41 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=12.17 $Y=1.295
+ $X2=12.185 $Y2=1.295
r88 19 20 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=11.76 $Y=1.295
+ $X2=12.17 $Y2=1.295
r89 18 19 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=11.28 $Y=1.295
+ $X2=11.76 $Y2=1.295
r90 17 18 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=10.78 $Y=1.295
+ $X2=11.28 $Y2=1.295
r91 17 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.78
+ $Y=1.295 $X2=10.78 $Y2=1.295
r92 16 17 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=10.32 $Y=1.295
+ $X2=10.78 $Y2=1.295
r93 15 20 30.1177 $w=3.08e-07 $l=7.75e-07 $layer=LI1_cond $X=12.27 $Y=0.435
+ $X2=12.27 $Y2=1.21
r94 13 39 146.063 $w=5e-07 $l=1.365e-06 $layer=POLY_cond $X=14.745 $Y=1.56
+ $X2=14.745 $Y2=2.925
r95 13 35 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=14.745 $Y=1.56
+ $X2=14.745 $Y2=1.075
r96 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.68
+ $Y=1.56 $X2=14.68 $Y2=1.56
r97 10 12 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=14.17 $Y=1.535
+ $X2=14.68 $Y2=1.535
r98 9 10 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=14.085 $Y=1.425
+ $X2=14.17 $Y2=1.535
r99 8 9 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=14.085 $Y=0.435
+ $X2=14.085 $Y2=1.425
r100 7 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.355 $Y=0.35
+ $X2=12.27 $Y2=0.435
r101 6 8 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14 $Y=0.35
+ $X2=14.085 $Y2=0.435
r102 6 7 107.321 $w=1.68e-07 $l=1.645e-06 $layer=LI1_cond $X=14 $Y=0.35
+ $X2=12.355 $Y2=0.35
r103 5 32 11.7706 $w=5e-07 $l=1.1e-07 $layer=POLY_cond $X=10.845 $Y=1.405
+ $X2=10.845 $Y2=1.295
r104 1 5 58.0257 $w=6.23e-07 $l=8.41873e-07 $layer=POLY_cond $X=10.65 $Y=2.155
+ $X2=10.845 $Y2=1.405
r105 1 3 89.3499 $w=5e-07 $l=8.35e-07 $layer=POLY_cond $X=10.65 $Y=2.155
+ $X2=10.65 $Y2=2.99
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%A_2729_463# 1 2 9 12 13 20 28
r44 20 23 38.4148 $w=3.28e-07 $l=1.1e-06 $layer=LI1_cond $X=15.895 $Y=1.075
+ $X2=15.895 $Y2=2.175
r45 16 28 126.802 $w=5e-07 $l=1.185e-06 $layer=POLY_cond $X=14.035 $Y=2.26
+ $X2=14.035 $Y2=1.075
r46 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.1
+ $Y=2.26 $X2=14.1 $Y2=2.26
r47 13 25 5.07075 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=15.872 $Y=2.26
+ $X2=15.872 $Y2=2.425
r48 13 23 2.80732 $w=3.73e-07 $l=8.5e-08 $layer=LI1_cond $X=15.872 $Y=2.26
+ $X2=15.872 $Y2=2.175
r49 13 15 103.406 $w=1.68e-07 $l=1.585e-06 $layer=LI1_cond $X=15.685 $Y=2.26
+ $X2=14.1 $Y2=2.26
r50 11 16 5.88532 $w=5e-07 $l=5.5e-08 $layer=POLY_cond $X=14.035 $Y=2.315
+ $X2=14.035 $Y2=2.26
r51 11 12 24.2435 $w=6.4e-07 $l=2.9e-07 $layer=POLY_cond $X=13.965 $Y=2.315
+ $X2=13.965 $Y2=2.605
r52 9 12 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=13.895 $Y=2.925
+ $X2=13.895 $Y2=2.605
r53 2 25 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=15.705
+ $Y=2.215 $X2=15.85 $Y2=2.425
r54 1 20 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=15.75
+ $Y=0.865 $X2=15.895 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%A_2501_543# 1 2 3 10 12 13 15 18 20 22 23
+ 24 27 31 33 38 41 47 48 49 52 54 55 57 61 63 65 69 70 71
c140 69 0 2.22566e-19 $X=12.82 $Y=0.7
c141 38 0 1.88329e-19 $X=18.58 $Y=1.845
r142 66 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.38
+ $Y=1.91 $X2=15.38 $Y2=1.91
r143 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.38
+ $Y=1.57 $X2=15.38 $Y2=1.57
r144 63 73 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.38 $Y=1.825
+ $X2=15.38 $Y2=1.91
r145 63 65 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=15.38 $Y=1.825
+ $X2=15.38 $Y2=1.57
r146 59 61 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=15.135 $Y=2.695
+ $X2=15.135 $Y2=2.925
r147 58 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.755 $Y=2.61
+ $X2=13.67 $Y2=2.61
r148 57 59 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=14.97 $Y=2.61
+ $X2=15.135 $Y2=2.695
r149 57 58 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=14.97 $Y=2.61
+ $X2=13.755 $Y2=2.61
r150 56 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.755 $Y=1.91
+ $X2=13.67 $Y2=1.91
r151 55 73 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.215 $Y=1.91
+ $X2=15.38 $Y2=1.91
r152 55 56 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=15.215 $Y=1.91
+ $X2=13.755 $Y2=1.91
r153 54 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.67 $Y=2.525
+ $X2=13.67 $Y2=2.61
r154 53 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.67 $Y=1.995
+ $X2=13.67 $Y2=1.91
r155 53 54 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=13.67 $Y=1.995
+ $X2=13.67 $Y2=2.525
r156 52 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.67 $Y=1.825
+ $X2=13.67 $Y2=1.91
r157 51 52 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=13.67 $Y=0.785
+ $X2=13.67 $Y2=1.825
r158 50 69 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.985 $Y=0.7
+ $X2=12.82 $Y2=0.7
r159 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.585 $Y=0.7
+ $X2=13.67 $Y2=0.785
r160 49 50 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=13.585 $Y=0.7
+ $X2=12.985 $Y2=0.7
r161 47 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.585 $Y=2.61
+ $X2=13.67 $Y2=2.61
r162 47 48 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=13.585 $Y=2.61
+ $X2=12.845 $Y2=2.61
r163 41 43 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=12.68 $Y=2.84
+ $X2=12.68 $Y2=3.215
r164 39 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.68 $Y=2.695
+ $X2=12.845 $Y2=2.61
r165 39 41 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=12.68 $Y=2.695
+ $X2=12.68 $Y2=2.84
r166 34 35 5.9297 $w=5.69e-07 $l=7e-08 $layer=POLY_cond $X=16.285 $Y=1.745
+ $X2=16.355 $Y2=1.745
r167 33 66 48.1118 $w=7e-07 $l=6.55e-07 $layer=POLY_cond $X=16.035 $Y=1.745
+ $X2=15.38 $Y2=1.745
r168 33 34 19.0441 $w=7e-07 $l=2.5e-07 $layer=POLY_cond $X=16.035 $Y=1.745
+ $X2=16.285 $Y2=1.745
r169 29 38 20.4101 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=18.58 $Y=2.095
+ $X2=18.58 $Y2=1.845
r170 29 31 72.229 $w=5e-07 $l=6.75e-07 $layer=POLY_cond $X=18.58 $Y=2.095
+ $X2=18.58 $Y2=2.77
r171 25 38 20.4101 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=18.58 $Y=1.595
+ $X2=18.58 $Y2=1.845
r172 25 27 55.6431 $w=5e-07 $l=5.2e-07 $layer=POLY_cond $X=18.58 $Y=1.595
+ $X2=18.58 $Y2=1.075
r173 24 37 22.0092 $w=5.69e-07 $l=2.95804e-07 $layer=POLY_cond $X=17.48 $Y=1.845
+ $X2=17.23 $Y2=1.745
r174 23 38 5.30422 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=18.33 $Y=1.845
+ $X2=18.58 $Y2=1.845
r175 23 24 90.955 $w=5e-07 $l=8.5e-07 $layer=POLY_cond $X=18.33 $Y=1.845
+ $X2=17.48 $Y2=1.845
r176 20 37 5.89942 $w=5e-07 $l=3.5e-07 $layer=POLY_cond $X=17.23 $Y=2.095
+ $X2=17.23 $Y2=1.745
r177 20 22 83.868 $w=5e-07 $l=8.7e-07 $layer=POLY_cond $X=17.23 $Y=2.095
+ $X2=17.23 $Y2=2.965
r178 16 37 4.2355 $w=5.69e-07 $l=5e-08 $layer=POLY_cond $X=17.18 $Y=1.745
+ $X2=17.23 $Y2=1.745
r179 16 35 69.8858 $w=5.69e-07 $l=8.25e-07 $layer=POLY_cond $X=17.18 $Y=1.745
+ $X2=16.355 $Y2=1.745
r180 16 18 73.299 $w=5e-07 $l=6.85e-07 $layer=POLY_cond $X=17.18 $Y=1.595
+ $X2=17.18 $Y2=0.91
r181 13 35 5.89942 $w=5e-07 $l=3.5e-07 $layer=POLY_cond $X=16.355 $Y=2.095
+ $X2=16.355 $Y2=1.745
r182 13 15 31.812 $w=5e-07 $l=3.3e-07 $layer=POLY_cond $X=16.355 $Y=2.095
+ $X2=16.355 $Y2=2.425
r183 10 34 5.89942 $w=5e-07 $l=3.5e-07 $layer=POLY_cond $X=16.285 $Y=1.395
+ $X2=16.285 $Y2=1.745
r184 10 12 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=16.285 $Y=1.395
+ $X2=16.285 $Y2=1.075
r185 3 61 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=14.995
+ $Y=2.715 $X2=15.135 $Y2=2.925
r186 2 43 300 $w=1.7e-07 $l=5.80948e-07 $layer=licon1_PDIFF $count=2 $X=12.505
+ $Y=2.715 $X2=12.68 $Y2=3.215
r187 2 41 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=12.505
+ $Y=2.715 $X2=12.68 $Y2=2.84
r188 1 69 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=12.68
+ $Y=0.535 $X2=12.82 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%A_3609_173# 1 2 9 13 15 19 21 24 28
c41 19 0 1.88329e-19 $X=18.19 $Y=1.59
r42 22 28 131.082 $w=5e-07 $l=1.225e-06 $layer=POLY_cond $X=19.475 $Y=1.67
+ $X2=19.475 $Y2=2.895
r43 22 24 81.3245 $w=5e-07 $l=7.6e-07 $layer=POLY_cond $X=19.475 $Y=1.67
+ $X2=19.475 $Y2=0.91
r44 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=19.41
+ $Y=1.67 $X2=19.41 $Y2=1.67
r45 16 19 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.355 $Y=1.59
+ $X2=18.19 $Y2=1.59
r46 15 21 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.245 $Y=1.59
+ $X2=19.41 $Y2=1.59
r47 15 16 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=19.245 $Y=1.59
+ $X2=18.355 $Y2=1.59
r48 11 19 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.19 $Y=1.675
+ $X2=18.19 $Y2=1.59
r49 11 13 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=18.19 $Y=1.675
+ $X2=18.19 $Y2=2.52
r50 7 19 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.19 $Y=1.505
+ $X2=18.19 $Y2=1.59
r51 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=18.19 $Y=1.505
+ $X2=18.19 $Y2=1.075
r52 2 13 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=18.045
+ $Y=2.395 $X2=18.19 $Y2=2.52
r53 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=18.045
+ $Y=0.865 $X2=18.19 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%VPWR 1 2 3 4 5 6 7 8 25 28 37 48 55 69 73
+ 82 95 103
c118 103 0 3.3847e-20 $X=19.37 $Y=3.59
r119 101 103 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=18.65 $Y=3.63
+ $X2=19.37 $Y2=3.63
r120 100 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=19.37 $Y=3.59
+ $X2=19.37 $Y2=3.59
r121 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=18.65 $Y=3.59
+ $X2=18.65 $Y2=3.59
r122 98 100 4.10947 $w=9.48e-07 $l=3.2e-07 $layer=LI1_cond $X=19.01 $Y=3.27
+ $X2=19.01 $Y2=3.59
r123 95 98 9.63158 $w=9.48e-07 $l=7.5e-07 $layer=LI1_cond $X=19.01 $Y=2.52
+ $X2=19.01 $Y2=3.27
r124 92 101 0.604651 $w=3.7e-07 $l=1.575e-06 $layer=MET1_cond $X=17.075 $Y=3.63
+ $X2=18.65 $Y2=3.63
r125 90 92 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=16.355 $Y=3.63
+ $X2=17.075 $Y2=3.63
r126 89 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.075 $Y=3.59
+ $X2=17.075 $Y2=3.59
r127 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.355 $Y=3.59
+ $X2=16.355 $Y2=3.59
r128 87 89 0.256842 $w=9.48e-07 $l=2e-08 $layer=LI1_cond $X=16.715 $Y=3.57
+ $X2=16.715 $Y2=3.59
r129 85 87 10.4021 $w=9.48e-07 $l=8.1e-07 $layer=LI1_cond $X=16.715 $Y=2.76
+ $X2=16.715 $Y2=3.57
r130 82 85 5.13684 $w=9.48e-07 $l=4e-07 $layer=LI1_cond $X=16.715 $Y=2.36
+ $X2=16.715 $Y2=2.76
r131 79 90 0.775489 $w=3.7e-07 $l=2.02e-06 $layer=MET1_cond $X=14.335 $Y=3.63
+ $X2=16.355 $Y2=3.63
r132 77 79 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=13.615 $Y=3.63
+ $X2=14.335 $Y2=3.63
r133 76 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.335 $Y=3.59
+ $X2=14.335 $Y2=3.59
r134 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.615 $Y=3.59
+ $X2=13.615 $Y2=3.59
r135 73 76 7.76947 $w=9.48e-07 $l=6.05e-07 $layer=LI1_cond $X=13.975 $Y=2.985
+ $X2=13.975 $Y2=3.59
r136 70 77 0.700627 $w=3.7e-07 $l=1.825e-06 $layer=MET1_cond $X=11.79 $Y=3.63
+ $X2=13.615 $Y2=3.63
r137 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.79 $Y=3.59
+ $X2=11.79 $Y2=3.59
r138 65 70 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=11.07 $Y=3.63
+ $X2=11.79 $Y2=3.63
r139 64 69 20.4879 $w=4.03e-07 $l=7.2e-07 $layer=LI1_cond $X=11.07 $Y=3.552
+ $X2=11.79 $Y2=3.552
r140 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.07 $Y=3.59
+ $X2=11.07 $Y2=3.59
r141 59 61 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.73 $Y=3.63
+ $X2=9.45 $Y2=3.63
r142 58 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.45 $Y=3.59
+ $X2=9.45 $Y2=3.59
r143 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.73 $Y=3.59
+ $X2=8.73 $Y2=3.59
r144 55 58 6.80632 $w=9.48e-07 $l=5.3e-07 $layer=LI1_cond $X=9.09 $Y=3.06
+ $X2=9.09 $Y2=3.59
r145 52 59 1.13252 $w=3.7e-07 $l=2.95e-06 $layer=MET1_cond $X=5.78 $Y=3.63
+ $X2=8.73 $Y2=3.63
r146 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.78 $Y=3.59
+ $X2=5.78 $Y2=3.59
r147 48 51 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=5.78 $Y=2.565
+ $X2=5.78 $Y2=3.59
r148 45 52 0.598892 $w=3.7e-07 $l=1.56e-06 $layer=MET1_cond $X=4.22 $Y=3.63
+ $X2=5.78 $Y2=3.63
r149 43 45 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.5 $Y=3.63
+ $X2=4.22 $Y2=3.63
r150 42 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.22 $Y=3.59
+ $X2=4.22 $Y2=3.59
r151 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.5 $Y=3.59
+ $X2=3.5 $Y2=3.59
r152 40 42 1.64494 $w=8.88e-07 $l=1.2e-07 $layer=LI1_cond $X=3.86 $Y=3.47
+ $X2=3.86 $Y2=3.59
r153 37 40 6.85393 $w=8.88e-07 $l=5e-07 $layer=LI1_cond $X=3.86 $Y=2.97 $X2=3.86
+ $Y2=3.47
r154 34 43 0.777408 $w=3.7e-07 $l=2.025e-06 $layer=MET1_cond $X=1.475 $Y=3.63
+ $X2=3.5 $Y2=3.63
r155 32 34 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.755 $Y=3.63
+ $X2=1.475 $Y2=3.63
r156 31 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.475 $Y=3.59
+ $X2=1.475 $Y2=3.59
r157 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.755 $Y=3.59
+ $X2=0.755 $Y2=3.59
r158 28 31 6.87053 $w=9.48e-07 $l=5.35e-07 $layer=LI1_cond $X=1.115 $Y=3.055
+ $X2=1.115 $Y2=3.59
r159 25 65 0.380066 $w=3.7e-07 $l=9.9e-07 $layer=MET1_cond $X=10.08 $Y=3.63
+ $X2=11.07 $Y2=3.63
r160 25 61 0.24186 $w=3.7e-07 $l=6.3e-07 $layer=MET1_cond $X=10.08 $Y=3.63
+ $X2=9.45 $Y2=3.63
r161 8 98 600 $w=1.7e-07 $l=9.94359e-07 $layer=licon1_PDIFF $count=1 $X=18.83
+ $Y=2.395 $X2=19.085 $Y2=3.27
r162 8 95 300 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=2 $X=18.83
+ $Y=2.395 $X2=19.085 $Y2=2.52
r163 7 87 400 $w=1.7e-07 $l=1.4678e-06 $layer=licon1_PDIFF $count=1 $X=16.605
+ $Y=2.215 $X2=16.84 $Y2=3.57
r164 7 85 400 $w=1.7e-07 $l=6.51997e-07 $layer=licon1_PDIFF $count=1 $X=16.605
+ $Y=2.215 $X2=16.84 $Y2=2.76
r165 7 82 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=16.605
+ $Y=2.215 $X2=16.84 $Y2=2.36
r166 6 73 600 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=14.145
+ $Y=2.715 $X2=14.285 $Y2=2.985
r167 5 64 600 $w=1.7e-07 $l=8.47968e-07 $layer=licon1_PDIFF $count=1 $X=10.9
+ $Y=2.78 $X2=11.155 $Y2=3.51
r168 4 55 600 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=9.26
+ $Y=2.78 $X2=9.4 $Y2=3.06
r169 3 48 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=5.635
+ $Y=2.44 $X2=5.78 $Y2=2.565
r170 2 40 600 $w=1.7e-07 $l=7.62398e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=2.845 $X2=4.22 $Y2=3.47
r171 2 37 600 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=2.845 $X2=4.22 $Y2=2.97
r172 1 28 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=2.845 $X2=1.075 $Y2=3.055
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%A_485_569# 1 2 3 4 13 15 18 20 21 24 25 26
+ 28 29 30 32 33 34 37 41 44 45 51 55 56 57
c143 55 0 4.65845e-20 $X=3.185 $Y=2.54
r144 56 57 109.604 $w=1.68e-07 $l=1.68e-06 $layer=LI1_cond $X=6.925 $Y=1.06
+ $X2=6.925 $Y2=2.74
r145 51 53 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=0.745
+ $X2=2.59 $Y2=0.83
r146 45 48 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=2.97
+ $X2=2.565 $Y2=3.055
r147 42 44 10.515 $w=4.53e-07 $l=4e-07 $layer=LI1_cond $X=7.067 $Y=3.39
+ $X2=7.067 $Y2=2.99
r148 41 57 10.8817 $w=4.53e-07 $l=2.27e-07 $layer=LI1_cond $X=7.067 $Y=2.967
+ $X2=7.067 $Y2=2.74
r149 41 44 0.604611 $w=4.53e-07 $l=2.3e-08 $layer=LI1_cond $X=7.067 $Y=2.967
+ $X2=7.067 $Y2=2.99
r150 35 56 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.885 $Y=0.935
+ $X2=6.885 $Y2=1.06
r151 35 37 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=6.885 $Y=0.935
+ $X2=6.885 $Y2=0.835
r152 33 42 8.8478 $w=1.7e-07 $l=2.66128e-07 $layer=LI1_cond $X=6.84 $Y=3.475
+ $X2=7.067 $Y2=3.39
r153 33 34 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.84 $Y=3.475
+ $X2=6.215 $Y2=3.475
r154 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.13 $Y=3.39
+ $X2=6.215 $Y2=3.475
r155 31 32 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=6.13 $Y=2.22
+ $X2=6.13 $Y2=3.39
r156 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.045 $Y=2.135
+ $X2=6.13 $Y2=2.22
r157 29 30 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.045 $Y=2.135
+ $X2=5.515 $Y2=2.135
r158 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.43 $Y=2.22
+ $X2=5.515 $Y2=2.135
r159 27 28 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=5.43 $Y=2.22
+ $X2=5.43 $Y2=3.635
r160 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.345 $Y=3.72
+ $X2=5.43 $Y2=3.635
r161 25 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.345 $Y=3.72
+ $X2=4.655 $Y2=3.72
r162 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.57 $Y=3.635
+ $X2=4.655 $Y2=3.72
r163 23 24 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=4.57 $Y=2.625
+ $X2=4.57 $Y2=3.635
r164 22 55 1.34256 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.305 $Y=2.54
+ $X2=3.185 $Y2=2.54
r165 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.485 $Y=2.54
+ $X2=4.57 $Y2=2.625
r166 21 22 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=4.485 $Y=2.54
+ $X2=3.305 $Y2=2.54
r167 20 55 5.16603 $w=1.7e-07 $l=1.00995e-07 $layer=LI1_cond $X=3.22 $Y=2.455
+ $X2=3.185 $Y2=2.54
r168 19 20 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=3.22 $Y=0.915
+ $X2=3.22 $Y2=2.455
r169 17 55 5.16603 $w=1.7e-07 $l=1.00995e-07 $layer=LI1_cond $X=3.15 $Y=2.625
+ $X2=3.185 $Y2=2.54
r170 17 18 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.15 $Y=2.625
+ $X2=3.15 $Y2=2.885
r171 16 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=0.83
+ $X2=2.59 $Y2=0.83
r172 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.135 $Y=0.83
+ $X2=3.22 $Y2=0.915
r173 15 16 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.135 $Y=0.83
+ $X2=2.755 $Y2=0.83
r174 14 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=2.97
+ $X2=2.565 $Y2=2.97
r175 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.065 $Y=2.97
+ $X2=3.15 $Y2=2.885
r176 13 14 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.065 $Y=2.97
+ $X2=2.73 $Y2=2.97
r177 4 44 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=6.985
+ $Y=2.78 $X2=7.13 $Y2=2.99
r178 3 48 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=2.845 $X2=2.565 $Y2=3.055
r179 2 37 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=6.78
+ $Y=0.6 $X2=6.925 $Y2=0.835
r180 1 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.45
+ $Y=0.535 $X2=2.59 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%Q_N 1 2 7 8 9 10 11 12 13 22
r18 13 41 12.8892 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=17.595 $Y=3.145
+ $X2=17.595 $Y2=3.57
r19 12 13 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=17.595 $Y=2.775
+ $X2=17.595 $Y2=3.145
r20 11 12 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=17.595 $Y=2.405
+ $X2=17.595 $Y2=2.775
r21 11 33 1.36474 $w=3.78e-07 $l=4.5e-08 $layer=LI1_cond $X=17.595 $Y=2.405
+ $X2=17.595 $Y2=2.36
r22 10 33 9.85642 $w=3.78e-07 $l=3.25e-07 $layer=LI1_cond $X=17.595 $Y=2.035
+ $X2=17.595 $Y2=2.36
r23 9 10 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=17.595 $Y=1.665
+ $X2=17.595 $Y2=2.035
r24 8 9 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=17.595 $Y=1.295
+ $X2=17.595 $Y2=1.665
r25 7 8 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=17.595 $Y=0.925
+ $X2=17.595 $Y2=1.295
r26 7 22 8.03677 $w=3.78e-07 $l=2.65e-07 $layer=LI1_cond $X=17.595 $Y=0.925
+ $X2=17.595 $Y2=0.66
r27 2 41 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=17.48
+ $Y=2.215 $X2=17.62 $Y2=3.57
r28 2 33 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=17.48
+ $Y=2.215 $X2=17.62 $Y2=2.36
r29 1 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=17.43
+ $Y=0.535 $X2=17.57 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%Q 1 2 7 8 9 10 11 12 13 25 47 50
r16 50 51 2.86126 $w=3.33e-07 $l=5e-08 $layer=LI1_cond $X=19.867 $Y=2.405
+ $X2=19.867 $Y2=2.355
r17 47 48 2.17324 $w=3.33e-07 $l=3e-08 $layer=LI1_cond $X=19.867 $Y=1.295
+ $X2=19.867 $Y2=1.325
r18 37 54 0.0688026 $w=3.33e-07 $l=2e-09 $layer=LI1_cond $X=19.867 $Y=2.522
+ $X2=19.867 $Y2=2.52
r19 13 43 4.30016 $w=3.33e-07 $l=1.25e-07 $layer=LI1_cond $X=19.867 $Y=3.145
+ $X2=19.867 $Y2=3.27
r20 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=19.867 $Y=2.775
+ $X2=19.867 $Y2=3.145
r21 12 37 8.70352 $w=3.33e-07 $l=2.53e-07 $layer=LI1_cond $X=19.867 $Y=2.775
+ $X2=19.867 $Y2=2.522
r22 11 54 3.37133 $w=3.33e-07 $l=9.8e-08 $layer=LI1_cond $X=19.867 $Y=2.422
+ $X2=19.867 $Y2=2.52
r23 11 50 0.584822 $w=3.33e-07 $l=1.7e-08 $layer=LI1_cond $X=19.867 $Y=2.422
+ $X2=19.867 $Y2=2.405
r24 11 51 0.901912 $w=2.28e-07 $l=1.8e-08 $layer=LI1_cond $X=19.92 $Y=2.337
+ $X2=19.92 $Y2=2.355
r25 10 11 15.1321 $w=2.28e-07 $l=3.02e-07 $layer=LI1_cond $X=19.92 $Y=2.035
+ $X2=19.92 $Y2=2.337
r26 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=19.92 $Y=1.665
+ $X2=19.92 $Y2=2.035
r27 8 47 0.963236 $w=3.33e-07 $l=2.8e-08 $layer=LI1_cond $X=19.867 $Y=1.267
+ $X2=19.867 $Y2=1.295
r28 8 23 3.74974 $w=3.33e-07 $l=1.09e-07 $layer=LI1_cond $X=19.867 $Y=1.267
+ $X2=19.867 $Y2=1.158
r29 8 9 15.6832 $w=2.28e-07 $l=3.13e-07 $layer=LI1_cond $X=19.92 $Y=1.352
+ $X2=19.92 $Y2=1.665
r30 8 48 1.35287 $w=2.28e-07 $l=2.7e-08 $layer=LI1_cond $X=19.92 $Y=1.352
+ $X2=19.92 $Y2=1.325
r31 7 23 8.0155 $w=3.33e-07 $l=2.33e-07 $layer=LI1_cond $X=19.867 $Y=0.925
+ $X2=19.867 $Y2=1.158
r32 7 25 9.11634 $w=3.33e-07 $l=2.65e-07 $layer=LI1_cond $X=19.867 $Y=0.925
+ $X2=19.867 $Y2=0.66
r33 2 54 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=19.725
+ $Y=2.395 $X2=19.865 $Y2=2.52
r34 2 43 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=19.725
+ $Y=2.395 $X2=19.865 $Y2=3.27
r35 1 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=19.725
+ $Y=0.535 $X2=19.865 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSBP_1%VGND 1 2 3 4 5 6 7 8 25 28 37 46 53 62 71
+ 80 91 95
r133 97 99 6.42105 $w=9.48e-07 $l=5e-07 $layer=LI1_cond $X=19.01 $Y=0.66
+ $X2=19.01 $Y2=1.16
r134 92 95 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=18.65 $Y=0.44
+ $X2=19.37 $Y2=0.44
r135 91 97 2.31158 $w=9.48e-07 $l=1.8e-07 $layer=LI1_cond $X=19.01 $Y=0.48
+ $X2=19.01 $Y2=0.66
r136 91 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=19.37 $Y=0.48
+ $X2=19.37 $Y2=0.48
r137 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=18.65 $Y=0.48
+ $X2=18.65 $Y2=0.48
r138 86 88 6.42105 $w=9.48e-07 $l=5e-07 $layer=LI1_cond $X=16.715 $Y=0.66
+ $X2=16.715 $Y2=1.16
r139 84 92 0.604651 $w=3.7e-07 $l=1.575e-06 $layer=MET1_cond $X=17.075 $Y=0.44
+ $X2=18.65 $Y2=0.44
r140 81 84 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=16.355 $Y=0.44
+ $X2=17.075 $Y2=0.44
r141 80 86 2.31158 $w=9.48e-07 $l=1.8e-07 $layer=LI1_cond $X=16.715 $Y=0.48
+ $X2=16.715 $Y2=0.66
r142 80 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.075 $Y=0.48
+ $X2=17.075 $Y2=0.48
r143 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.355 $Y=0.48
+ $X2=16.355 $Y2=0.48
r144 75 81 0.449169 $w=3.7e-07 $l=1.17e-06 $layer=MET1_cond $X=15.185 $Y=0.44
+ $X2=16.355 $Y2=0.44
r145 72 75 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=14.465 $Y=0.44
+ $X2=15.185 $Y2=0.44
r146 71 77 7.64105 $w=9.48e-07 $l=5.95e-07 $layer=LI1_cond $X=14.825 $Y=0.48
+ $X2=14.825 $Y2=1.075
r147 71 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.185 $Y=0.48
+ $X2=15.185 $Y2=0.48
r148 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.465 $Y=0.48
+ $X2=14.465 $Y2=0.48
r149 66 72 1.18435 $w=3.7e-07 $l=3.085e-06 $layer=MET1_cond $X=11.38 $Y=0.44
+ $X2=14.465 $Y2=0.44
r150 63 66 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.66 $Y=0.44
+ $X2=11.38 $Y2=0.44
r151 62 68 4.23789 $w=9.48e-07 $l=3.3e-07 $layer=LI1_cond $X=11.02 $Y=0.48
+ $X2=11.02 $Y2=0.81
r152 62 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.38 $Y=0.48
+ $X2=11.38 $Y2=0.48
r153 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.66 $Y=0.48
+ $X2=10.66 $Y2=0.48
r154 54 57 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.525 $Y=0.44
+ $X2=9.245 $Y2=0.44
r155 53 59 4.23789 $w=9.48e-07 $l=3.3e-07 $layer=LI1_cond $X=8.885 $Y=0.48
+ $X2=8.885 $Y2=0.81
r156 53 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.245 $Y=0.48
+ $X2=9.245 $Y2=0.48
r157 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.525 $Y=0.48
+ $X2=8.525 $Y2=0.48
r158 47 54 1.02887 $w=3.7e-07 $l=2.68e-06 $layer=MET1_cond $X=5.845 $Y=0.44
+ $X2=8.525 $Y2=0.44
r159 46 50 6.28448 $w=5.88e-07 $l=3.1e-07 $layer=LI1_cond $X=5.665 $Y=0.48
+ $X2=5.665 $Y2=0.79
r160 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.845 $Y=0.48
+ $X2=5.845 $Y2=0.48
r161 41 47 0.449169 $w=3.7e-07 $l=1.17e-06 $layer=MET1_cond $X=4.675 $Y=0.44
+ $X2=5.845 $Y2=0.44
r162 38 41 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.955 $Y=0.44
+ $X2=4.675 $Y2=0.44
r163 37 43 3.63258 $w=8.88e-07 $l=2.65e-07 $layer=LI1_cond $X=4.315 $Y=0.48
+ $X2=4.315 $Y2=0.745
r164 37 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.675 $Y=0.48
+ $X2=4.675 $Y2=0.48
r165 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.955 $Y=0.48
+ $X2=3.955 $Y2=0.48
r166 32 38 0.942488 $w=3.7e-07 $l=2.455e-06 $layer=MET1_cond $X=1.5 $Y=0.44
+ $X2=3.955 $Y2=0.44
r167 29 32 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.78 $Y=0.44
+ $X2=1.5 $Y2=0.44
r168 28 34 3.40316 $w=9.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.14 $Y=0.48
+ $X2=1.14 $Y2=0.745
r169 28 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.5 $Y=0.48
+ $X2=1.5 $Y2=0.48
r170 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.78 $Y=0.48
+ $X2=0.78 $Y2=0.48
r171 25 63 0.222665 $w=3.7e-07 $l=5.8e-07 $layer=MET1_cond $X=10.08 $Y=0.44
+ $X2=10.66 $Y2=0.44
r172 25 57 0.320561 $w=3.7e-07 $l=8.35e-07 $layer=MET1_cond $X=10.08 $Y=0.44
+ $X2=9.245 $Y2=0.44
r173 8 99 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=18.83
+ $Y=0.865 $X2=19.085 $Y2=1.16
r174 8 97 182 $w=1.7e-07 $l=3.42491e-07 $layer=licon1_NDIFF $count=1 $X=18.83
+ $Y=0.865 $X2=19.085 $Y2=0.66
r175 7 88 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=16.535
+ $Y=0.865 $X2=16.79 $Y2=1.16
r176 7 86 182 $w=1.7e-07 $l=3.42491e-07 $layer=licon1_NDIFF $count=1 $X=16.535
+ $Y=0.865 $X2=16.79 $Y2=0.66
r177 6 77 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=14.995
+ $Y=0.865 $X2=15.135 $Y2=1.075
r178 5 68 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=11.095
+ $Y=0.535 $X2=11.33 $Y2=0.81
r179 4 59 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.055
+ $Y=0.6 $X2=9.195 $Y2=0.81
r180 3 50 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.45
+ $Y=0.58 $X2=5.575 $Y2=0.79
r181 2 43 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.94
+ $Y=0.535 $X2=4.08 $Y2=0.745
r182 1 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.535 $X2=1.1 $Y2=0.745
.ends

