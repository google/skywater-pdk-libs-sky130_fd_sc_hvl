* File: sky130_fd_sc_hvl__buf_16.spice
* Created: Wed Sep  2 09:03:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__buf_16.pex.spice"
.subckt sky130_fd_sc_hvl__buf_16  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_183_141#_M1006_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250016 A=0.375 P=2.5 MULT=1
MM1016 N_VGND_M1016_d N_A_M1016_g N_A_183_141#_M1006_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250001
+ SB=250016 A=0.375 P=2.5 MULT=1
MM1019 N_VGND_M1016_d N_A_M1019_g N_A_183_141#_M1019_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250002
+ SB=250015 A=0.375 P=2.5 MULT=1
MM1026 N_VGND_M1026_d N_A_M1026_g N_A_183_141#_M1019_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250002
+ SB=250014 A=0.375 P=2.5 MULT=1
MM1040 N_VGND_M1026_d N_A_M1040_g N_A_183_141#_M1040_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250003
+ SB=250013 A=0.375 P=2.5 MULT=1
MM1043 N_VGND_M1043_d N_A_M1043_g N_A_183_141#_M1040_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250004
+ SB=250012 A=0.375 P=2.5 MULT=1
MM1002 N_VGND_M1043_d N_A_183_141#_M1002_g N_X_M1002_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250005
+ SB=250012 A=0.375 P=2.5 MULT=1
MM1004 N_VGND_M1004_d N_A_183_141#_M1004_g N_X_M1002_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250005
+ SB=250011 A=0.375 P=2.5 MULT=1
MM1007 N_VGND_M1004_d N_A_183_141#_M1007_g N_X_M1007_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250006
+ SB=250010 A=0.375 P=2.5 MULT=1
MM1009 N_VGND_M1009_d N_A_183_141#_M1009_g N_X_M1007_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250007
+ SB=250009 A=0.375 P=2.5 MULT=1
MM1014 N_VGND_M1009_d N_A_183_141#_M1014_g N_X_M1014_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250008
+ SB=250009 A=0.375 P=2.5 MULT=1
MM1017 N_VGND_M1017_d N_A_183_141#_M1017_g N_X_M1014_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250009
+ SB=250008 A=0.375 P=2.5 MULT=1
MM1020 N_VGND_M1017_d N_A_183_141#_M1020_g N_X_M1020_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250009
+ SB=250007 A=0.375 P=2.5 MULT=1
MM1024 N_VGND_M1024_d N_A_183_141#_M1024_g N_X_M1020_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250010
+ SB=250006 A=0.375 P=2.5 MULT=1
MM1027 N_VGND_M1024_d N_A_183_141#_M1027_g N_X_M1027_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250011
+ SB=250005 A=0.375 P=2.5 MULT=1
MM1028 N_VGND_M1028_d N_A_183_141#_M1028_g N_X_M1027_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250012
+ SB=250005 A=0.375 P=2.5 MULT=1
MM1030 N_VGND_M1028_d N_A_183_141#_M1030_g N_X_M1030_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250012
+ SB=250004 A=0.375 P=2.5 MULT=1
MM1032 N_VGND_M1032_d N_A_183_141#_M1032_g N_X_M1030_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250013
+ SB=250003 A=0.375 P=2.5 MULT=1
MM1034 N_VGND_M1032_d N_A_183_141#_M1034_g N_X_M1034_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250014
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1035 N_VGND_M1035_d N_A_183_141#_M1035_g N_X_M1034_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250015
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1037 N_VGND_M1035_d N_A_183_141#_M1037_g N_X_M1037_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250016
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1041 N_VGND_M1041_d N_A_183_141#_M1041_g N_X_M1037_s N_VNB_M1006_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250016
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_183_141#_M1000_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250016 A=0.75 P=4 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_A_183_141#_M1000_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001 SB=250016
+ A=0.75 P=4 MULT=1
MM1011 N_VPWR_M1005_d N_A_M1011_g N_A_183_141#_M1011_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002 SB=250015
+ A=0.75 P=4 MULT=1
MM1023 N_VPWR_M1023_d N_A_M1023_g N_A_183_141#_M1011_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002 SB=250014
+ A=0.75 P=4 MULT=1
MM1029 N_VPWR_M1023_d N_A_M1029_g N_A_183_141#_M1029_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250003 SB=250013
+ A=0.75 P=4 MULT=1
MM1036 N_VPWR_M1036_d N_A_M1036_g N_A_183_141#_M1029_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250004 SB=250012
+ A=0.75 P=4 MULT=1
MM1001 N_X_M1001_d N_A_183_141#_M1001_g N_VPWR_M1036_d N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250005 SB=250012
+ A=0.75 P=4 MULT=1
MM1003 N_X_M1001_d N_A_183_141#_M1003_g N_VPWR_M1003_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250005 SB=250011
+ A=0.75 P=4 MULT=1
MM1008 N_X_M1008_d N_A_183_141#_M1008_g N_VPWR_M1003_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250006 SB=250010
+ A=0.75 P=4 MULT=1
MM1010 N_X_M1008_d N_A_183_141#_M1010_g N_VPWR_M1010_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250007 SB=250009
+ A=0.75 P=4 MULT=1
MM1012 N_X_M1012_d N_A_183_141#_M1012_g N_VPWR_M1010_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250008 SB=250009
+ A=0.75 P=4 MULT=1
MM1013 N_X_M1012_d N_A_183_141#_M1013_g N_VPWR_M1013_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250009 SB=250008
+ A=0.75 P=4 MULT=1
MM1015 N_X_M1015_d N_A_183_141#_M1015_g N_VPWR_M1013_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250009 SB=250007
+ A=0.75 P=4 MULT=1
MM1018 N_X_M1015_d N_A_183_141#_M1018_g N_VPWR_M1018_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250010 SB=250006
+ A=0.75 P=4 MULT=1
MM1021 N_X_M1021_d N_A_183_141#_M1021_g N_VPWR_M1018_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250011 SB=250005
+ A=0.75 P=4 MULT=1
MM1022 N_X_M1021_d N_A_183_141#_M1022_g N_VPWR_M1022_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250012 SB=250005
+ A=0.75 P=4 MULT=1
MM1025 N_X_M1025_d N_A_183_141#_M1025_g N_VPWR_M1022_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250012 SB=250004
+ A=0.75 P=4 MULT=1
MM1031 N_X_M1025_d N_A_183_141#_M1031_g N_VPWR_M1031_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250013 SB=250003
+ A=0.75 P=4 MULT=1
MM1033 N_X_M1033_d N_A_183_141#_M1033_g N_VPWR_M1031_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250014 SB=250002
+ A=0.75 P=4 MULT=1
MM1038 N_X_M1033_d N_A_183_141#_M1038_g N_VPWR_M1038_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250015 SB=250002
+ A=0.75 P=4 MULT=1
MM1039 N_X_M1039_d N_A_183_141#_M1039_g N_VPWR_M1038_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250016 SB=250001
+ A=0.75 P=4 MULT=1
MM1042 N_X_M1039_d N_A_183_141#_M1042_g N_VPWR_M1042_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 M=1 R=3 SA=250016
+ SB=250000 A=0.75 P=4 MULT=1
DX44_noxref N_VNB_M1006_b N_VPB_M1000_b NWDIODE A=47.892 P=42.04
*
.include "sky130_fd_sc_hvl__buf_16.pxi.spice"
*
.ends
*
*
