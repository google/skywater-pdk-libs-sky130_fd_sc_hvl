* File: sky130_fd_sc_hvl__dlxtp_1.pxi.spice
* Created: Fri Aug 28 09:35:18 2020
* 
x_PM_SKY130_FD_SC_HVL__DLXTP_1%VNB N_VNB_M1010_b VNB N_VNB_c_3_p VNB
+ PM_SKY130_FD_SC_HVL__DLXTP_1%VNB
x_PM_SKY130_FD_SC_HVL__DLXTP_1%VPB N_VPB_M1005_b VPB N_VPB_c_71_p VPB
+ PM_SKY130_FD_SC_HVL__DLXTP_1%VPB
x_PM_SKY130_FD_SC_HVL__DLXTP_1%GATE N_GATE_M1005_g N_GATE_M1010_g GATE
+ N_GATE_c_140_n PM_SKY130_FD_SC_HVL__DLXTP_1%GATE
x_PM_SKY130_FD_SC_HVL__DLXTP_1%A_30_443# N_A_30_443#_M1010_s N_A_30_443#_M1005_s
+ N_A_30_443#_M1000_g N_A_30_443#_M1011_g N_A_30_443#_c_169_n
+ N_A_30_443#_c_178_n N_A_30_443#_c_179_n N_A_30_443#_c_203_n
+ N_A_30_443#_c_170_n N_A_30_443#_c_208_n N_A_30_443#_c_181_n
+ N_A_30_443#_c_214_p N_A_30_443#_c_182_n N_A_30_443#_c_185_n
+ N_A_30_443#_c_226_p N_A_30_443#_c_217_p N_A_30_443#_c_187_n
+ N_A_30_443#_c_171_n N_A_30_443#_c_172_n N_A_30_443#_c_189_n
+ N_A_30_443#_c_244_p N_A_30_443#_c_190_n N_A_30_443#_M1006_g
+ N_A_30_443#_M1007_g PM_SKY130_FD_SC_HVL__DLXTP_1%A_30_443#
x_PM_SKY130_FD_SC_HVL__DLXTP_1%D N_D_M1004_g N_D_c_313_n N_D_M1013_g N_D_c_317_n
+ D N_D_c_311_n N_D_c_312_n PM_SKY130_FD_SC_HVL__DLXTP_1%D
x_PM_SKY130_FD_SC_HVL__DLXTP_1%A_384_107# N_A_384_107#_M1000_d
+ N_A_384_107#_M1011_d N_A_384_107#_M1015_g N_A_384_107#_c_359_n
+ N_A_384_107#_c_367_n N_A_384_107#_c_368_n N_A_384_107#_c_369_n
+ N_A_384_107#_M1014_g N_A_384_107#_c_360_n N_A_384_107#_c_362_n
+ N_A_384_107#_c_373_n N_A_384_107#_c_363_n N_A_384_107#_c_364_n
+ N_A_384_107#_c_414_n N_A_384_107#_c_365_n
+ PM_SKY130_FD_SC_HVL__DLXTP_1%A_384_107#
x_PM_SKY130_FD_SC_HVL__DLXTP_1%A_1004_81# N_A_1004_81#_M1003_s
+ N_A_1004_81#_M1008_s N_A_1004_81#_c_455_n N_A_1004_81#_M1012_g
+ N_A_1004_81#_c_486_p N_A_1004_81#_c_487_p N_A_1004_81#_c_457_n
+ N_A_1004_81#_c_458_n N_A_1004_81#_c_459_n N_A_1004_81#_c_463_n
+ N_A_1004_81#_c_460_n N_A_1004_81#_c_464_n N_A_1004_81#_c_461_n
+ N_A_1004_81#_c_467_n N_A_1004_81#_c_462_n N_A_1004_81#_M1001_g
+ PM_SKY130_FD_SC_HVL__DLXTP_1%A_1004_81#
x_PM_SKY130_FD_SC_HVL__DLXTP_1%A_806_107# N_A_806_107#_M1015_d
+ N_A_806_107#_M1006_d N_A_806_107#_M1008_g N_A_806_107#_M1003_g
+ N_A_806_107#_M1002_g N_A_806_107#_M1009_g N_A_806_107#_c_541_n
+ N_A_806_107#_c_542_n N_A_806_107#_c_530_n N_A_806_107#_c_545_n
+ N_A_806_107#_c_531_n N_A_806_107#_c_546_n N_A_806_107#_c_532_n
+ N_A_806_107#_c_534_n N_A_806_107#_c_591_n N_A_806_107#_c_535_n
+ N_A_806_107#_c_536_n PM_SKY130_FD_SC_HVL__DLXTP_1%A_806_107#
x_PM_SKY130_FD_SC_HVL__DLXTP_1%VPWR N_VPWR_M1005_d N_VPWR_M1013_s N_VPWR_M1001_d
+ N_VPWR_M1008_d VPWR N_VPWR_c_633_n N_VPWR_c_636_n N_VPWR_c_639_n
+ N_VPWR_c_642_n N_VPWR_c_645_n PM_SKY130_FD_SC_HVL__DLXTP_1%VPWR
x_PM_SKY130_FD_SC_HVL__DLXTP_1%A_650_107# N_A_650_107#_M1004_d
+ N_A_650_107#_M1013_d N_A_650_107#_c_687_n N_A_650_107#_c_688_n
+ N_A_650_107#_c_692_n N_A_650_107#_c_700_n N_A_650_107#_c_693_n
+ N_A_650_107#_c_694_n N_A_650_107#_c_690_n N_A_650_107#_c_691_n
+ N_A_650_107#_c_696_n PM_SKY130_FD_SC_HVL__DLXTP_1%A_650_107#
x_PM_SKY130_FD_SC_HVL__DLXTP_1%Q N_Q_M1009_d N_Q_M1002_d Q Q N_Q_c_751_n
+ PM_SKY130_FD_SC_HVL__DLXTP_1%Q
x_PM_SKY130_FD_SC_HVL__DLXTP_1%VGND N_VGND_M1010_d N_VGND_M1004_s N_VGND_M1012_d
+ N_VGND_M1003_d VGND N_VGND_c_766_n N_VGND_c_768_n N_VGND_c_770_n
+ N_VGND_c_772_n N_VGND_c_774_n PM_SKY130_FD_SC_HVL__DLXTP_1%VGND
cc_1 N_VNB_M1010_b N_GATE_M1005_g 0.00826652f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=2.59
cc_2 N_VNB_M1010_b N_GATE_M1010_g 0.0467682f $X=-0.33 $Y=-0.265 $X2=0.89
+ $Y2=0.745
cc_3 N_VNB_c_3_p N_GATE_M1010_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.89 $Y2=0.745
cc_4 N_VNB_M1010_b N_GATE_c_140_n 0.0991461f $X=-0.33 $Y=-0.265 $X2=0.705
+ $Y2=1.28
cc_5 N_VNB_M1010_b N_A_30_443#_M1000_g 0.0681875f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.21
cc_6 N_VNB_c_3_p N_A_30_443#_M1000_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.635 $Y2=1.21
cc_7 N_VNB_M1010_b N_A_30_443#_c_169_n 0.0467693f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_8 N_VNB_M1010_b N_A_30_443#_c_170_n 0.0646286f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_M1010_b N_A_30_443#_c_171_n 0.00156806f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_10 N_VNB_M1010_b N_A_30_443#_c_172_n 0.0450392f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_c_3_p N_A_30_443#_c_172_n 0.00135547f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_12 N_VNB_M1010_b N_A_30_443#_M1007_g 0.116159f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_13 N_VNB_c_3_p N_A_30_443#_M1007_g 0.0023273f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_14 N_VNB_M1010_b N_D_M1004_g 0.118641f $X=-0.33 $Y=-0.265 $X2=0.665 $Y2=2.59
cc_15 N_VNB_c_3_p N_D_M1004_g 0.00119158f $X=0.24 $Y=0 $X2=0.665 $Y2=2.59
cc_16 N_VNB_M1010_b N_D_c_311_n 0.0135335f $X=-0.33 $Y=-0.265 $X2=0.777
+ $Y2=1.805
cc_17 N_VNB_M1010_b N_D_c_312_n 0.0030442f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_18 N_VNB_M1010_b N_A_384_107#_M1015_g 0.0728286f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.21
cc_19 N_VNB_c_3_p N_A_384_107#_M1015_g 0.0023273f $X=0.24 $Y=0 $X2=0.635
+ $Y2=1.21
cc_20 N_VNB_M1010_b N_A_384_107#_c_359_n 0.0247731f $X=-0.33 $Y=-0.265 $X2=0.705
+ $Y2=1.28
cc_21 N_VNB_M1010_b N_A_384_107#_c_360_n 0.0244242f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_22 N_VNB_c_3_p N_A_384_107#_c_360_n 5.64934e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_23 N_VNB_M1010_b N_A_384_107#_c_362_n 0.0286877f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_24 N_VNB_M1010_b N_A_384_107#_c_363_n 0.00433715f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_25 N_VNB_M1010_b N_A_384_107#_c_364_n 0.00343325f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_26 N_VNB_M1010_b N_A_384_107#_c_365_n 0.0246928f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_27 N_VNB_M1010_b N_A_1004_81#_c_455_n 0.0445791f $X=-0.33 $Y=-0.265 $X2=0.89
+ $Y2=0.745
cc_28 N_VNB_c_3_p N_A_1004_81#_c_455_n 0.00116831f $X=0.24 $Y=0 $X2=0.89
+ $Y2=0.745
cc_29 N_VNB_M1010_b N_A_1004_81#_c_457_n 0.0724593f $X=-0.33 $Y=-0.265 $X2=0.705
+ $Y2=1.28
cc_30 N_VNB_M1010_b N_A_1004_81#_c_458_n 0.0108041f $X=-0.33 $Y=-0.265 $X2=0.777
+ $Y2=1.805
cc_31 N_VNB_M1010_b N_A_1004_81#_c_459_n 0.0103809f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_32 N_VNB_M1010_b N_A_1004_81#_c_460_n 0.00338411f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_33 N_VNB_M1010_b N_A_1004_81#_c_461_n 0.0338447f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_M1010_b N_A_1004_81#_c_462_n 0.00369881f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_35 N_VNB_M1010_b N_A_806_107#_M1003_g 0.0464881f $X=-0.33 $Y=-0.265 $X2=0.705
+ $Y2=1.28
cc_36 N_VNB_M1010_b N_A_806_107#_M1009_g 0.0677643f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_37 N_VNB_c_3_p N_A_806_107#_M1009_g 0.00112176f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_38 N_VNB_M1010_b N_A_806_107#_c_530_n 0.00710823f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_39 N_VNB_M1010_b N_A_806_107#_c_531_n 0.00871571f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_M1010_b N_A_806_107#_c_532_n 0.0109104f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_41 N_VNB_c_3_p N_A_806_107#_c_532_n 8.65969e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_42 N_VNB_M1010_b N_A_806_107#_c_534_n 4.78778e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_M1010_b N_A_806_107#_c_535_n 0.00802934f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_44 N_VNB_M1010_b N_A_806_107#_c_536_n 0.0845961f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_45 N_VNB_M1010_b N_A_650_107#_c_687_n 0.0061186f $X=-0.33 $Y=-0.265 $X2=0.89
+ $Y2=0.745
cc_46 N_VNB_M1010_b N_A_650_107#_c_688_n 0.0109585f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.21
cc_47 N_VNB_c_3_p N_A_650_107#_c_688_n 8.6949e-19 $X=0.24 $Y=0 $X2=0.635
+ $Y2=1.21
cc_48 N_VNB_M1010_b N_A_650_107#_c_690_n 0.00316667f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_49 N_VNB_M1010_b N_A_650_107#_c_691_n 0.0106031f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_M1010_b N_Q_c_751_n 0.0638623f $X=-0.33 $Y=-0.265 $X2=0.705 $Y2=1.28
cc_51 N_VNB_c_3_p N_Q_c_751_n 8.87563e-19 $X=0.24 $Y=0 $X2=0.705 $Y2=1.28
cc_52 N_VNB_M1010_b N_VGND_c_766_n 0.0580926f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_53 N_VNB_c_3_p N_VGND_c_766_n 0.00269373f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_54 N_VNB_M1010_b N_VGND_c_768_n 0.0406436f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_55 N_VNB_c_3_p N_VGND_c_768_n 0.00167165f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_56 N_VNB_M1010_b N_VGND_c_770_n 0.0418101f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_57 N_VNB_c_3_p N_VGND_c_770_n 0.00167538f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_58 N_VNB_M1010_b N_VGND_c_772_n 0.0578394f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_59 N_VNB_c_3_p N_VGND_c_772_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_60 N_VNB_M1010_b N_VGND_c_774_n 0.140178f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_61 N_VNB_c_3_p N_VGND_c_774_n 0.872906f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_62 N_VPB_M1005_b N_GATE_M1005_g 0.0659414f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=2.59
cc_63 N_VPB_M1005_b N_A_30_443#_M1011_g 0.0482669f $X=-0.33 $Y=1.885 $X2=0.705
+ $Y2=1.28
cc_64 N_VPB_M1005_b N_A_30_443#_c_169_n 9.52481e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_65 N_VPB_M1005_b N_A_30_443#_c_178_n 0.0405221f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_66 N_VPB_M1005_b N_A_30_443#_c_179_n 0.0210265f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_67 N_VPB_M1005_b N_A_30_443#_c_170_n 0.0253283f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_68 N_VPB_M1005_b N_A_30_443#_c_181_n 0.0179059f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_69 N_VPB_M1005_b N_A_30_443#_c_182_n 0.00127674f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_70 VPB N_A_30_443#_c_182_n 0.00347996f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_71 N_VPB_c_71_p N_A_30_443#_c_182_n 0.0551782f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_72 VPB N_A_30_443#_c_185_n 8.21022e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_73 N_VPB_c_71_p N_A_30_443#_c_185_n 0.0108189f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_74 N_VPB_M1005_b N_A_30_443#_c_187_n 0.00714214f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_75 N_VPB_M1005_b N_A_30_443#_c_171_n 0.00689372f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_76 N_VPB_M1005_b N_A_30_443#_c_189_n 0.00770964f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_77 N_VPB_M1005_b N_A_30_443#_c_190_n 0.0874174f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_78 VPB N_A_30_443#_c_190_n 0.00282611f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_79 N_VPB_c_71_p N_A_30_443#_c_190_n 0.010545f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_80 N_VPB_M1005_b N_D_c_313_n 0.0519002f $X=-0.33 $Y=1.885 $X2=0.89 $Y2=0.745
cc_81 N_VPB_M1005_b N_D_M1013_g 0.0465925f $X=-0.33 $Y=1.885 $X2=0.635 $Y2=1.21
cc_82 VPB N_D_M1013_g 0.00282611f $X=0 $Y=3.955 $X2=0.635 $Y2=1.21
cc_83 N_VPB_c_71_p N_D_M1013_g 0.0112133f $X=7.92 $Y=4.07 $X2=0.635 $Y2=1.21
cc_84 N_VPB_M1005_b N_D_c_317_n 0.0369051f $X=-0.33 $Y=1.885 $X2=0.777 $Y2=1.28
cc_85 N_VPB_M1005_b N_D_c_311_n 0.0185447f $X=-0.33 $Y=1.885 $X2=0.777 $Y2=1.805
cc_86 N_VPB_M1005_b N_D_c_312_n 0.00792337f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_87 N_VPB_M1005_b N_A_384_107#_c_359_n 0.00962522f $X=-0.33 $Y=1.885 $X2=0.705
+ $Y2=1.28
cc_88 N_VPB_M1005_b N_A_384_107#_c_367_n 0.0344101f $X=-0.33 $Y=1.885 $X2=0.705
+ $Y2=1.28
cc_89 N_VPB_M1005_b N_A_384_107#_c_368_n 0.0245246f $X=-0.33 $Y=1.885 $X2=0.777
+ $Y2=1.085
cc_90 N_VPB_M1005_b N_A_384_107#_c_369_n 0.0808305f $X=-0.33 $Y=1.885 $X2=0.777
+ $Y2=1.805
cc_91 N_VPB_M1005_b N_A_384_107#_M1014_g 0.0395797f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_92 VPB N_A_384_107#_M1014_g 0.00190694f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_93 N_VPB_c_71_p N_A_384_107#_M1014_g 0.00837567f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_94 N_VPB_M1005_b N_A_384_107#_c_373_n 0.00294837f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_95 N_VPB_M1005_b N_A_384_107#_c_363_n 0.00385334f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_96 N_VPB_M1005_b N_A_1004_81#_c_463_n 7.06744e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_97 N_VPB_M1005_b N_A_1004_81#_c_464_n 0.00188754f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_98 N_VPB_M1005_b N_A_1004_81#_c_461_n 0.132553f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_99 N_VPB_c_71_p N_A_1004_81#_c_461_n 0.0017044f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_100 N_VPB_M1005_b N_A_1004_81#_c_467_n 0.0152312f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_101 N_VPB_M1005_b N_A_806_107#_M1008_g 0.0451831f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.21
cc_102 N_VPB_M1005_b N_A_806_107#_M1002_g 0.0425053f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_103 VPB N_A_806_107#_M1002_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_104 N_VPB_c_71_p N_A_806_107#_M1002_g 0.0162989f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_105 N_VPB_M1005_b N_A_806_107#_c_541_n 0.0024757f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_106 N_VPB_M1005_b N_A_806_107#_c_542_n 0.00642854f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_107 VPB N_A_806_107#_c_542_n 7.25672e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_108 N_VPB_c_71_p N_A_806_107#_c_542_n 0.0115764f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_109 N_VPB_M1005_b N_A_806_107#_c_545_n 8.87644e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_110 N_VPB_M1005_b N_A_806_107#_c_546_n 0.00864329f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_111 N_VPB_M1005_b N_A_806_107#_c_534_n 9.57556e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_112 N_VPB_M1005_b N_A_806_107#_c_535_n 0.0186217f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_113 N_VPB_M1005_b N_A_806_107#_c_536_n 0.0475855f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_114 N_VPB_M1005_b N_VPWR_c_633_n 0.047351f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_633_n 0.00252021f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_116 N_VPB_c_71_p N_VPWR_c_633_n 0.0384021f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_117 N_VPB_M1005_b N_VPWR_c_636_n 0.0309249f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_636_n 0.00272896f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_119 N_VPB_c_71_p N_VPWR_c_636_n 0.0408779f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_120 N_VPB_M1005_b N_VPWR_c_639_n 0.0357629f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_639_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_122 N_VPB_c_71_p N_VPWR_c_639_n 0.0409968f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_123 N_VPB_M1005_b N_VPWR_c_642_n 0.0278947f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_642_n 0.00335473f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_125 N_VPB_c_71_p N_VPWR_c_642_n 0.0490696f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_126 N_VPB_M1005_b N_VPWR_c_645_n 0.112253f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_645_n 0.869942f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_128 N_VPB_c_71_p N_VPWR_c_645_n 0.0405284f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_129 N_VPB_M1005_b N_A_650_107#_c_692_n 0.00187603f $X=-0.33 $Y=1.885
+ $X2=0.705 $Y2=1.28
cc_130 N_VPB_M1005_b N_A_650_107#_c_693_n 0.00622092f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_131 N_VPB_M1005_b N_A_650_107#_c_694_n 0.00367553f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_132 N_VPB_M1005_b N_A_650_107#_c_691_n 0.00152241f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_133 N_VPB_M1005_b N_A_650_107#_c_696_n 0.0132212f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_134 N_VPB_M1005_b N_Q_c_751_n 0.0678887f $X=-0.33 $Y=1.885 $X2=0.705 $Y2=1.28
cc_135 VPB N_Q_c_751_n 0.00110823f $X=0 $Y=3.955 $X2=0.705 $Y2=1.28
cc_136 N_VPB_c_71_p N_Q_c_751_n 0.0182942f $X=7.92 $Y=4.07 $X2=0.705 $Y2=1.28
cc_137 N_GATE_M1010_g N_A_30_443#_M1000_g 0.027146f $X=0.89 $Y=0.745 $X2=0 $Y2=0
cc_138 GATE N_A_30_443#_M1000_g 0.00185351f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_139 N_GATE_M1005_g N_A_30_443#_M1011_g 0.0116868f $X=0.665 $Y=2.59 $X2=0
+ $Y2=0
cc_140 N_GATE_M1010_g N_A_30_443#_c_169_n 0.00327546f $X=0.89 $Y=0.745 $X2=7.92
+ $Y2=0
cc_141 GATE N_A_30_443#_c_169_n 0.0407856f $X=0.635 $Y=1.21 $X2=7.92 $Y2=0
cc_142 N_GATE_c_140_n N_A_30_443#_c_169_n 0.0297595f $X=0.705 $Y=1.28 $X2=7.92
+ $Y2=0
cc_143 N_GATE_M1005_g N_A_30_443#_c_178_n 0.0088236f $X=0.665 $Y=2.59 $X2=0
+ $Y2=0
cc_144 N_GATE_M1005_g N_A_30_443#_c_179_n 0.0373789f $X=0.665 $Y=2.59 $X2=4.08
+ $Y2=0
cc_145 GATE N_A_30_443#_c_179_n 0.0234404f $X=0.635 $Y=1.21 $X2=4.08 $Y2=0
cc_146 N_GATE_c_140_n N_A_30_443#_c_179_n 0.010077f $X=0.705 $Y=1.28 $X2=4.08
+ $Y2=0
cc_147 N_GATE_M1005_g N_A_30_443#_c_203_n 5.15034e-19 $X=0.665 $Y=2.59 $X2=4.08
+ $Y2=0.058
cc_148 GATE N_A_30_443#_c_203_n 0.00887751f $X=0.635 $Y=1.21 $X2=4.08 $Y2=0.058
cc_149 N_GATE_c_140_n N_A_30_443#_c_203_n 0.00202248f $X=0.705 $Y=1.28 $X2=4.08
+ $Y2=0.058
cc_150 N_GATE_M1005_g N_A_30_443#_c_170_n 0.00659872f $X=0.665 $Y=2.59 $X2=0
+ $Y2=0
cc_151 N_GATE_c_140_n N_A_30_443#_c_170_n 0.027146f $X=0.705 $Y=1.28 $X2=0 $Y2=0
cc_152 N_GATE_M1005_g N_A_30_443#_c_208_n 8.69114e-19 $X=0.665 $Y=2.59 $X2=0
+ $Y2=0
cc_153 N_GATE_M1010_g N_A_30_443#_c_172_n 0.0106459f $X=0.89 $Y=0.745 $X2=0
+ $Y2=0
cc_154 GATE N_A_30_443#_c_172_n 0.00968915f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_155 N_GATE_c_140_n N_A_30_443#_c_172_n 0.00932901f $X=0.705 $Y=1.28 $X2=0
+ $Y2=0
cc_156 N_GATE_M1005_g N_VPWR_c_633_n 0.0594475f $X=0.665 $Y=2.59 $X2=7.92 $Y2=0
cc_157 N_GATE_M1005_g N_VPWR_c_645_n 0.00357298f $X=0.665 $Y=2.59 $X2=0 $Y2=0
cc_158 N_GATE_M1010_g N_VGND_c_766_n 0.0457062f $X=0.89 $Y=0.745 $X2=7.92 $Y2=0
cc_159 GATE N_VGND_c_766_n 0.00175812f $X=0.635 $Y=1.21 $X2=7.92 $Y2=0
cc_160 N_GATE_M1010_g N_VGND_c_774_n 0.00627686f $X=0.89 $Y=0.745 $X2=0 $Y2=0
cc_161 GATE N_VGND_c_774_n 0.00623385f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_162 N_A_30_443#_c_190_n N_D_c_313_n 0.0385587f $X=3.885 $Y=2.61 $X2=0 $Y2=0
cc_163 N_A_30_443#_c_181_n N_D_M1013_g 0.00876749f $X=3.02 $Y=2.73 $X2=0 $Y2=0
cc_164 N_A_30_443#_c_214_p N_D_M1013_g 0.0365907f $X=3.105 $Y=3.635 $X2=0 $Y2=0
cc_165 N_A_30_443#_c_182_n N_D_M1013_g 0.00767174f $X=3.88 $Y=3.72 $X2=0 $Y2=0
cc_166 N_A_30_443#_c_185_n N_D_M1013_g 0.00547635f $X=3.19 $Y=3.72 $X2=0 $Y2=0
cc_167 N_A_30_443#_c_217_p N_D_M1013_g 0.00124415f $X=3.965 $Y=3.635 $X2=0 $Y2=0
cc_168 N_A_30_443#_c_181_n N_D_c_317_n 0.0225367f $X=3.02 $Y=2.73 $X2=0.24 $Y2=0
cc_169 N_A_30_443#_c_170_n N_D_c_312_n 0.00222299f $X=1.705 $Y=1.51 $X2=7.92
+ $Y2=0
cc_170 N_A_30_443#_c_181_n N_D_c_312_n 0.0440693f $X=3.02 $Y=2.73 $X2=7.92 $Y2=0
cc_171 N_A_30_443#_c_181_n N_A_384_107#_M1011_d 0.00532528f $X=3.02 $Y=2.73
+ $X2=0 $Y2=0
cc_172 N_A_30_443#_M1007_g N_A_384_107#_M1015_g 0.0280825f $X=4.56 $Y=0.745
+ $X2=0 $Y2=0
cc_173 N_A_30_443#_c_187_n N_A_384_107#_c_367_n 0.00601317f $X=4.41 $Y=2.615
+ $X2=0 $Y2=0
cc_174 N_A_30_443#_c_171_n N_A_384_107#_c_367_n 0.0101445f $X=4.575 $Y=1.25
+ $X2=0 $Y2=0
cc_175 N_A_30_443#_M1007_g N_A_384_107#_c_367_n 0.0350844f $X=4.56 $Y=0.745
+ $X2=0 $Y2=0
cc_176 N_A_30_443#_c_226_p N_A_384_107#_c_368_n 2.82903e-19 $X=3.965 $Y=2.715
+ $X2=0 $Y2=0
cc_177 N_A_30_443#_c_190_n N_A_384_107#_c_368_n 0.0328499f $X=3.885 $Y=2.61
+ $X2=0 $Y2=0
cc_178 N_A_30_443#_c_217_p N_A_384_107#_c_369_n 4.94666e-19 $X=3.965 $Y=3.635
+ $X2=0 $Y2=0
cc_179 N_A_30_443#_c_187_n N_A_384_107#_c_369_n 0.0123142f $X=4.41 $Y=2.615
+ $X2=0 $Y2=0
cc_180 N_A_30_443#_c_171_n N_A_384_107#_c_369_n 0.0234062f $X=4.575 $Y=1.25
+ $X2=0 $Y2=0
cc_181 N_A_30_443#_c_190_n N_A_384_107#_c_369_n 0.0130105f $X=3.885 $Y=2.61
+ $X2=0 $Y2=0
cc_182 N_A_30_443#_c_217_p N_A_384_107#_M1014_g 7.10852e-19 $X=3.965 $Y=3.635
+ $X2=7.92 $Y2=0
cc_183 N_A_30_443#_c_190_n N_A_384_107#_M1014_g 0.0132701f $X=3.885 $Y=2.61
+ $X2=7.92 $Y2=0
cc_184 N_A_30_443#_M1000_g N_A_384_107#_c_360_n 0.0177317f $X=1.67 $Y=0.745
+ $X2=0 $Y2=0
cc_185 N_A_30_443#_c_203_n N_A_384_107#_c_360_n 0.00684578f $X=1.705 $Y=1.51
+ $X2=0 $Y2=0
cc_186 N_A_30_443#_c_170_n N_A_384_107#_c_360_n 0.00490064f $X=1.705 $Y=1.51
+ $X2=0 $Y2=0
cc_187 N_A_30_443#_M1011_g N_A_384_107#_c_373_n 0.00586228f $X=1.735 $Y=2.59
+ $X2=0 $Y2=0
cc_188 N_A_30_443#_c_208_n N_A_384_107#_c_373_n 0.0184176f $X=1.695 $Y=2.645
+ $X2=0 $Y2=0
cc_189 N_A_30_443#_c_181_n N_A_384_107#_c_373_n 0.0210092f $X=3.02 $Y=2.73 $X2=0
+ $Y2=0
cc_190 N_A_30_443#_M1011_g N_A_384_107#_c_363_n 0.00390292f $X=1.735 $Y=2.59
+ $X2=0 $Y2=0
cc_191 N_A_30_443#_c_203_n N_A_384_107#_c_363_n 0.0202415f $X=1.705 $Y=1.51
+ $X2=0 $Y2=0
cc_192 N_A_30_443#_c_170_n N_A_384_107#_c_363_n 0.0166644f $X=1.705 $Y=1.51
+ $X2=0 $Y2=0
cc_193 N_A_30_443#_c_208_n N_A_384_107#_c_363_n 0.00752177f $X=1.695 $Y=2.645
+ $X2=0 $Y2=0
cc_194 N_A_30_443#_c_244_p N_A_384_107#_c_363_n 0.012631f $X=1.54 $Y=1.905 $X2=0
+ $Y2=0
cc_195 N_A_30_443#_c_203_n N_A_384_107#_c_364_n 0.0127216f $X=1.705 $Y=1.51
+ $X2=0 $Y2=0
cc_196 N_A_30_443#_c_170_n N_A_384_107#_c_364_n 0.00694394f $X=1.705 $Y=1.51
+ $X2=0 $Y2=0
cc_197 N_A_30_443#_M1007_g N_A_384_107#_c_365_n 0.0204894f $X=4.56 $Y=0.745
+ $X2=0 $Y2=0
cc_198 N_A_30_443#_M1007_g N_A_1004_81#_c_455_n 0.0773152f $X=4.56 $Y=0.745
+ $X2=0 $Y2=0
cc_199 N_A_30_443#_c_171_n N_A_1004_81#_c_457_n 4.30005e-19 $X=4.575 $Y=1.25
+ $X2=0 $Y2=0
cc_200 N_A_30_443#_c_171_n N_A_1004_81#_c_461_n 7.34845e-19 $X=4.575 $Y=1.25
+ $X2=0 $Y2=0
cc_201 N_A_30_443#_M1007_g N_A_1004_81#_c_461_n 0.00413645f $X=4.56 $Y=0.745
+ $X2=0 $Y2=0
cc_202 N_A_30_443#_c_217_p N_A_806_107#_c_541_n 0.00727363f $X=3.965 $Y=3.635
+ $X2=4.08 $Y2=0.057
cc_203 N_A_30_443#_c_187_n N_A_806_107#_c_541_n 0.0209769f $X=4.41 $Y=2.615
+ $X2=4.08 $Y2=0.057
cc_204 N_A_30_443#_c_190_n N_A_806_107#_c_541_n 4.57034e-19 $X=3.885 $Y=2.61
+ $X2=4.08 $Y2=0.057
cc_205 N_A_30_443#_c_182_n N_A_806_107#_c_542_n 0.00497652f $X=3.88 $Y=3.72
+ $X2=4.08 $Y2=0.058
cc_206 N_A_30_443#_c_217_p N_A_806_107#_c_542_n 0.0212598f $X=3.965 $Y=3.635
+ $X2=4.08 $Y2=0.058
cc_207 N_A_30_443#_c_190_n N_A_806_107#_c_542_n 0.00199868f $X=3.885 $Y=2.61
+ $X2=4.08 $Y2=0.058
cc_208 N_A_30_443#_c_171_n N_A_806_107#_c_530_n 0.0226757f $X=4.575 $Y=1.25
+ $X2=0 $Y2=0
cc_209 N_A_30_443#_M1007_g N_A_806_107#_c_530_n 0.0304819f $X=4.56 $Y=0.745
+ $X2=0 $Y2=0
cc_210 N_A_30_443#_c_187_n N_A_806_107#_c_545_n 0.0194512f $X=4.41 $Y=2.615
+ $X2=0 $Y2=0
cc_211 N_A_30_443#_c_171_n N_A_806_107#_c_531_n 0.0534801f $X=4.575 $Y=1.25
+ $X2=0 $Y2=0
cc_212 N_A_30_443#_M1007_g N_A_806_107#_c_531_n 0.00918915f $X=4.56 $Y=0.745
+ $X2=0 $Y2=0
cc_213 N_A_30_443#_c_187_n N_A_806_107#_c_546_n 0.0145485f $X=4.41 $Y=2.615
+ $X2=0 $Y2=0
cc_214 N_A_30_443#_c_171_n N_A_806_107#_c_546_n 0.0347205f $X=4.575 $Y=1.25
+ $X2=0 $Y2=0
cc_215 N_A_30_443#_M1007_g N_A_806_107#_c_532_n 0.0090244f $X=4.56 $Y=0.745
+ $X2=0 $Y2=0
cc_216 N_A_30_443#_c_171_n N_A_806_107#_c_534_n 0.0142666f $X=4.575 $Y=1.25
+ $X2=0 $Y2=0
cc_217 N_A_30_443#_M1011_g N_VPWR_c_633_n 0.0101281f $X=1.735 $Y=2.59 $X2=7.92
+ $Y2=0
cc_218 N_A_30_443#_c_178_n N_VPWR_c_633_n 0.0299621f $X=0.275 $Y=2.36 $X2=7.92
+ $Y2=0
cc_219 N_A_30_443#_c_179_n N_VPWR_c_633_n 0.0654022f $X=1.54 $Y=1.99 $X2=7.92
+ $Y2=0
cc_220 N_A_30_443#_c_170_n N_VPWR_c_633_n 2.43438e-19 $X=1.705 $Y=1.51 $X2=7.92
+ $Y2=0
cc_221 N_A_30_443#_M1011_g N_VPWR_c_636_n 0.00904199f $X=1.735 $Y=2.59 $X2=0
+ $Y2=0
cc_222 N_A_30_443#_c_181_n N_VPWR_c_636_n 0.070712f $X=3.02 $Y=2.73 $X2=0 $Y2=0
cc_223 N_A_30_443#_c_214_p N_VPWR_c_636_n 0.0443401f $X=3.105 $Y=3.635 $X2=0
+ $Y2=0
cc_224 N_A_30_443#_c_185_n N_VPWR_c_636_n 0.00430349f $X=3.19 $Y=3.72 $X2=0
+ $Y2=0
cc_225 N_A_30_443#_M1011_g N_VPWR_c_645_n 0.0114846f $X=1.735 $Y=2.59 $X2=0
+ $Y2=0
cc_226 N_A_30_443#_c_178_n N_VPWR_c_645_n 0.0107528f $X=0.275 $Y=2.36 $X2=0
+ $Y2=0
cc_227 N_A_30_443#_c_214_p N_VPWR_c_645_n 0.0199533f $X=3.105 $Y=3.635 $X2=0
+ $Y2=0
cc_228 N_A_30_443#_c_182_n N_VPWR_c_645_n 0.0308119f $X=3.88 $Y=3.72 $X2=0 $Y2=0
cc_229 N_A_30_443#_c_185_n N_VPWR_c_645_n 0.0069161f $X=3.19 $Y=3.72 $X2=0 $Y2=0
cc_230 N_A_30_443#_c_217_p N_VPWR_c_645_n 0.0199629f $X=3.965 $Y=3.635 $X2=0
+ $Y2=0
cc_231 N_A_30_443#_c_190_n N_VPWR_c_645_n 0.0174165f $X=3.885 $Y=2.61 $X2=0
+ $Y2=0
cc_232 N_A_30_443#_c_182_n N_A_650_107#_M1013_d 0.0012031f $X=3.88 $Y=3.72 $X2=0
+ $Y2=0
cc_233 N_A_30_443#_c_217_p N_A_650_107#_c_692_n 0.038092f $X=3.965 $Y=3.635
+ $X2=0 $Y2=0
cc_234 N_A_30_443#_c_190_n N_A_650_107#_c_692_n 0.00480908f $X=3.885 $Y=2.61
+ $X2=0 $Y2=0
cc_235 N_A_30_443#_c_182_n N_A_650_107#_c_700_n 0.0195527f $X=3.88 $Y=3.72 $X2=0
+ $Y2=0
cc_236 N_A_30_443#_c_190_n N_A_650_107#_c_700_n 0.00718685f $X=3.885 $Y=2.61
+ $X2=0 $Y2=0
cc_237 N_A_30_443#_c_226_p N_A_650_107#_c_693_n 0.0241533f $X=3.965 $Y=2.715
+ $X2=7.92 $Y2=0
cc_238 N_A_30_443#_c_187_n N_A_650_107#_c_693_n 0.0140271f $X=4.41 $Y=2.615
+ $X2=7.92 $Y2=0
cc_239 N_A_30_443#_c_171_n N_A_650_107#_c_693_n 0.0140042f $X=4.575 $Y=1.25
+ $X2=7.92 $Y2=0
cc_240 N_A_30_443#_c_190_n N_A_650_107#_c_693_n 0.00408185f $X=3.885 $Y=2.61
+ $X2=7.92 $Y2=0
cc_241 N_A_30_443#_c_171_n N_A_650_107#_c_690_n 0.0137305f $X=4.575 $Y=1.25
+ $X2=0 $Y2=0
cc_242 N_A_30_443#_M1007_g N_A_650_107#_c_690_n 0.0015524f $X=4.56 $Y=0.745
+ $X2=0 $Y2=0
cc_243 N_A_30_443#_c_171_n N_A_650_107#_c_691_n 0.0649104f $X=4.575 $Y=1.25
+ $X2=0 $Y2=0
cc_244 N_A_30_443#_M1007_g N_A_650_107#_c_691_n 0.00388756f $X=4.56 $Y=0.745
+ $X2=0 $Y2=0
cc_245 N_A_30_443#_c_181_n N_A_650_107#_c_696_n 0.0129653f $X=3.02 $Y=2.73
+ $X2=4.08 $Y2=0.058
cc_246 N_A_30_443#_c_214_p N_A_650_107#_c_696_n 0.0252495f $X=3.105 $Y=3.635
+ $X2=4.08 $Y2=0.058
cc_247 N_A_30_443#_c_226_p N_A_650_107#_c_696_n 0.0153021f $X=3.965 $Y=2.715
+ $X2=4.08 $Y2=0.058
cc_248 N_A_30_443#_c_217_p N_A_650_107#_c_696_n 0.00764029f $X=3.965 $Y=3.635
+ $X2=4.08 $Y2=0.058
cc_249 N_A_30_443#_c_190_n N_A_650_107#_c_696_n 0.00562354f $X=3.885 $Y=2.61
+ $X2=4.08 $Y2=0.058
cc_250 N_A_30_443#_M1000_g N_VGND_c_766_n 0.0453952f $X=1.67 $Y=0.745 $X2=7.92
+ $Y2=0
cc_251 N_A_30_443#_c_203_n N_VGND_c_766_n 0.0118731f $X=1.705 $Y=1.51 $X2=7.92
+ $Y2=0
cc_252 N_A_30_443#_c_172_n N_VGND_c_766_n 0.037224f $X=0.5 $Y=0.745 $X2=7.92
+ $Y2=0
cc_253 N_A_30_443#_M1000_g N_VGND_c_768_n 0.00200035f $X=1.67 $Y=0.745 $X2=4.08
+ $Y2=0.058
cc_254 N_A_30_443#_M1007_g N_VGND_c_770_n 0.00217486f $X=4.56 $Y=0.745 $X2=0
+ $Y2=0
cc_255 N_A_30_443#_M1000_g N_VGND_c_774_n 0.00936553f $X=1.67 $Y=0.745 $X2=0
+ $Y2=0
cc_256 N_A_30_443#_c_169_n N_VGND_c_774_n 6.69455e-19 $X=0.235 $Y=1.905 $X2=0
+ $Y2=0
cc_257 N_A_30_443#_c_172_n N_VGND_c_774_n 0.0337119f $X=0.5 $Y=0.745 $X2=0 $Y2=0
cc_258 N_A_30_443#_M1007_g N_VGND_c_774_n 0.0151022f $X=4.56 $Y=0.745 $X2=0
+ $Y2=0
cc_259 N_D_M1004_g N_A_384_107#_M1015_g 0.0489374f $X=3 $Y=0.745 $X2=0 $Y2=0
cc_260 N_D_c_311_n N_A_384_107#_c_359_n 0.015806f $X=2.935 $Y=1.96 $X2=0 $Y2=0
cc_261 N_D_c_312_n N_A_384_107#_c_359_n 0.00138349f $X=2.935 $Y=1.96 $X2=0 $Y2=0
cc_262 N_D_c_313_n N_A_384_107#_c_368_n 0.015806f $X=3.035 $Y=2.52 $X2=0 $Y2=0
cc_263 N_D_M1004_g N_A_384_107#_c_360_n 0.0140384f $X=3 $Y=0.745 $X2=0 $Y2=0
cc_264 N_D_M1004_g N_A_384_107#_c_362_n 0.0422921f $X=3 $Y=0.745 $X2=0 $Y2=0
cc_265 N_D_c_311_n N_A_384_107#_c_362_n 0.00293702f $X=2.935 $Y=1.96 $X2=0 $Y2=0
cc_266 N_D_c_312_n N_A_384_107#_c_362_n 0.0434591f $X=2.935 $Y=1.96 $X2=0 $Y2=0
cc_267 N_D_c_313_n N_A_384_107#_c_373_n 0.0014694f $X=3.035 $Y=2.52 $X2=0 $Y2=0
cc_268 N_D_M1004_g N_A_384_107#_c_363_n 0.00561103f $X=3 $Y=0.745 $X2=0 $Y2=0
cc_269 N_D_c_311_n N_A_384_107#_c_363_n 0.0014694f $X=2.935 $Y=1.96 $X2=0 $Y2=0
cc_270 N_D_c_312_n N_A_384_107#_c_363_n 0.0463343f $X=2.935 $Y=1.96 $X2=0 $Y2=0
cc_271 N_D_M1004_g N_A_384_107#_c_414_n 0.00108234f $X=3 $Y=0.745 $X2=0 $Y2=0
cc_272 N_D_c_311_n N_A_384_107#_c_414_n 9.53483e-19 $X=2.935 $Y=1.96 $X2=0 $Y2=0
cc_273 N_D_c_312_n N_A_384_107#_c_414_n 0.00672602f $X=2.935 $Y=1.96 $X2=0 $Y2=0
cc_274 N_D_M1013_g N_VPWR_c_636_n 0.0126198f $X=3.07 $Y=3.31 $X2=0 $Y2=0
cc_275 N_D_c_317_n N_VPWR_c_636_n 3.52969e-19 $X=3.035 $Y=2.805 $X2=0 $Y2=0
cc_276 N_D_M1013_g N_VPWR_c_645_n 0.017461f $X=3.07 $Y=3.31 $X2=0 $Y2=0
cc_277 N_D_M1004_g N_A_650_107#_c_687_n 0.0122636f $X=3 $Y=0.745 $X2=0 $Y2=0
cc_278 N_D_M1004_g N_A_650_107#_c_688_n 0.00626181f $X=3 $Y=0.745 $X2=0 $Y2=0
cc_279 N_D_c_317_n N_A_650_107#_c_692_n 0.00482713f $X=3.035 $Y=2.805 $X2=0
+ $Y2=0
cc_280 N_D_M1013_g N_A_650_107#_c_700_n 0.00482713f $X=3.07 $Y=3.31 $X2=0 $Y2=0
cc_281 N_D_c_313_n N_A_650_107#_c_694_n 0.00436425f $X=3.035 $Y=2.52 $X2=0 $Y2=0
cc_282 N_D_c_312_n N_A_650_107#_c_694_n 0.0105728f $X=2.935 $Y=1.96 $X2=0 $Y2=0
cc_283 N_D_c_313_n N_A_650_107#_c_696_n 0.00482713f $X=3.035 $Y=2.52 $X2=4.08
+ $Y2=0.058
cc_284 N_D_c_312_n N_A_650_107#_c_696_n 0.00714931f $X=2.935 $Y=1.96 $X2=4.08
+ $Y2=0.058
cc_285 N_D_M1004_g N_VGND_c_768_n 0.0354518f $X=3 $Y=0.745 $X2=4.08 $Y2=0.058
cc_286 N_D_M1004_g N_VGND_c_774_n 0.0140308f $X=3 $Y=0.745 $X2=0 $Y2=0
cc_287 N_A_384_107#_c_369_n N_A_1004_81#_c_457_n 8.69855e-19 $X=4.82 $Y=2.805
+ $X2=0 $Y2=0
cc_288 N_A_384_107#_c_369_n N_A_1004_81#_c_461_n 0.0951576f $X=4.82 $Y=2.805
+ $X2=0 $Y2=0
cc_289 N_A_384_107#_c_367_n N_A_806_107#_c_541_n 4.53651e-19 $X=4.54 $Y=2.1
+ $X2=4.08 $Y2=0.057
cc_290 N_A_384_107#_M1014_g N_A_806_107#_c_542_n 0.0113374f $X=4.82 $Y=3.145
+ $X2=4.08 $Y2=0.058
cc_291 N_A_384_107#_c_369_n N_A_806_107#_c_545_n 8.72107e-19 $X=4.82 $Y=2.805
+ $X2=0 $Y2=0
cc_292 N_A_384_107#_M1014_g N_A_806_107#_c_545_n 0.0303122f $X=4.82 $Y=3.145
+ $X2=0 $Y2=0
cc_293 N_A_384_107#_c_369_n N_A_806_107#_c_546_n 0.0266789f $X=4.82 $Y=2.805
+ $X2=0 $Y2=0
cc_294 N_A_384_107#_M1014_g N_A_806_107#_c_546_n 0.00495557f $X=4.82 $Y=3.145
+ $X2=0 $Y2=0
cc_295 N_A_384_107#_M1015_g N_A_806_107#_c_532_n 0.0112382f $X=3.78 $Y=0.745
+ $X2=0 $Y2=0
cc_296 N_A_384_107#_c_369_n N_A_806_107#_c_534_n 0.00357117f $X=4.82 $Y=2.805
+ $X2=0 $Y2=0
cc_297 N_A_384_107#_M1014_g N_VPWR_c_639_n 0.00423015f $X=4.82 $Y=3.145 $X2=0
+ $Y2=0
cc_298 N_A_384_107#_M1014_g N_VPWR_c_645_n 0.0140817f $X=4.82 $Y=3.145 $X2=0
+ $Y2=0
cc_299 N_A_384_107#_M1015_g N_A_650_107#_c_687_n 0.0138045f $X=3.78 $Y=0.745
+ $X2=0 $Y2=0
cc_300 N_A_384_107#_c_362_n N_A_650_107#_c_687_n 0.0196839f $X=3.55 $Y=1.53
+ $X2=0 $Y2=0
cc_301 N_A_384_107#_c_414_n N_A_650_107#_c_687_n 3.98497e-19 $X=3.715 $Y=1.545
+ $X2=0 $Y2=0
cc_302 N_A_384_107#_M1015_g N_A_650_107#_c_688_n 0.00864664f $X=3.78 $Y=0.745
+ $X2=0 $Y2=0
cc_303 N_A_384_107#_c_368_n N_A_650_107#_c_692_n 7.18317e-19 $X=4.06 $Y=2.1
+ $X2=0 $Y2=0
cc_304 N_A_384_107#_c_367_n N_A_650_107#_c_693_n 0.00301882f $X=4.54 $Y=2.1
+ $X2=7.92 $Y2=0
cc_305 N_A_384_107#_c_368_n N_A_650_107#_c_693_n 0.0193005f $X=4.06 $Y=2.1
+ $X2=7.92 $Y2=0
cc_306 N_A_384_107#_c_369_n N_A_650_107#_c_693_n 6.88575e-19 $X=4.82 $Y=2.805
+ $X2=7.92 $Y2=0
cc_307 N_A_384_107#_c_362_n N_A_650_107#_c_693_n 2.32646e-19 $X=3.55 $Y=1.53
+ $X2=7.92 $Y2=0
cc_308 N_A_384_107#_c_414_n N_A_650_107#_c_693_n 0.0234047f $X=3.715 $Y=1.545
+ $X2=7.92 $Y2=0
cc_309 N_A_384_107#_c_368_n N_A_650_107#_c_694_n 8.70892e-19 $X=4.06 $Y=2.1
+ $X2=0 $Y2=0
cc_310 N_A_384_107#_c_362_n N_A_650_107#_c_694_n 0.00626001f $X=3.55 $Y=1.53
+ $X2=0 $Y2=0
cc_311 N_A_384_107#_M1015_g N_A_650_107#_c_690_n 0.0301256f $X=3.78 $Y=0.745
+ $X2=0 $Y2=0
cc_312 N_A_384_107#_c_414_n N_A_650_107#_c_690_n 0.0231595f $X=3.715 $Y=1.545
+ $X2=0 $Y2=0
cc_313 N_A_384_107#_c_365_n N_A_650_107#_c_690_n 0.00133216f $X=3.715 $Y=1.545
+ $X2=0 $Y2=0
cc_314 N_A_384_107#_M1015_g N_A_650_107#_c_691_n 0.00244788f $X=3.78 $Y=0.745
+ $X2=0 $Y2=0
cc_315 N_A_384_107#_c_367_n N_A_650_107#_c_691_n 0.0169658f $X=4.54 $Y=2.1 $X2=0
+ $Y2=0
cc_316 N_A_384_107#_c_414_n N_A_650_107#_c_691_n 0.0395283f $X=3.715 $Y=1.545
+ $X2=0 $Y2=0
cc_317 N_A_384_107#_c_365_n N_A_650_107#_c_691_n 0.0115865f $X=3.715 $Y=1.545
+ $X2=0 $Y2=0
cc_318 N_A_384_107#_c_360_n N_VGND_c_766_n 0.0218749f $X=2.06 $Y=0.745 $X2=7.92
+ $Y2=0
cc_319 N_A_384_107#_M1015_g N_VGND_c_768_n 7.89605e-19 $X=3.78 $Y=0.745 $X2=4.08
+ $Y2=0.058
cc_320 N_A_384_107#_c_360_n N_VGND_c_768_n 0.0362217f $X=2.06 $Y=0.745 $X2=4.08
+ $Y2=0.058
cc_321 N_A_384_107#_c_362_n N_VGND_c_768_n 0.0222591f $X=3.55 $Y=1.53 $X2=4.08
+ $Y2=0.058
cc_322 N_A_384_107#_M1000_d N_VGND_c_774_n 0.00221032f $X=1.92 $Y=0.535 $X2=0
+ $Y2=0
cc_323 N_A_384_107#_M1015_g N_VGND_c_774_n 0.0152606f $X=3.78 $Y=0.745 $X2=0
+ $Y2=0
cc_324 N_A_384_107#_c_360_n N_VGND_c_774_n 0.0236764f $X=2.06 $Y=0.745 $X2=0
+ $Y2=0
cc_325 N_A_1004_81#_c_463_n N_A_806_107#_M1008_g 0.0299853f $X=6.86 $Y=2.27
+ $X2=0 $Y2=0
cc_326 N_A_1004_81#_c_464_n N_A_806_107#_M1008_g 0.00277582f $X=6.945 $Y=2.185
+ $X2=0 $Y2=0
cc_327 N_A_1004_81#_c_461_n N_A_806_107#_M1008_g 0.0134164f $X=5.595 $Y=1.57
+ $X2=0 $Y2=0
cc_328 N_A_1004_81#_c_467_n N_A_806_107#_M1008_g 0.014644f $X=6.19 $Y=2.27 $X2=0
+ $Y2=0
cc_329 N_A_1004_81#_c_457_n N_A_806_107#_M1003_g 0.00395573f $X=5.595 $Y=1.23
+ $X2=0 $Y2=0
cc_330 N_A_1004_81#_c_459_n N_A_806_107#_M1003_g 0.0179641f $X=6.21 $Y=1.075
+ $X2=0 $Y2=0
cc_331 N_A_1004_81#_c_463_n N_A_806_107#_M1002_g 0.002554f $X=6.86 $Y=2.27
+ $X2=7.92 $Y2=0
cc_332 N_A_1004_81#_c_464_n N_A_806_107#_M1002_g 0.00123404f $X=6.945 $Y=2.185
+ $X2=7.92 $Y2=0
cc_333 N_A_1004_81#_c_460_n N_A_806_107#_M1009_g 0.00233299f $X=6.86 $Y=1.51
+ $X2=4.08 $Y2=0
cc_334 N_A_1004_81#_c_455_n N_A_806_107#_c_530_n 0.00732214f $X=5.27 $Y=1.065
+ $X2=0 $Y2=0
cc_335 N_A_1004_81#_c_461_n N_A_806_107#_c_545_n 2.35572e-19 $X=5.595 $Y=1.57
+ $X2=0 $Y2=0
cc_336 N_A_1004_81#_c_455_n N_A_806_107#_c_531_n 0.00770148f $X=5.27 $Y=1.065
+ $X2=0 $Y2=0
cc_337 N_A_1004_81#_c_486_p N_A_806_107#_c_531_n 0.0101969f $X=5.595 $Y=1.425
+ $X2=0 $Y2=0
cc_338 N_A_1004_81#_c_487_p N_A_806_107#_c_531_n 0.014319f $X=5.595 $Y=1.23
+ $X2=0 $Y2=0
cc_339 N_A_1004_81#_c_457_n N_A_806_107#_c_531_n 0.0170514f $X=5.595 $Y=1.23
+ $X2=0 $Y2=0
cc_340 N_A_1004_81#_c_461_n N_A_806_107#_c_531_n 0.0060798f $X=5.595 $Y=1.57
+ $X2=0 $Y2=0
cc_341 N_A_1004_81#_c_461_n N_A_806_107#_c_546_n 0.0180546f $X=5.595 $Y=1.57
+ $X2=0 $Y2=0
cc_342 N_A_1004_81#_c_455_n N_A_806_107#_c_532_n 9.82792e-19 $X=5.27 $Y=1.065
+ $X2=0 $Y2=0
cc_343 N_A_1004_81#_c_463_n N_A_806_107#_c_591_n 0.0215422f $X=6.86 $Y=2.27
+ $X2=0 $Y2=0
cc_344 N_A_1004_81#_c_460_n N_A_806_107#_c_591_n 0.0201841f $X=6.86 $Y=1.51
+ $X2=0 $Y2=0
cc_345 N_A_1004_81#_c_464_n N_A_806_107#_c_591_n 0.016338f $X=6.945 $Y=2.185
+ $X2=0 $Y2=0
cc_346 N_A_1004_81#_c_461_n N_A_806_107#_c_591_n 3.51214e-19 $X=5.595 $Y=1.57
+ $X2=0 $Y2=0
cc_347 N_A_1004_81#_c_462_n N_A_806_107#_c_591_n 0.00181701f $X=6.21 $Y=1.51
+ $X2=0 $Y2=0
cc_348 N_A_1004_81#_c_486_p N_A_806_107#_c_535_n 0.0236895f $X=5.595 $Y=1.425
+ $X2=0 $Y2=0
cc_349 N_A_1004_81#_c_457_n N_A_806_107#_c_535_n 0.00706945f $X=5.595 $Y=1.23
+ $X2=0 $Y2=0
cc_350 N_A_1004_81#_c_458_n N_A_806_107#_c_535_n 0.0166624f $X=6.045 $Y=1.51
+ $X2=0 $Y2=0
cc_351 N_A_1004_81#_c_461_n N_A_806_107#_c_535_n 0.0481206f $X=5.595 $Y=1.57
+ $X2=0 $Y2=0
cc_352 N_A_1004_81#_c_467_n N_A_806_107#_c_535_n 0.0256738f $X=6.19 $Y=2.27
+ $X2=0 $Y2=0
cc_353 N_A_1004_81#_c_462_n N_A_806_107#_c_535_n 0.0200298f $X=6.21 $Y=1.51
+ $X2=0 $Y2=0
cc_354 N_A_1004_81#_c_486_p N_A_806_107#_c_536_n 3.77595e-19 $X=5.595 $Y=1.425
+ $X2=0 $Y2=0
cc_355 N_A_1004_81#_c_457_n N_A_806_107#_c_536_n 0.0134164f $X=5.595 $Y=1.23
+ $X2=0 $Y2=0
cc_356 N_A_1004_81#_c_459_n N_A_806_107#_c_536_n 0.00103646f $X=6.21 $Y=1.075
+ $X2=0 $Y2=0
cc_357 N_A_1004_81#_c_460_n N_A_806_107#_c_536_n 0.0323416f $X=6.86 $Y=1.51
+ $X2=0 $Y2=0
cc_358 N_A_1004_81#_c_464_n N_A_806_107#_c_536_n 0.0381632f $X=6.945 $Y=2.185
+ $X2=0 $Y2=0
cc_359 N_A_1004_81#_c_462_n N_A_806_107#_c_536_n 0.00456343f $X=6.21 $Y=1.51
+ $X2=0 $Y2=0
cc_360 N_A_1004_81#_c_463_n N_VPWR_M1008_d 0.00389977f $X=6.86 $Y=2.27 $X2=0
+ $Y2=0
cc_361 N_A_1004_81#_c_461_n N_VPWR_c_639_n 0.0682898f $X=5.595 $Y=1.57 $X2=0
+ $Y2=0
cc_362 N_A_1004_81#_c_467_n N_VPWR_c_639_n 0.0147064f $X=6.19 $Y=2.27 $X2=0
+ $Y2=0
cc_363 N_A_1004_81#_c_463_n N_VPWR_c_642_n 0.0337366f $X=6.86 $Y=2.27 $X2=0
+ $Y2=0
cc_364 N_A_1004_81#_c_467_n N_VPWR_c_642_n 0.0106243f $X=6.19 $Y=2.27 $X2=0
+ $Y2=0
cc_365 N_A_1004_81#_c_463_n N_Q_c_751_n 0.00478277f $X=6.86 $Y=2.27 $X2=0 $Y2=0
cc_366 N_A_1004_81#_c_460_n N_Q_c_751_n 0.00498425f $X=6.86 $Y=1.51 $X2=0 $Y2=0
cc_367 N_A_1004_81#_c_464_n N_Q_c_751_n 0.0137606f $X=6.945 $Y=2.185 $X2=0 $Y2=0
cc_368 N_A_1004_81#_c_455_n N_VGND_c_770_n 0.0364619f $X=5.27 $Y=1.065 $X2=0
+ $Y2=0
cc_369 N_A_1004_81#_c_487_p N_VGND_c_770_n 0.0227087f $X=5.595 $Y=1.23 $X2=0
+ $Y2=0
cc_370 N_A_1004_81#_c_457_n N_VGND_c_770_n 0.0070093f $X=5.595 $Y=1.23 $X2=0
+ $Y2=0
cc_371 N_A_1004_81#_c_458_n N_VGND_c_770_n 0.00357969f $X=6.045 $Y=1.51 $X2=0
+ $Y2=0
cc_372 N_A_1004_81#_c_459_n N_VGND_c_770_n 0.00410271f $X=6.21 $Y=1.075 $X2=0
+ $Y2=0
cc_373 N_A_1004_81#_c_459_n N_VGND_c_772_n 0.0303552f $X=6.21 $Y=1.075 $X2=0
+ $Y2=0
cc_374 N_A_1004_81#_c_460_n N_VGND_c_772_n 0.0346705f $X=6.86 $Y=1.51 $X2=0
+ $Y2=0
cc_375 N_A_1004_81#_c_455_n N_VGND_c_774_n 0.0140312f $X=5.27 $Y=1.065 $X2=0
+ $Y2=0
cc_376 N_A_1004_81#_c_487_p N_VGND_c_774_n 0.00139698f $X=5.595 $Y=1.23 $X2=0
+ $Y2=0
cc_377 N_A_1004_81#_c_459_n N_VGND_c_774_n 0.0177898f $X=6.21 $Y=1.075 $X2=0
+ $Y2=0
cc_378 N_A_806_107#_c_545_n N_VPWR_c_639_n 0.0034929f $X=4.92 $Y=2.98 $X2=0
+ $Y2=0
cc_379 N_A_806_107#_M1008_g N_VPWR_c_642_n 0.0279548f $X=6.58 $Y=2.425 $X2=0
+ $Y2=0
cc_380 N_A_806_107#_M1002_g N_VPWR_c_642_n 0.0675823f $X=7.475 $Y=2.965 $X2=0
+ $Y2=0
cc_381 N_A_806_107#_c_536_n N_VPWR_c_642_n 0.00412544f $X=7.475 $Y=1.75 $X2=0
+ $Y2=0
cc_382 N_A_806_107#_M1006_d N_VPWR_c_645_n 0.00221032f $X=4.175 $Y=2.935 $X2=0
+ $Y2=0
cc_383 N_A_806_107#_M1002_g N_VPWR_c_645_n 0.0130327f $X=7.475 $Y=2.965 $X2=0
+ $Y2=0
cc_384 N_A_806_107#_c_542_n N_VPWR_c_645_n 0.0353966f $X=4.315 $Y=3.56 $X2=0
+ $Y2=0
cc_385 N_A_806_107#_c_545_n N_VPWR_c_645_n 0.0220484f $X=4.92 $Y=2.98 $X2=0
+ $Y2=0
cc_386 N_A_806_107#_c_532_n N_A_650_107#_c_687_n 0.00290563f $X=4.17 $Y=0.745
+ $X2=0 $Y2=0
cc_387 N_A_806_107#_c_532_n N_A_650_107#_c_688_n 0.00941113f $X=4.17 $Y=0.745
+ $X2=0 $Y2=0
cc_388 N_A_806_107#_c_532_n N_A_650_107#_c_690_n 0.0152474f $X=4.17 $Y=0.745
+ $X2=0 $Y2=0
cc_389 N_A_806_107#_M1002_g N_Q_c_751_n 0.0413252f $X=7.475 $Y=2.965 $X2=0 $Y2=0
cc_390 N_A_806_107#_M1009_g N_Q_c_751_n 0.0350576f $X=7.495 $Y=0.91 $X2=0 $Y2=0
cc_391 N_A_806_107#_c_536_n N_Q_c_751_n 0.0276045f $X=7.475 $Y=1.75 $X2=0 $Y2=0
cc_392 N_A_806_107#_M1003_g N_VGND_c_770_n 0.00373023f $X=6.6 $Y=1.075 $X2=0
+ $Y2=0
cc_393 N_A_806_107#_c_530_n N_VGND_c_770_n 0.0119358f $X=4.92 $Y=0.83 $X2=0
+ $Y2=0
cc_394 N_A_806_107#_M1003_g N_VGND_c_772_n 0.0436966f $X=6.6 $Y=1.075 $X2=0
+ $Y2=0
cc_395 N_A_806_107#_M1009_g N_VGND_c_772_n 0.0553663f $X=7.495 $Y=0.91 $X2=0
+ $Y2=0
cc_396 N_A_806_107#_c_536_n N_VGND_c_772_n 0.00536236f $X=7.475 $Y=1.75 $X2=0
+ $Y2=0
cc_397 N_A_806_107#_M1003_g N_VGND_c_774_n 0.00672879f $X=6.6 $Y=1.075 $X2=0
+ $Y2=0
cc_398 N_A_806_107#_M1009_g N_VGND_c_774_n 0.0129444f $X=7.495 $Y=0.91 $X2=0
+ $Y2=0
cc_399 N_A_806_107#_c_530_n N_VGND_c_774_n 0.02665f $X=4.92 $Y=0.83 $X2=0 $Y2=0
cc_400 N_A_806_107#_c_532_n N_VGND_c_774_n 0.0250024f $X=4.17 $Y=0.745 $X2=0
+ $Y2=0
cc_401 N_A_806_107#_c_530_n A_962_107# 0.00361414f $X=4.92 $Y=0.83 $X2=0 $Y2=0
cc_402 N_A_806_107#_c_531_n A_962_107# 4.37085e-19 $X=5.005 $Y=1.835 $X2=0 $Y2=0
cc_403 N_VPWR_c_645_n N_A_650_107#_M1013_d 0.0020435f $X=7.37 $Y=3.59 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_645_n N_A_650_107#_c_700_n 0.0221201f $X=7.37 $Y=3.59 $X2=7.92
+ $Y2=4.07
cc_405 N_VPWR_c_642_n N_Q_c_751_n 0.0758093f $X=7.085 $Y=2.62 $X2=0.24 $Y2=4.07
cc_406 N_VPWR_c_645_n N_Q_c_751_n 0.0452076f $X=7.37 $Y=3.59 $X2=0.24 $Y2=4.07
cc_407 N_A_650_107#_c_687_n N_VGND_c_768_n 0.00897815f $X=3.39 $Y=0.83 $X2=4.08
+ $Y2=0.058
cc_408 N_A_650_107#_c_688_n N_VGND_c_768_n 0.0186857f $X=3.39 $Y=0.745 $X2=4.08
+ $Y2=0.058
cc_409 N_A_650_107#_c_688_n N_VGND_c_774_n 0.0317667f $X=3.39 $Y=0.745 $X2=0
+ $Y2=0
cc_410 N_A_650_107#_c_690_n N_VGND_c_774_n 0.0146091f $X=4.06 $Y=1.18 $X2=0
+ $Y2=0
cc_411 N_Q_c_751_n N_VGND_c_772_n 0.0505052f $X=7.885 $Y=0.68 $X2=0 $Y2=0
cc_412 N_Q_c_751_n N_VGND_c_774_n 0.0337877f $X=7.885 $Y=0.68 $X2=0 $Y2=0
cc_413 N_VGND_c_774_n A_962_107# 0.00173335f $X=7.39 $Y=0.48 $X2=0 $Y2=0
