* File: sky130_fd_sc_hvl__dfrbp_1.spice
* Created: Fri Aug 28 09:33:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__dfrbp_1.pex.spice"
.subckt sky130_fd_sc_hvl__dfrbp_1  VNB VPB CLK RESET_B D VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* D	D
* RESET_B	RESET_B
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_CLK_M1020_g N_A_37_107#_M1020_s N_VNB_M1020_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1003 N_A_350_107#_M1003_d N_A_37_107#_M1003_g N_VGND_M1020_d N_VNB_M1020_b NHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1013 A_728_173# N_RESET_B_M1013_g N_VGND_M1013_s N_VNB_M1020_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250000 SB=250007 A=0.21 P=1.84 MULT=1
MM1014 N_A_509_608#_M1014_d N_D_M1014_g A_728_173# N_VNB_M1020_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250001 SB=250006 A=0.21 P=1.84 MULT=1
MM1006 N_A_978_608#_M1006_d N_A_37_107#_M1006_g N_A_509_608#_M1014_d
+ N_VNB_M1020_b NHV L=0.5 W=0.42 AD=0.09345 AS=0.0588 PD=0.865 PS=0.7
+ NRD=44.7792 NRS=0 M=1 R=0.84 SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1028 A_1215_173# N_A_350_107#_M1028_g N_A_978_608#_M1006_d N_VNB_M1020_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.09345 PD=0.63 PS=0.865 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250004 A=0.21 P=1.84 MULT=1
MM1031 A_1357_173# N_A_1176_466#_M1031_g A_1215_173# N_VNB_M1020_b NHV L=0.5
+ W=0.42 AD=0.0483 AS=0.0441 PD=0.65 PS=0.63 NRD=16.2792 NRS=13.566 M=1 R=0.84
+ SA=250003 SB=250003 A=0.21 P=1.84 MULT=1
MM1029 N_VGND_M1029_d N_RESET_B_M1029_g A_1357_173# N_VNB_M1020_b NHV L=0.5
+ W=0.42 AD=0.149531 AS=0.0483 PD=1.04462 PS=0.65 NRD=81.7038 NRS=16.2792 M=1
+ R=0.84 SA=250004 SB=250003 A=0.21 P=1.84 MULT=1
MM1032 N_A_1176_466#_M1032_d N_A_978_608#_M1032_g N_VGND_M1029_d N_VNB_M1020_b
+ NHV L=0.5 W=0.75 AD=0.105 AS=0.267019 PD=1.03 PS=1.86538 NRD=0 NRS=12.1524 M=1
+ R=1.5 SA=250003 SB=250003 A=0.375 P=2.5 MULT=1
MM1016 N_A_1900_107#_M1016_d N_A_350_107#_M1016_g N_A_1176_466#_M1032_d
+ N_VNB_M1020_b NHV L=0.5 W=0.75 AD=0.206346 AS=0.105 PD=1.69231 PS=1.03
+ NRD=15.96 NRS=0 M=1 R=1.5 SA=250004 SB=250002 A=0.375 P=2.5 MULT=1
MM1005 A_2114_107# N_A_37_107#_M1005_g N_A_1900_107#_M1016_d N_VNB_M1020_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.115554 PD=0.63 PS=0.947692 NRD=13.566 NRS=50.2056
+ M=1 R=0.84 SA=250003 SB=250002 A=0.21 P=1.84 MULT=1
MM1007 N_VGND_M1007_d N_A_2122_348#_M1007_g A_2114_107# N_VNB_M1020_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250004 SB=250002 A=0.21 P=1.84 MULT=1
MM1000 A_2412_107# N_RESET_B_M1000_g N_VGND_M1007_d N_VNB_M1020_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250005 SB=250001 A=0.21 P=1.84 MULT=1
MM1001 N_A_2122_348#_M1001_d N_A_1900_107#_M1001_g A_2412_107# N_VNB_M1020_b NHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250005 SB=250000 A=0.21 P=1.84 MULT=1
MM1017 N_Q_N_M1017_d N_A_1900_107#_M1017_g N_VGND_M1017_s N_VNB_M1020_b NHV
+ L=0.5 W=0.75 AD=0.21375 AS=0.21375 PD=2.07 PS=2.07 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1024 N_VGND_M1024_d N_A_1900_107#_M1024_g N_A_2937_443#_M1024_s N_VNB_M1020_b
+ NHV L=0.5 W=0.42 AD=0.0933154 AS=0.1197 PD=0.822051 PS=1.41 NRD=31.2132 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1021 N_Q_M1021_d N_A_2937_443#_M1021_g N_VGND_M1024_d N_VNB_M1020_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.166635 PD=2.03 PS=1.46795 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_CLK_M1004_g N_A_37_107#_M1004_s N_VPB_M1004_b PHV L=0.5
+ W=0.75 AD=0.18375 AS=0.21375 PD=1.24 PS=2.07 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1026 N_A_350_107#_M1026_d N_A_37_107#_M1026_g N_VPWR_M1004_d N_VPB_M1004_b PHV
+ L=0.5 W=0.75 AD=0.21375 AS=0.18375 PD=2.07 PS=1.24 NRD=0 NRS=53.4609 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1018 N_VPWR_M1018_d N_RESET_B_M1018_g N_A_509_608#_M1018_s N_VPB_M1004_b PHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250004 A=0.21 P=1.84 MULT=1
MM1008 N_A_509_608#_M1008_d N_D_M1008_g N_VPWR_M1018_d N_VPB_M1004_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250001
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1030 N_A_978_608#_M1030_d N_A_350_107#_M1030_g N_A_509_608#_M1008_d
+ N_VPB_M1004_b PHV L=0.5 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0
+ M=1 R=0.84 SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1019 A_1134_608# N_A_37_107#_M1019_g N_A_978_608#_M1030_d N_VPB_M1004_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1022 N_VPWR_M1022_d N_A_1176_466#_M1022_g A_1134_608# N_VPB_M1004_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250003 SB=250001 A=0.21 P=1.84 MULT=1
MM1011 N_A_978_608#_M1011_d N_RESET_B_M1011_g N_VPWR_M1022_d N_VPB_M1004_b PHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250004 SB=250000 A=0.21 P=1.84 MULT=1
MM1009 N_A_1176_466#_M1009_d N_A_978_608#_M1009_g N_VPWR_M1009_s N_VPB_M1004_b
+ PHV L=0.5 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=2 SA=250000
+ SB=250003 A=0.5 P=3 MULT=1
MM1002 N_A_1900_107#_M1002_d N_A_37_107#_M1002_g N_A_1176_466#_M1009_d
+ N_VPB_M1004_b PHV L=0.5 W=1 AD=0.233239 AS=0.14 PD=1.96479 PS=1.28 NRD=0 NRS=0
+ M=1 R=2 SA=250001 SB=250002 A=0.5 P=3 MULT=1
MM1015 A_2079_462# N_A_350_107#_M1015_g N_A_1900_107#_M1002_d N_VPB_M1004_b PHV
+ L=0.5 W=0.42 AD=0.04515 AS=0.0979606 PD=0.635 PS=0.825211 NRD=23.8559
+ NRS=52.2958 M=1 R=0.84 SA=250002 SB=250004 A=0.21 P=1.84 MULT=1
MM1027 N_VPWR_M1027_d N_A_2122_348#_M1027_g A_2079_462# N_VPB_M1004_b PHV L=0.5
+ W=0.42 AD=0.0798 AS=0.04515 PD=0.8 PS=0.635 NRD=0 NRS=23.8559 M=1 R=0.84
+ SA=250002 SB=250003 A=0.21 P=1.84 MULT=1
MM1025 N_A_2122_348#_M1025_d N_RESET_B_M1025_g N_VPWR_M1027_d N_VPB_M1004_b PHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.0798 PD=0.7 PS=0.8 NRD=0 NRS=45.458 M=1 R=0.84
+ SA=250003 SB=250002 A=0.21 P=1.84 MULT=1
MM1012 N_VPWR_M1012_d N_A_1900_107#_M1012_g N_A_2122_348#_M1025_d N_VPB_M1004_b
+ PHV L=0.5 W=0.42 AD=0.141291 AS=0.0588 PD=1.00844 PS=0.7 NRD=507.048 NRS=0 M=1
+ R=0.84 SA=250004 SB=250001 A=0.21 P=1.84 MULT=1
MM1023 N_Q_N_M1023_d N_A_1900_107#_M1023_g N_VPWR_M1012_d N_VPB_M1004_b PHV
+ L=0.5 W=1.5 AD=0.4275 AS=0.504609 PD=3.57 PS=3.60156 NRD=0 NRS=0 M=1 R=3
+ SA=250002 SB=250000 A=0.75 P=4 MULT=1
MM1033 N_VPWR_M1033_d N_A_1900_107#_M1033_g N_A_2937_443#_M1033_s N_VPB_M1004_b
+ PHV L=0.5 W=0.75 AD=0.17 AS=0.21375 PD=1.26333 PS=2.07 NRD=29.2803 NRS=0 M=1
+ R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1010 N_Q_M1010_d N_A_2937_443#_M1010_g N_VPWR_M1033_d N_VPB_M1004_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.34 PD=3.57 PS=2.52667 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
DX34_noxref N_VNB_M1020_b N_VPB_M1004_b NWDIODE A=45.396 P=40.12
*
.include "sky130_fd_sc_hvl__dfrbp_1.pxi.spice"
*
.ends
*
*
