* File: sky130_fd_sc_hvl__schmittbuf_1.pex.spice
* Created: Wed Sep  2 09:09:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%VNB 5 7 11 25
r29 7 25 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=0.057
+ $X2=2.64 $Y2=0.058
r30 7 11 0.00134943 $w=5.28e-06 $l=5.7e-08 $layer=MET1_cond $X=2.64 $Y=0.057
+ $X2=2.64 $Y2=0
r31 5 11 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r32 5 11 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%VPB 4 6 14 21
r43 10 21 0.00134943 $w=5.28e-06 $l=5.7e-08 $layer=MET1_cond $X=2.64 $Y=4.07
+ $X2=2.64 $Y2=4.013
r44 10 14 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=4.07
+ $X2=5.04 $Y2=4.07
r45 9 14 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=5.04
+ $Y2=4.07
r46 9 10 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r47 6 21 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=4.012
+ $X2=2.64 $Y2=4.013
r48 4 14 33.0909 $w=1.7e-07 $l=5.08232e-06 $layer=licon1_NTAP_notbjt $count=5
+ $X=0 $Y=3.985 $X2=5.04 $Y2=4.07
r49 4 9 33.0909 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=5
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_117_181# 1 2 7 9 11 13 17 20 23 26
+ 28 36 44 45 46 47
c86 26 0 1.14034e-19 $X=1.47 $Y=1.82
r87 46 47 13.6649 $w=4.08e-07 $l=3.55e-07 $layer=LI1_cond $X=3.855 $Y=1.78
+ $X2=4.21 $Y2=1.78
r88 44 45 7.01511 $w=3.53e-07 $l=1.3e-07 $layer=LI1_cond $X=1.832 $Y=2.46
+ $X2=1.832 $Y2=2.33
r89 40 41 8.14726 $w=2.92e-07 $l=1.95e-07 $layer=LI1_cond $X=1.77 $Y=1.4
+ $X2=1.77 $Y2=1.595
r90 36 47 11.1028 $w=4.08e-07 $l=3.95e-07 $layer=LI1_cond $X=4.605 $Y=1.85
+ $X2=4.21 $Y2=1.85
r91 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.605
+ $Y=1.89 $X2=4.605 $Y2=1.89
r92 33 41 3.56764 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=1.94 $Y=1.595
+ $X2=1.77 $Y2=1.595
r93 33 46 117.995 $w=1.78e-07 $l=1.915e-06 $layer=LI1_cond $X=1.94 $Y=1.595
+ $X2=3.855 $Y2=1.595
r94 28 45 21.2576 $w=1.78e-07 $l=3.45e-07 $layer=LI1_cond $X=1.745 $Y=1.985
+ $X2=1.745 $Y2=2.33
r95 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.47
+ $Y=1.82 $X2=1.47 $Y2=1.82
r96 23 28 8.67714 $w=2.92e-07 $l=1.77059e-07 $layer=LI1_cond $X=1.77 $Y=1.82
+ $X2=1.745 $Y2=1.985
r97 23 41 9.40069 $w=2.92e-07 $l=2.25e-07 $layer=LI1_cond $X=1.77 $Y=1.82
+ $X2=1.77 $Y2=1.595
r98 23 25 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.6 $Y=1.82 $X2=1.47
+ $Y2=1.82
r99 22 26 53.4613 $w=3.4e-07 $l=3.15e-07 $layer=POLY_cond $X=1.155 $Y=1.815
+ $X2=1.47 $Y2=1.815
r100 21 22 11.6485 $w=3.4e-07 $l=2.85e-07 $layer=POLY_cond $X=0.87 $Y=1.815
+ $X2=1.155 $Y2=1.815
r101 20 21 55.3911 $w=4.96e-07 $l=5.7e-07 $layer=POLY_cond $X=0.87 $Y=1.245
+ $X2=0.87 $Y2=1.815
r102 11 37 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=4.615 $Y=1.89
+ $X2=4.605 $Y2=1.89
r103 11 17 97.3754 $w=5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.615 $Y=2.055
+ $X2=4.615 $Y2=2.965
r104 11 13 87.2098 $w=5e-07 $l=8.15e-07 $layer=POLY_cond $X=4.615 $Y=1.725
+ $X2=4.615 $Y2=0.91
r105 7 21 16.388 $w=5e-07 $l=1.86682e-07 $layer=POLY_cond $X=0.905 $Y=1.985
+ $X2=0.87 $Y2=1.815
r106 7 9 75.4392 $w=5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.905 $Y=1.985
+ $X2=0.905 $Y2=2.69
r107 2 44 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.72
+ $Y=2.315 $X2=1.845 $Y2=2.46
r108 1 40 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.65
+ $Y=1.125 $X2=1.775 $Y2=1.4
.ends

.subckt PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A 3 7 9 11 15 17 18 19
c40 19 0 1.14034e-19 $X=3.12 $Y=2.035
c41 11 0 7.68622e-20 $X=2.945 $Y=1.335
c42 3 0 2.80268e-20 $X=2.165 $Y=1.335
r43 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.87
+ $Y=1.94 $X2=2.87 $Y2=1.94
r44 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.19
+ $Y=1.94 $X2=2.19 $Y2=1.94
r45 19 30 9.76647 $w=2.93e-07 $l=2.5e-07 $layer=LI1_cond $X=3.12 $Y=2.002
+ $X2=2.87 $Y2=2.002
r46 18 30 8.98515 $w=2.93e-07 $l=2.3e-07 $layer=LI1_cond $X=2.64 $Y=2.002
+ $X2=2.87 $Y2=2.002
r47 18 26 17.5796 $w=2.93e-07 $l=4.5e-07 $layer=LI1_cond $X=2.64 $Y=2.002
+ $X2=2.19 $Y2=2.002
r48 17 26 1.17198 $w=2.93e-07 $l=3e-08 $layer=LI1_cond $X=2.16 $Y=2.002 $X2=2.19
+ $Y2=2.002
r49 13 15 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.015 $Y=2.14
+ $X2=3.015 $Y2=2.69
r50 9 13 8.99733 $w=3.75e-07 $l=7e-08 $layer=POLY_cond $X=2.945 $Y=1.932
+ $X2=3.015 $Y2=1.932
r51 9 29 9.64 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=2.945 $Y=1.932 $X2=2.87
+ $Y2=1.932
r52 9 11 41.7323 $w=5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.945 $Y=1.725
+ $X2=2.945 $Y2=1.335
r53 5 29 81.6187 $w=3.75e-07 $l=6.35e-07 $layer=POLY_cond $X=2.235 $Y=1.932
+ $X2=2.87 $Y2=1.932
r54 5 25 5.784 $w=3.75e-07 $l=4.5e-08 $layer=POLY_cond $X=2.235 $Y=1.932
+ $X2=2.19 $Y2=1.932
r55 5 7 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.235 $Y=2.14 $X2=2.235
+ $Y2=2.69
r56 1 25 3.21333 $w=3.75e-07 $l=2.5e-08 $layer=POLY_cond $X=2.165 $Y=1.932
+ $X2=2.19 $Y2=1.932
r57 1 3 41.7323 $w=5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.165 $Y=1.725 $X2=2.165
+ $Y2=1.335
.ends

.subckt PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_78_463# 1 2 9 12 13 15 19
r31 13 15 49.6831 $w=2.23e-07 $l=9.7e-07 $layer=LI1_cond $X=0.875 $Y=0.682
+ $X2=1.845 $Y2=0.682
r32 12 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=2.165
+ $X2=0.79 $Y2=2.25
r33 11 13 6.9898 $w=2.25e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.79 $Y=0.795
+ $X2=0.875 $Y2=0.682
r34 11 12 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=0.79 $Y=0.795
+ $X2=0.79 $Y2=2.165
r35 7 19 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.555 $Y=2.25
+ $X2=0.79 $Y2=2.25
r36 7 9 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.555 $Y=2.335
+ $X2=0.555 $Y2=2.46
r37 2 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.39
+ $Y=2.315 $X2=0.515 $Y2=2.46
r38 1 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.72
+ $Y=0.535 $X2=1.845 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_64_207# 1 2 8 9 10 11 13 20
r32 11 15 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.405 $Y=1.89
+ $X2=0.17 $Y2=1.89
r33 11 13 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=0.405 $Y=1.805
+ $X2=0.405 $Y2=1.255
r34 9 20 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.74 $Y=3.57
+ $X2=0.905 $Y2=3.57
r35 9 10 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=0.74 $Y=3.57
+ $X2=0.255 $Y2=3.57
r36 8 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=3.485
+ $X2=0.255 $Y2=3.57
r37 7 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.17 $Y=1.975
+ $X2=0.17 $Y2=1.89
r38 7 8 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=0.17 $Y=1.975
+ $X2=0.17 $Y2=3.485
r39 2 20 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.78
+ $Y=3.425 $X2=0.905 $Y2=3.57
r40 1 13 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=0.32
+ $Y=1.035 $X2=0.445 $Y2=1.255
.ends

.subckt PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_231_463# 1 2 9 11 12 15
r25 13 15 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=2.625 $Y=3.235
+ $X2=2.625 $Y2=2.45
r26 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.46 $Y=3.32
+ $X2=2.625 $Y2=3.235
r27 11 12 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=2.46 $Y=3.32 $X2=1.46
+ $Y2=3.32
r28 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.33 $Y=3.235
+ $X2=1.46 $Y2=3.32
r29 7 9 34.3517 $w=2.58e-07 $l=7.75e-07 $layer=LI1_cond $X=1.33 $Y=3.235
+ $X2=1.33 $Y2=2.46
r30 2 15 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=2.485
+ $Y=2.315 $X2=2.625 $Y2=2.45
r31 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.155
+ $Y=2.315 $X2=1.295 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%VPWR 1 4 12 15
r27 13 15 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=3.31 $Y=3.63
+ $X2=4.39 $Y2=3.63
r28 12 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.39 $Y=3.56
+ $X2=4.39 $Y2=3.56
r29 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.31 $Y=3.56
+ $X2=3.31 $Y2=3.56
r30 10 12 3.23179 $w=1.359e-06 $l=3.6e-07 $layer=LI1_cond $X=3.85 $Y=3.2
+ $X2=3.85 $Y2=3.56
r31 7 10 6.82266 $w=1.359e-06 $l=7.6e-07 $layer=LI1_cond $X=3.85 $Y=2.44
+ $X2=3.85 $Y2=3.2
r32 4 13 0.257217 $w=3.7e-07 $l=6.7e-07 $layer=MET1_cond $X=2.64 $Y=3.63
+ $X2=3.31 $Y2=3.63
r33 1 12 600 $w=1.7e-07 $l=1.73599e-06 $layer=licon1_PDIFF $count=1 $X=2.56
+ $Y=3.425 $X2=4.225 $Y2=3.57
r34 1 10 600 $w=1.7e-07 $l=1.77394e-06 $layer=licon1_PDIFF $count=1 $X=2.56
+ $Y=3.425 $X2=4.225 $Y2=3.2
r35 1 7 300 $w=1.7e-07 $l=2.10054e-06 $layer=licon1_PDIFF $count=2 $X=2.56
+ $Y=3.425 $X2=4.225 $Y2=2.44
r36 1 7 150 $w=1.7e-07 $l=1.68708e-06 $layer=licon1_PDIFF $count=4 $X=2.56
+ $Y=3.425 $X2=3.825 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%X 1 2 7 8 9 10 11 12 13 22
r14 13 40 13.9325 $w=3.33e-07 $l=4.05e-07 $layer=LI1_cond $X=5.027 $Y=3.145
+ $X2=5.027 $Y2=3.55
r15 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=5.027 $Y=2.775
+ $X2=5.027 $Y2=3.145
r16 11 12 13.9325 $w=3.33e-07 $l=4.05e-07 $layer=LI1_cond $X=5.027 $Y=2.37
+ $X2=5.027 $Y2=2.775
r17 10 11 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=5.027 $Y=2.035
+ $X2=5.027 $Y2=2.37
r18 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=5.027 $Y=1.665
+ $X2=5.027 $Y2=2.035
r19 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=5.027 $Y=1.295
+ $X2=5.027 $Y2=1.665
r20 7 8 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=5.027 $Y=0.925
+ $X2=5.027 $Y2=1.295
r21 7 22 8.42831 $w=3.33e-07 $l=2.45e-07 $layer=LI1_cond $X=5.027 $Y=0.925
+ $X2=5.027 $Y2=0.68
r22 2 40 300 $w=1.7e-07 $l=1.40326e-06 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=2.215 $X2=5.005 $Y2=3.55
r23 2 11 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=2.215 $X2=5.005 $Y2=2.37
r24 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.865
+ $Y=0.535 $X2=5.005 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%A_217_207# 1 2 7 9 14
c26 7 0 7.68622e-20 $X=2.39 $Y=1.06
r27 14 17 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.555 $Y=1.06
+ $X2=2.555 $Y2=1.25
r28 9 12 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.225 $Y=1.06
+ $X2=1.225 $Y2=1.245
r29 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=1.06 $X2=1.225
+ $Y2=1.06
r30 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=1.06
+ $X2=2.555 $Y2=1.06
r31 7 8 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=2.39 $Y=1.06 $X2=1.39
+ $Y2=1.06
r32 2 17 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=1.125 $X2=2.555 $Y2=1.25
r33 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=1.035 $X2=1.225 $Y2=1.245
.ends

.subckt PM_SKY130_FD_SC_HVL__SCHMITTBUF_1%VGND 1 4 7 11
c23 11 0 2.80268e-20 $X=4.495 $Y=0.51
r24 8 11 0.460686 $w=3.7e-07 $l=1.2e-06 $layer=MET1_cond $X=3.295 $Y=0.44
+ $X2=4.495 $Y2=0.44
r25 7 13 2.18146 $w=1.508e-06 $l=2.7e-07 $layer=LI1_cond $X=3.875 $Y=0.51
+ $X2=3.875 $Y2=0.78
r26 7 11 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.495 $Y=0.51
+ $X2=4.495 $Y2=0.51
r27 7 8 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.295 $Y=0.51
+ $X2=3.295 $Y2=0.51
r28 4 8 0.251458 $w=3.7e-07 $l=6.55e-07 $layer=MET1_cond $X=2.64 $Y=0.44
+ $X2=3.295 $Y2=0.44
r29 1 13 60.6667 $w=1.7e-07 $l=1.72315e-06 $layer=licon1_NDIFF $count=3 $X=2.62
+ $Y=0.535 $X2=4.225 $Y2=0.78
r30 1 13 60.6667 $w=1.7e-07 $l=9.0424e-07 $layer=licon1_NDIFF $count=3 $X=2.62
+ $Y=0.535 $X2=3.41 $Y2=0.78
.ends

