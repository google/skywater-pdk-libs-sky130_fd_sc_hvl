* File: sky130_fd_sc_hvl__sdfxbp_1.spice
* Created: Wed Sep  2 09:10:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__sdfxbp_1.pex.spice"
.subckt sky130_fd_sc_hvl__sdfxbp_1  VNB VPB SCE SCD D CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* D	D
* SCD	SCD
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1028 N_VGND_M1028_d N_SCE_M1028_g N_A_30_515#_M1028_s N_VNB_M1028_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1019 A_425_107# N_SCD_M1019_g N_VGND_M1028_d N_VNB_M1028_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84 SA=250001
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1020 N_A_567_107#_M1020_d N_SCE_M1020_g A_425_107# N_VNB_M1028_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1013 A_723_107# N_A_30_515#_M1013_g N_A_567_107#_M1020_d N_VNB_M1028_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1014 N_VGND_M1014_d N_D_M1014_g A_723_107# N_VNB_M1028_b NHV L=0.5 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250003
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1003 N_VGND_M1003_d N_A_1124_81#_M1003_g N_A_1067_107#_M1003_s N_VNB_M1028_b
+ NHV L=0.5 W=0.75 AD=0.252212 AS=0.21375 PD=1.79487 PS=2.07 NRD=12.1524 NRS=0
+ M=1 R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1012 N_A_1454_173#_M1012_d N_A_1067_107#_M1012_g N_VGND_M1003_d N_VNB_M1028_b
+ NHV L=0.5 W=0.42 AD=0.1197 AS=0.141238 PD=1.41 PS=1.00513 NRD=0 NRS=76.3458
+ M=1 R=0.84 SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1017 N_A_1124_81#_M1017_d N_A_1570_457#_M1017_g N_A_567_107#_M1017_s
+ N_VNB_M1028_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1030 N_A_1454_173#_M1030_d N_A_1726_453#_M1030_g N_A_1124_81#_M1017_d
+ N_VNB_M1028_b NHV L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0
+ M=1 R=0.84 SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1004 N_VGND_M1004_d N_A_1570_457#_M1004_g N_A_1726_453#_M1004_s N_VNB_M1028_b
+ NHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1026 N_A_1570_457#_M1026_d N_CLK_M1026_g N_VGND_M1004_d N_VNB_M1028_b NHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1005 N_A_2518_445#_M1005_d N_A_1726_453#_M1005_g N_A_1067_107#_M1005_s
+ N_VNB_M1028_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1029 A_2747_173# N_A_1570_457#_M1029_g N_A_2518_445#_M1005_d N_VNB_M1028_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250001 SB=250002 A=0.21 P=1.84 MULT=1
MM1031 N_VGND_M1031_d N_A_2789_147#_M1031_g A_2747_173# N_VNB_M1028_b NHV L=0.5
+ W=0.42 AD=0.0933154 AS=0.0441 PD=0.822051 PS=0.63 NRD=31.2132 NRS=13.566 M=1
+ R=0.84 SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1006 N_A_2789_147#_M1006_d N_A_2518_445#_M1006_g N_VGND_M1031_d N_VNB_M1028_b
+ NHV L=0.5 W=0.75 AD=0.21375 AS=0.166635 PD=2.07 PS=1.46795 NRD=0 NRS=0 M=1
+ R=1.5 SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1010 N_VGND_M1010_d N_A_2789_147#_M1010_g N_Q_M1010_s N_VNB_M1028_b NHV L=0.5
+ W=0.75 AD=0.166635 AS=0.21375 PD=1.46795 PS=2.07 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1032 N_A_3531_107#_M1032_d N_A_2789_147#_M1032_g N_VGND_M1010_d N_VNB_M1028_b
+ NHV L=0.5 W=0.42 AD=0.1197 AS=0.0933154 PD=1.41 PS=0.822051 NRD=0 NRS=31.2132
+ M=1 R=0.84 SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1011 N_Q_N_M1011_d N_A_3531_107#_M1011_g N_VGND_M1011_s N_VNB_M1028_b NHV
+ L=0.5 W=0.75 AD=0.21375 AS=0.21375 PD=2.07 PS=2.07 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1022 N_VPWR_M1022_d N_SCE_M1022_g N_A_30_515#_M1022_s N_VPB_M1022_b PHV L=0.5
+ W=0.42 AD=0.1197 AS=0.1113 PD=1.41 PS=1.37 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1000 N_VPWR_M1000_d N_SCD_M1000_g N_A_268_659#_M1000_s N_VPB_M1022_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1018 N_A_581_659#_M1018_d N_SCE_M1018_g N_VPWR_M1000_d N_VPB_M1022_b PHV L=0.5
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250001
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1016 N_A_567_107#_M1016_d N_A_30_515#_M1016_g N_A_268_659#_M1016_s
+ N_VPB_M1022_b PHV L=0.5 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1007 N_A_581_659#_M1007_d N_D_M1007_g N_A_567_107#_M1016_d N_VPB_M1022_b PHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1035 N_VPWR_M1035_d N_A_1124_81#_M1035_g N_A_1067_107#_M1035_s N_VPB_M1022_b
+ PHV L=0.5 W=1 AD=0.351549 AS=0.265 PD=2.52817 PS=2.53 NRD=0 NRS=0 M=1 R=2
+ SA=250000 SB=250001 A=0.5 P=3 MULT=1
MM1001 A_1528_579# N_A_1067_107#_M1001_g N_VPWR_M1035_d N_VPB_M1022_b PHV L=0.5
+ W=0.42 AD=0.0441 AS=0.147651 PD=0.63 PS=1.06183 NRD=22.729 NRS=134.846 M=1
+ R=0.84 SA=250001 SB=250002 A=0.21 P=1.84 MULT=1
MM1002 N_A_1124_81#_M1002_d N_A_1570_457#_M1002_g A_1528_579# N_VPB_M1022_b PHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1027 N_A_567_107#_M1027_d N_A_1726_453#_M1027_g N_A_1124_81#_M1002_d
+ N_VPB_M1022_b PHV L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0
+ M=1 R=0.84 SA=250003 SB=250000 A=0.21 P=1.84 MULT=1
MM1024 N_VPWR_M1024_d N_A_1570_457#_M1024_g N_A_1726_453#_M1024_s N_VPB_M1022_b
+ PHV L=0.5 W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1008 N_A_1570_457#_M1008_d N_CLK_M1008_g N_VPWR_M1024_d N_VPB_M1022_b PHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1034 N_A_2518_445#_M1034_d N_A_1726_453#_M1034_g N_A_2365_445#_M1034_s
+ N_VPB_M1022_b PHV L=0.5 W=0.42 AD=0.0920451 AS=0.1113 PD=0.81338 PS=1.37
+ NRD=43.1851 NRS=0 M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1025 N_A_1067_107#_M1025_d N_A_1570_457#_M1025_g N_A_2518_445#_M1034_d
+ N_VPB_M1022_b PHV L=0.5 W=1 AD=0.285 AS=0.219155 PD=2.57 PS=1.93662 NRD=0
+ NRS=0 M=1 R=2 SA=250000 SB=250000 A=0.5 P=3 MULT=1
MM1023 N_VPWR_M1023_d N_A_2789_147#_M1023_g N_A_2365_445#_M1023_s N_VPB_M1022_b
+ PHV L=0.5 W=0.42 AD=0.0920451 AS=0.1113 PD=0.81338 PS=1.37 NRD=43.1851 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1015 N_A_2789_147#_M1015_d N_A_2518_445#_M1015_g N_VPWR_M1023_d N_VPB_M1022_b
+ PHV L=0.5 W=1 AD=0.265 AS=0.219155 PD=2.53 PS=1.93662 NRD=0 NRS=0 M=1 R=2
+ SA=250000 SB=250000 A=0.5 P=3 MULT=1
MM1009 N_VPWR_M1009_d N_A_2789_147#_M1009_g N_Q_M1009_s N_VPB_M1022_b PHV L=0.5
+ W=1.5 AD=0.32 AS=0.3975 PD=2.5 PS=3.53 NRD=0 NRS=0 M=1 R=3 SA=250000 SB=250000
+ A=0.75 P=4 MULT=1
MM1033 N_A_3531_107#_M1033_d N_A_2789_147#_M1033_g N_VPWR_M1009_d N_VPB_M1022_b
+ PHV L=0.5 W=0.75 AD=0.19875 AS=0.16 PD=2.03 PS=1.25 NRD=0 NRS=24.1806 M=1
+ R=1.5 SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1021 N_Q_N_M1021_d N_A_3531_107#_M1021_g N_VPWR_M1021_s N_VPB_M1022_b PHV
+ L=0.5 W=1.5 AD=0.4275 AS=0.4275 PD=3.57 PS=3.57 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
DX36_noxref N_VNB_M1028_b N_VPB_M1022_b NWDIODE A=53.32 P=46.22
*
.include "sky130_fd_sc_hvl__sdfxbp_1.pxi.spice"
*
.ends
*
*
