* File: sky130_fd_sc_hvl__and3_1.pex.spice
* Created: Fri Aug 28 09:32:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__AND3_1%VNB 5 7 11 25
r20 7 25 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=0.057
+ $X2=1.92 $Y2=0.058
r21 7 11 0.00185547 $w=3.84e-06 $l=5.7e-08 $layer=MET1_cond $X=1.92 $Y=0.057
+ $X2=1.92 $Y2=0
r22 5 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r23 5 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__AND3_1%VPB 4 6 14 21
r29 10 21 0.00185547 $w=3.84e-06 $l=5.7e-08 $layer=MET1_cond $X=1.92 $Y=4.07
+ $X2=1.92 $Y2=4.013
r30 10 14 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=4.07
+ $X2=3.6 $Y2=4.07
r31 9 14 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=3.6
+ $Y2=4.07
r32 9 10 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r33 6 21 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=4.012
+ $X2=1.92 $Y2=4.013
r34 4 14 45.5 $w=1.7e-07 $l=3.64225e-06 $layer=licon1_NTAP_notbjt $count=4 $X=0
+ $Y=3.985 $X2=3.6 $Y2=4.07
r35 4 9 45.5 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=4 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__AND3_1%A 3 7 8 9 13 15
r22 13 16 32.3893 $w=5.7e-07 $l=3.35e-07 $layer=POLY_cond $X=0.72 $Y=1.56
+ $X2=0.72 $Y2=1.895
r23 13 15 16.4322 $w=5.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.72 $Y=1.56
+ $X2=0.72 $Y2=1.395
r24 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.56 $X2=0.77 $Y2=1.56
r25 9 14 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.77 $Y=1.295
+ $X2=0.77 $Y2=1.56
r26 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.77 $Y=0.925 $X2=0.77
+ $Y2=1.295
r27 7 15 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.755 $Y=1.075 $X2=0.755
+ $Y2=1.395
r28 3 16 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=0.685 $Y=2.795 $X2=0.685
+ $Y2=1.895
.ends

.subckt PM_SKY130_FD_SC_HVL__AND3_1%B 1 2 6 10 12
r22 9 12 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.465 $Y=2.26
+ $X2=1.465 $Y2=2.795
r23 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.4 $Y=2.26
+ $X2=1.4 $Y2=2.26
r24 6 9 126.802 $w=5e-07 $l=1.185e-06 $layer=POLY_cond $X=1.465 $Y=1.075
+ $X2=1.465 $Y2=2.26
r25 2 10 7.3171 $w=3.13e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=2.332 $X2=1.4
+ $Y2=2.332
r26 1 2 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=2.332 $X2=1.2
+ $Y2=2.332
.ends

.subckt PM_SKY130_FD_SC_HVL__AND3_1%C 3 6 8 10 12 21 23
r35 21 24 32.3893 $w=5.7e-07 $l=3.35e-07 $layer=POLY_cond $X=2.21 $Y=1.56
+ $X2=2.21 $Y2=1.895
r36 21 23 16.4322 $w=5.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.56
+ $X2=2.21 $Y2=1.395
r37 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.09
+ $Y=1.56 $X2=2.09 $Y2=1.56
r38 12 22 1.0027 $w=8.33e-07 $l=7e-08 $layer=LI1_cond $X=2.16 $Y=1.227 $X2=2.09
+ $Y2=1.227
r39 10 22 5.87296 $w=8.33e-07 $l=4.1e-07 $layer=LI1_cond $X=1.68 $Y=1.227
+ $X2=2.09 $Y2=1.227
r40 8 10 6.87566 $w=8.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.227 $X2=1.68
+ $Y2=1.227
r41 6 24 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=2.245 $Y=2.795 $X2=2.245
+ $Y2=1.895
r42 3 23 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.175 $Y=1.075 $X2=2.175
+ $Y2=1.395
.ends

.subckt PM_SKY130_FD_SC_HVL__AND3_1%A_30_517# 1 2 3 12 16 20 24 26 30 32 34 35
+ 37 38
r67 38 44 25.8045 $w=5.35e-07 $l=2.55e-07 $layer=POLY_cond $X=3.157 $Y=1.83
+ $X2=3.157 $Y2=2.085
r68 38 43 41.8054 $w=5.35e-07 $l=4.15e-07 $layer=POLY_cond $X=3.157 $Y=1.83
+ $X2=3.157 $Y2=1.415
r69 37 40 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.075 $Y=1.83 $X2=3.075
+ $Y2=1.91
r70 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.075
+ $Y=1.83 $X2=3.075 $Y2=1.83
r71 33 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.02 $Y=1.91
+ $X2=1.895 $Y2=1.91
r72 32 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.91 $Y=1.91
+ $X2=3.075 $Y2=1.91
r73 32 33 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.91 $Y=1.91
+ $X2=2.02 $Y2=1.91
r74 28 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=1.995
+ $X2=1.895 $Y2=1.91
r75 28 30 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=1.895 $Y=1.995
+ $X2=1.895 $Y2=2.795
r76 27 34 3.08518 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.425 $Y=1.91
+ $X2=0.277 $Y2=1.91
r77 26 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.77 $Y=1.91
+ $X2=1.895 $Y2=1.91
r78 26 27 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=1.77 $Y=1.91
+ $X2=0.425 $Y2=1.91
r79 22 34 3.43356 $w=2.72e-07 $l=9.53677e-08 $layer=LI1_cond $X=0.255 $Y=1.995
+ $X2=0.277 $Y2=1.91
r80 22 24 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=0.255 $Y=1.995
+ $X2=0.255 $Y2=2.795
r81 18 34 3.43356 $w=2.72e-07 $l=8.5e-08 $layer=LI1_cond $X=0.277 $Y=1.825
+ $X2=0.277 $Y2=1.91
r82 18 20 29.2994 $w=2.93e-07 $l=7.5e-07 $layer=LI1_cond $X=0.277 $Y=1.825
+ $X2=0.277 $Y2=1.075
r83 16 43 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.175 $Y=0.91
+ $X2=3.175 $Y2=1.415
r84 12 44 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.14 $Y=2.965 $X2=3.14
+ $Y2=2.085
r85 3 30 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.715
+ $Y=2.585 $X2=1.855 $Y2=2.795
r86 2 24 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.585 $X2=0.295 $Y2=2.795
r87 1 20 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.195
+ $Y=0.865 $X2=0.34 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__AND3_1%VPWR 1 2 7 10 19 29
r30 27 29 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.315 $Y=3.63
+ $X2=3.035 $Y2=3.63
r31 26 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.035 $Y=3.59
+ $X2=3.035 $Y2=3.59
r32 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.315 $Y=3.59
+ $X2=2.315 $Y2=3.59
r33 24 26 5.32947 $w=9.48e-07 $l=4.15e-07 $layer=LI1_cond $X=2.675 $Y=3.175
+ $X2=2.675 $Y2=3.59
r34 22 24 5.39368 $w=9.48e-07 $l=4.2e-07 $layer=LI1_cond $X=2.675 $Y=2.755
+ $X2=2.675 $Y2=3.175
r35 19 22 5.32947 $w=9.48e-07 $l=4.15e-07 $layer=LI1_cond $X=2.675 $Y=2.34
+ $X2=2.675 $Y2=2.755
r36 14 16 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.675 $Y=3.63
+ $X2=1.395 $Y2=3.63
r37 13 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.395 $Y=3.59
+ $X2=1.395 $Y2=3.59
r38 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.675 $Y=3.59
+ $X2=0.675 $Y2=3.59
r39 10 13 9.95263 $w=9.48e-07 $l=7.75e-07 $layer=LI1_cond $X=1.035 $Y=2.815
+ $X2=1.035 $Y2=3.59
r40 7 27 0.151643 $w=3.7e-07 $l=3.95e-07 $layer=MET1_cond $X=1.92 $Y=3.63
+ $X2=2.315 $Y2=3.63
r41 7 16 0.20155 $w=3.7e-07 $l=5.25e-07 $layer=MET1_cond $X=1.92 $Y=3.63
+ $X2=1.395 $Y2=3.63
r42 2 24 300 $w=1.7e-07 $l=7.06081e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=2.585 $X2=2.75 $Y2=3.175
r43 2 22 600 $w=1.7e-07 $l=3.29204e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=2.585 $X2=2.75 $Y2=2.755
r44 2 19 600 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=2.585 $X2=2.75 $Y2=2.34
r45 1 10 600 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=2.585 $X2=1.075 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HVL__AND3_1%X 1 2 7 8 9 10 11 12 13 24 36
r18 34 36 1.81098 $w=3.48e-07 $l=5.5e-08 $layer=LI1_cond $X=3.54 $Y=2.35
+ $X2=3.54 $Y2=2.405
r19 13 43 14.6525 $w=3.48e-07 $l=4.45e-07 $layer=LI1_cond $X=3.54 $Y=3.145
+ $X2=3.54 $Y2=3.59
r20 12 13 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.54 $Y=2.775
+ $X2=3.54 $Y2=3.145
r21 11 34 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=3.54 $Y=2.335
+ $X2=3.54 $Y2=2.35
r22 11 46 5.48937 $w=3.48e-07 $l=1.6e-07 $layer=LI1_cond $X=3.54 $Y=2.335
+ $X2=3.54 $Y2=2.175
r23 11 12 11.6891 $w=3.48e-07 $l=3.55e-07 $layer=LI1_cond $X=3.54 $Y=2.42
+ $X2=3.54 $Y2=2.775
r24 11 36 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=3.54 $Y=2.42
+ $X2=3.54 $Y2=2.405
r25 10 46 5.2899 $w=3.03e-07 $l=1.4e-07 $layer=LI1_cond $X=3.562 $Y=2.035
+ $X2=3.562 $Y2=2.175
r26 9 10 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=3.562 $Y=1.665
+ $X2=3.562 $Y2=2.035
r27 8 9 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=3.562 $Y=1.295
+ $X2=3.562 $Y2=1.665
r28 7 8 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=3.562 $Y=0.925
+ $X2=3.562 $Y2=1.295
r29 7 24 9.25733 $w=3.03e-07 $l=2.45e-07 $layer=LI1_cond $X=3.562 $Y=0.925
+ $X2=3.562 $Y2=0.68
r30 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=3.39
+ $Y=2.215 $X2=3.53 $Y2=2.34
r31 2 43 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=3.39
+ $Y=2.215 $X2=3.53 $Y2=3.59
r32 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.425
+ $Y=0.535 $X2=3.565 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__AND3_1%VGND 1 4 7 8
r20 11 13 7.42906 $w=8.03e-07 $l=5e-07 $layer=LI1_cond $X=2.837 $Y=0.66
+ $X2=2.837 $Y2=1.16
r21 7 11 2.67446 $w=8.03e-07 $l=1.8e-07 $layer=LI1_cond $X=2.837 $Y=0.48
+ $X2=2.837 $Y2=0.66
r22 7 8 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.1 $Y=0.48 $X2=3.1
+ $Y2=0.48
r23 4 8 0.453008 $w=3.7e-07 $l=1.18e-06 $layer=MET1_cond $X=1.92 $Y=0.44 $X2=3.1
+ $Y2=0.44
r24 1 13 182 $w=1.7e-07 $l=4.85592e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.865 $X2=2.785 $Y2=1.16
r25 1 11 182 $w=1.7e-07 $l=4.50999e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.865 $X2=2.785 $Y2=0.66
.ends

