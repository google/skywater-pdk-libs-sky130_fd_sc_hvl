* File: sky130_fd_sc_hvl__decap_8.pex.spice
* Created: Fri Aug 28 09:33:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__DECAP_8%VNB 5 7 11 25
r12 7 25 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=0.057
+ $X2=1.92 $Y2=0.058
r13 7 11 0.00185547 $w=3.84e-06 $l=5.7e-08 $layer=MET1_cond $X=1.92 $Y=0.057
+ $X2=1.92 $Y2=0
r14 5 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r15 5 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__DECAP_8%VPB 4 6 14 21
r18 10 21 0.00185547 $w=3.84e-06 $l=5.7e-08 $layer=MET1_cond $X=1.92 $Y=4.07
+ $X2=1.92 $Y2=4.013
r19 10 14 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=4.07
+ $X2=3.6 $Y2=4.07
r20 9 14 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=3.6
+ $Y2=4.07
r21 9 10 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r22 6 21 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=4.012
+ $X2=1.92 $Y2=4.013
r23 4 14 45.5 $w=1.7e-07 $l=3.64225e-06 $layer=licon1_NTAP_notbjt $count=4 $X=0
+ $Y=3.985 $X2=3.6 $Y2=4.07
r24 4 9 45.5 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=4 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__DECAP_8%VGND 1 12 17 22 23 27 28 30 50
r47 47 50 3.111 $w=9.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.965 $Y=0.86
+ $X2=3.22 $Y2=0.86
r48 45 47 9.577 $w=9.98e-07 $l=7.85e-07 $layer=LI1_cond $X=2.18 $Y=0.86
+ $X2=2.965 $Y2=0.86
r49 44 45 2.928 $w=9.98e-07 $l=2.4e-07 $layer=LI1_cond $X=1.94 $Y=0.86 $X2=2.18
+ $Y2=0.86
r50 42 44 12.688 $w=9.98e-07 $l=1.04e-06 $layer=LI1_cond $X=0.9 $Y=0.86 $X2=1.94
+ $Y2=0.86
r51 41 47 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.965 $Y=0.475
+ $X2=2.965 $Y2=0.475
r52 40 42 0.854 $w=9.98e-07 $l=7e-08 $layer=LI1_cond $X=0.83 $Y=0.86 $X2=0.9
+ $Y2=0.86
r53 40 41 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.83 $Y=0.475
+ $X2=0.83 $Y2=0.475
r54 37 40 2.074 $w=9.98e-07 $l=1.7e-07 $layer=LI1_cond $X=0.66 $Y=0.86 $X2=0.83
+ $Y2=0.86
r55 30 41 0.00113932 $w=3.84e-06 $l=3.5e-08 $layer=MET1_cond $X=1.92 $Y=0.44
+ $X2=1.92 $Y2=0.475
r56 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.18
+ $Y=1.86 $X2=2.18 $Y2=1.86
r57 25 45 7.34451 $w=3.3e-07 $l=5e-07 $layer=LI1_cond $X=2.18 $Y=1.36 $X2=2.18
+ $Y2=0.86
r58 25 27 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.18 $Y=1.36 $X2=2.18
+ $Y2=1.86
r59 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.9
+ $Y=1.86 $X2=0.9 $Y2=1.86
r60 20 42 7.34451 $w=3.3e-07 $l=5e-07 $layer=LI1_cond $X=0.9 $Y=1.36 $X2=0.9
+ $Y2=0.86
r61 20 22 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.9 $Y=1.36 $X2=0.9
+ $Y2=1.86
r62 18 28 124.152 $w=3.3e-07 $l=7.1e-07 $layer=POLY_cond $X=2.18 $Y=2.57
+ $X2=2.18 $Y2=1.86
r63 17 18 57.2398 $w=1e-06 $l=6.3e-07 $layer=POLY_cond $X=2.515 $Y=3.2 $X2=2.515
+ $Y2=2.57
r64 13 23 124.152 $w=3.3e-07 $l=7.1e-07 $layer=POLY_cond $X=0.9 $Y=2.57 $X2=0.9
+ $Y2=1.86
r65 12 13 57.2398 $w=1e-06 $l=6.3e-07 $layer=POLY_cond $X=1.235 $Y=3.2 $X2=1.235
+ $Y2=2.57
r66 1 50 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=3.08
+ $Y=0.59 $X2=3.22 $Y2=0.805
r67 1 44 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=1.8 $Y=0.59
+ $X2=1.94 $Y2=0.805
r68 1 37 91 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=2 $X=1.8 $Y=0.59
+ $X2=0.66 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_HVL__DECAP_8%VPWR 1 10 12 13 15 18 19 23 24 26 46 48
r45 45 48 2.62243 $w=1.068e-06 $l=2.3e-07 $layer=LI1_cond $X=2.925 $Y=3.215
+ $X2=3.155 $Y2=3.215
r46 45 46 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.925 $Y=3.64
+ $X2=2.925 $Y2=3.64
r47 43 45 0.114019 $w=1.068e-06 $l=1e-08 $layer=LI1_cond $X=2.915 $Y=3.215
+ $X2=2.925 $Y2=3.215
r48 41 43 11.8579 $w=1.068e-06 $l=1.04e-06 $layer=LI1_cond $X=1.875 $Y=3.215
+ $X2=2.915 $Y2=3.215
r49 39 41 2.73645 $w=1.068e-06 $l=2.4e-07 $layer=LI1_cond $X=1.635 $Y=3.215
+ $X2=1.875 $Y2=3.215
r50 37 39 9.63458 $w=1.068e-06 $l=8.45e-07 $layer=LI1_cond $X=0.79 $Y=3.215
+ $X2=1.635 $Y2=3.215
r51 37 38 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.79 $Y=3.64
+ $X2=0.79 $Y2=3.64
r52 33 37 2.33738 $w=1.068e-06 $l=2.05e-07 $layer=LI1_cond $X=0.585 $Y=3.215
+ $X2=0.79 $Y2=3.215
r53 26 46 0.385825 $w=3.7e-07 $l=1.005e-06 $layer=MET1_cond $X=1.92 $Y=3.63
+ $X2=2.925 $Y2=3.63
r54 26 38 0.433813 $w=3.7e-07 $l=1.13e-06 $layer=MET1_cond $X=1.92 $Y=3.63
+ $X2=0.79 $Y2=3.63
r55 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=1.86 $X2=2.915 $Y2=1.86
r56 21 43 7.77329 $w=3.3e-07 $l=5.35e-07 $layer=LI1_cond $X=2.915 $Y=2.68
+ $X2=2.915 $Y2=3.215
r57 21 23 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=2.915 $Y=2.68
+ $X2=2.915 $Y2=1.86
r58 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.635
+ $Y=1.86 $X2=1.635 $Y2=1.86
r59 16 39 7.77329 $w=3.3e-07 $l=5.35e-07 $layer=LI1_cond $X=1.635 $Y=2.68
+ $X2=1.635 $Y2=3.215
r60 16 18 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=1.635 $Y=2.68
+ $X2=1.635 $Y2=1.86
r61 13 24 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=2.915 $Y=1.47
+ $X2=2.915 $Y2=1.86
r62 13 15 47.6333 $w=1e-06 $l=5.4631e-07 $layer=POLY_cond $X=2.915 $Y=1.47
+ $X2=2.829 $Y2=0.965
r63 10 19 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=1.635 $Y=1.47
+ $X2=1.635 $Y2=1.86
r64 10 12 47.6333 $w=1e-06 $l=5.4631e-07 $layer=POLY_cond $X=1.635 $Y=1.47
+ $X2=1.549 $Y2=0.965
r65 1 48 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.015
+ $Y=2.7 $X2=3.155 $Y2=3.555
r66 1 48 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.015
+ $Y=2.7 $X2=3.155 $Y2=2.845
r67 1 41 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.735
+ $Y=2.7 $X2=1.875 $Y2=3.555
r68 1 41 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.735
+ $Y=2.7 $X2=1.875 $Y2=2.845
r69 1 33 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.735
+ $Y=2.7 $X2=0.585 $Y2=3.555
r70 1 33 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.735
+ $Y=2.7 $X2=0.585 $Y2=2.845
.ends

