* File: sky130_fd_sc_hvl__inv_8.spice
* Created: Fri Aug 28 09:36:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__inv_8.pex.spice"
.subckt sky130_fd_sc_hvl__inv_8  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s N_VNB_M1000_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000 SB=250006
+ A=0.375 P=2.5 MULT=1
MM1001 N_Y_M1000_d N_A_M1001_g N_VGND_M1001_s N_VNB_M1000_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250001 SB=250005
+ A=0.375 P=2.5 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1001_s N_VNB_M1000_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250002 SB=250004
+ A=0.375 P=2.5 MULT=1
MM1005 N_Y_M1002_d N_A_M1005_g N_VGND_M1005_s N_VNB_M1000_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250002 SB=250003
+ A=0.375 P=2.5 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VGND_M1005_s N_VNB_M1000_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250003 SB=250003
+ A=0.375 P=2.5 MULT=1
MM1008 N_Y_M1006_d N_A_M1008_g N_VGND_M1008_s N_VNB_M1000_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.1575 PD=1.03 PS=1.17 NRD=0 NRS=0 M=1 R=1.5 SA=250004 SB=250002
+ A=0.375 P=2.5 MULT=1
MM1010 N_Y_M1010_d N_A_M1010_g N_VGND_M1008_s N_VNB_M1000_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.1575 PD=1.03 PS=1.17 NRD=0 NRS=21.2724 M=1 R=1.5 SA=250005
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1013 N_Y_M1010_d N_A_M1013_g N_VGND_M1013_s N_VNB_M1000_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.20625 PD=1.03 PS=2.05 NRD=0 NRS=1.5162 M=1 R=1.5 SA=250006
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g N_VPWR_M1003_s N_VPB_M1003_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 M=1 R=3 SA=250000 SB=250005
+ A=0.75 P=4 MULT=1
MM1004 N_Y_M1003_d N_A_M1004_g N_VPWR_M1004_s N_VPB_M1003_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001 SB=250005 A=0.75
+ P=4 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_VPWR_M1004_s N_VPB_M1003_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002 SB=250004 A=0.75
+ P=4 MULT=1
MM1009 N_Y_M1007_d N_A_M1009_g N_VPWR_M1009_s N_VPB_M1003_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002 SB=250003 A=0.75
+ P=4 MULT=1
MM1011 N_Y_M1011_d N_A_M1011_g N_VPWR_M1009_s N_VPB_M1003_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250003 SB=250002 A=0.75
+ P=4 MULT=1
MM1012 N_Y_M1011_d N_A_M1012_g N_VPWR_M1012_s N_VPB_M1003_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250004 SB=250002 A=0.75
+ P=4 MULT=1
MM1014 N_Y_M1014_d N_A_M1014_g N_VPWR_M1012_s N_VPB_M1003_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250005 SB=250001 A=0.75
+ P=4 MULT=1
MM1015 N_Y_M1014_d N_A_M1015_g N_VPWR_M1015_s N_VPB_M1003_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 M=1 R=3 SA=250005 SB=250000
+ A=0.75 P=4 MULT=1
DX16_noxref N_VNB_M1000_b N_VPB_M1003_b NWDIODE A=20.436 P=20.92
*
.include "sky130_fd_sc_hvl__inv_8.pxi.spice"
*
.ends
*
*
