* File: sky130_fd_sc_hvl__a22o_1.pxi.spice
* Created: Fri Aug 28 09:32:22 2020
* 
x_PM_SKY130_FD_SC_HVL__A22O_1%VNB N_VNB_M1008_b VNB N_VNB_c_4_p VNB
+ PM_SKY130_FD_SC_HVL__A22O_1%VNB
x_PM_SKY130_FD_SC_HVL__A22O_1%VPB N_VPB_M1009_b VPB N_VPB_c_34_p VPB
+ PM_SKY130_FD_SC_HVL__A22O_1%VPB
x_PM_SKY130_FD_SC_HVL__A22O_1%A_83_81# N_A_83_81#_M1001_d N_A_83_81#_M1000_d
+ N_A_83_81#_M1008_g N_A_83_81#_M1009_g N_A_83_81#_c_76_n N_A_83_81#_c_91_p
+ N_A_83_81#_c_77_n N_A_83_81#_c_78_n N_A_83_81#_c_80_n N_A_83_81#_c_82_n
+ N_A_83_81#_c_115_p N_A_83_81#_c_83_n N_A_83_81#_c_84_n N_A_83_81#_c_85_n
+ N_A_83_81#_c_88_n PM_SKY130_FD_SC_HVL__A22O_1%A_83_81#
x_PM_SKY130_FD_SC_HVL__A22O_1%B2 N_B2_M1000_g N_B2_M1002_g B2 B2 B2 B2
+ N_B2_c_143_n N_B2_c_148_n PM_SKY130_FD_SC_HVL__A22O_1%B2
x_PM_SKY130_FD_SC_HVL__A22O_1%B1 B1 B1 B1 N_B1_M1001_g N_B1_M1004_g
+ PM_SKY130_FD_SC_HVL__A22O_1%B1
x_PM_SKY130_FD_SC_HVL__A22O_1%A1 N_A1_M1003_g N_A1_M1006_g A1 A1 A1 N_A1_c_207_n
+ PM_SKY130_FD_SC_HVL__A22O_1%A1
x_PM_SKY130_FD_SC_HVL__A22O_1%A2 N_A2_M1007_g N_A2_M1005_g A2 N_A2_c_239_n
+ PM_SKY130_FD_SC_HVL__A22O_1%A2
x_PM_SKY130_FD_SC_HVL__A22O_1%X N_X_M1008_s N_X_M1009_s X X X X X X X
+ N_X_c_259_n PM_SKY130_FD_SC_HVL__A22O_1%X
x_PM_SKY130_FD_SC_HVL__A22O_1%VPWR N_VPWR_M1009_d N_VPWR_M1003_d VPWR
+ N_VPWR_c_273_n N_VPWR_c_276_n N_VPWR_c_279_n PM_SKY130_FD_SC_HVL__A22O_1%VPWR
x_PM_SKY130_FD_SC_HVL__A22O_1%A_316_443# N_A_316_443#_M1000_s
+ N_A_316_443#_M1004_d N_A_316_443#_M1005_d N_A_316_443#_c_312_n
+ N_A_316_443#_c_313_n N_A_316_443#_c_316_n N_A_316_443#_c_319_n
+ N_A_316_443#_c_320_n N_A_316_443#_c_321_n N_A_316_443#_c_322_n
+ PM_SKY130_FD_SC_HVL__A22O_1%A_316_443#
x_PM_SKY130_FD_SC_HVL__A22O_1%VGND N_VGND_M1008_d N_VGND_M1007_d VGND
+ N_VGND_c_362_n N_VGND_c_364_n N_VGND_c_366_n PM_SKY130_FD_SC_HVL__A22O_1%VGND
cc_1 N_VNB_M1008_b N_A_83_81#_c_76_n 0.0364454f $X=-0.33 $Y=-0.265 $X2=2.5
+ $Y2=1.51
cc_2 N_VNB_M1008_b N_A_83_81#_c_77_n 0.001277f $X=-0.33 $Y=-0.265 $X2=2.77
+ $Y2=1.425
cc_3 N_VNB_M1008_b N_A_83_81#_c_78_n 0.0243114f $X=-0.33 $Y=-0.265 $X2=3.385
+ $Y2=0.545
cc_4 N_VNB_c_4_p N_A_83_81#_c_78_n 0.00265143f $X=0.24 $Y=0 $X2=3.385 $Y2=0.545
cc_5 N_VNB_M1008_b N_A_83_81#_c_80_n 0.00644733f $X=-0.33 $Y=-0.265 $X2=2.855
+ $Y2=0.545
cc_6 N_VNB_c_4_p N_A_83_81#_c_80_n 5.23982e-19 $X=0.24 $Y=0 $X2=2.855 $Y2=0.545
cc_7 N_VNB_M1008_b N_A_83_81#_c_82_n 0.00303989f $X=-0.33 $Y=-0.265 $X2=3.47
+ $Y2=0.66
cc_8 N_VNB_M1008_b N_A_83_81#_c_83_n 0.0613666f $X=-0.33 $Y=-0.265 $X2=0.75
+ $Y2=1.59
cc_9 N_VNB_M1008_b N_A_83_81#_c_84_n 0.00366547f $X=-0.33 $Y=-0.265 $X2=2.677
+ $Y2=1.51
cc_10 N_VNB_M1008_b N_A_83_81#_c_85_n 0.0491296f $X=-0.33 $Y=-0.265 $X2=0.675
+ $Y2=1.395
cc_11 N_VNB_c_4_p N_A_83_81#_c_85_n 6.33027e-19 $X=0.24 $Y=0 $X2=0.675 $Y2=1.395
cc_12 N_VNB_M1008_b N_B2_M1002_g 0.0525062f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=1.395
cc_13 N_VNB_c_4_p N_B2_M1002_g 0.00156395f $X=0.24 $Y=0 $X2=0.665 $Y2=1.395
cc_14 N_VNB_M1008_b N_B2_c_143_n 0.0605127f $X=-0.33 $Y=-0.265 $X2=2.665
+ $Y2=3.37
cc_15 N_VNB_M1008_b N_B1_M1001_g 0.0843442f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=0.91
cc_16 N_VNB_c_4_p N_B1_M1001_g 0.0023273f $X=0.24 $Y=0 $X2=0.665 $Y2=0.91
cc_17 N_VNB_M1008_b N_A1_M1006_g 0.0425572f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=1.395
cc_18 N_VNB_c_4_p N_A1_M1006_g 9.54195e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=1.395
cc_19 N_VNB_M1008_b A1 0.00761266f $X=-0.33 $Y=-0.265 $X2=0.685 $Y2=2.965
cc_20 N_VNB_M1008_b N_A1_c_207_n 0.040872f $X=-0.33 $Y=-0.265 $X2=2.665 $Y2=2.34
cc_21 N_VNB_M1008_b N_A2_M1007_g 0.0432009f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_22 N_VNB_M1008_b N_A2_c_239_n 0.0853623f $X=-0.33 $Y=-0.265 $X2=2.665
+ $Y2=1.595
cc_23 N_VNB_M1008_b N_X_c_259_n 0.069541f $X=-0.33 $Y=-0.265 $X2=2.77 $Y2=1.425
cc_24 N_VNB_c_4_p N_X_c_259_n 6.39784e-19 $X=0.24 $Y=0 $X2=2.77 $Y2=1.425
cc_25 N_VNB_M1008_b N_VGND_c_362_n 0.089026f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.105
cc_26 N_VNB_c_4_p N_VGND_c_362_n 0.00484742f $X=0.24 $Y=0 $X2=0.685 $Y2=2.105
cc_27 N_VNB_M1008_b N_VGND_c_364_n 0.101071f $X=-0.33 $Y=-0.265 $X2=3.51
+ $Y2=0.66
cc_28 N_VNB_c_4_p N_VGND_c_364_n 0.00371223f $X=0.24 $Y=0 $X2=3.51 $Y2=0.66
cc_29 N_VNB_M1008_b N_VGND_c_366_n 0.0884645f $X=-0.33 $Y=-0.265 $X2=3.47
+ $Y2=0.66
cc_30 N_VNB_c_4_p N_VGND_c_366_n 0.564589f $X=0.24 $Y=0 $X2=3.47 $Y2=0.66
cc_31 N_VPB_M1009_b N_A_83_81#_c_83_n 0.030304f $X=-0.33 $Y=1.885 $X2=0.75
+ $Y2=1.59
cc_32 N_VPB_M1009_b N_A_83_81#_c_88_n 0.0426348f $X=-0.33 $Y=1.885 $X2=0.675
+ $Y2=2.105
cc_33 VPB N_A_83_81#_c_88_n 0.00970178f $X=0 $Y=3.955 $X2=0.675 $Y2=2.105
cc_34 N_VPB_c_34_p N_A_83_81#_c_88_n 0.0152133f $X=5.04 $Y=4.07 $X2=0.675
+ $Y2=2.105
cc_35 N_VPB_M1009_b N_B2_M1000_g 0.0382985f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_36 VPB N_B2_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_37 N_VPB_c_34_p N_B2_M1000_g 0.0134686f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_38 N_VPB_M1009_b N_B2_c_143_n 0.0303133f $X=-0.33 $Y=1.885 $X2=2.665 $Y2=3.37
cc_39 N_VPB_M1009_b N_B2_c_148_n 0.00372366f $X=-0.33 $Y=1.885 $X2=2.665
+ $Y2=3.37
cc_40 N_VPB_M1009_b N_B1_M1001_g 0.0494779f $X=-0.33 $Y=1.885 $X2=0.665 $Y2=0.91
cc_41 VPB N_B1_M1001_g 0.00970178f $X=0 $Y=3.955 $X2=0.665 $Y2=0.91
cc_42 N_VPB_c_34_p N_B1_M1001_g 0.0134683f $X=5.04 $Y=4.07 $X2=0.665 $Y2=0.91
cc_43 N_VPB_M1009_b N_A1_M1003_g 0.0353896f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_44 VPB N_A1_M1003_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_45 N_VPB_c_34_p N_A1_M1003_g 0.0152133f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_46 N_VPB_M1009_b N_A1_c_207_n 0.0171659f $X=-0.33 $Y=1.885 $X2=2.665 $Y2=2.34
cc_47 N_VPB_M1009_b N_A2_M1005_g 0.0394876f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=1.395
cc_48 VPB N_A2_M1005_g 0.00970178f $X=0 $Y=3.955 $X2=0.665 $Y2=1.395
cc_49 N_VPB_c_34_p N_A2_M1005_g 0.015886f $X=5.04 $Y=4.07 $X2=0.665 $Y2=1.395
cc_50 N_VPB_M1009_b N_A2_c_239_n 0.0418169f $X=-0.33 $Y=1.885 $X2=2.665
+ $Y2=1.595
cc_51 N_VPB_M1009_b N_X_c_259_n 0.0713924f $X=-0.33 $Y=1.885 $X2=2.77 $Y2=1.425
cc_52 VPB N_X_c_259_n 8.36738e-19 $X=0 $Y=3.955 $X2=2.77 $Y2=1.425
cc_53 N_VPB_c_34_p N_X_c_259_n 0.014426f $X=5.04 $Y=4.07 $X2=2.77 $Y2=1.425
cc_54 N_VPB_M1009_b N_VPWR_c_273_n 0.0359502f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.105
cc_55 VPB N_VPWR_c_273_n 0.0034009f $X=0 $Y=3.955 $X2=0.685 $Y2=2.105
cc_56 N_VPB_c_34_p N_VPWR_c_273_n 0.0459724f $X=5.04 $Y=4.07 $X2=0.685 $Y2=2.105
cc_57 N_VPB_M1009_b N_VPWR_c_276_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_276_n 0.00406397f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_59 N_VPB_c_34_p N_VPWR_c_276_n 0.047451f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_60 N_VPB_M1009_b N_VPWR_c_279_n 0.0529852f $X=-0.33 $Y=1.885 $X2=3.47
+ $Y2=0.66
cc_61 VPB N_VPWR_c_279_n 0.56003f $X=0 $Y=3.955 $X2=3.47 $Y2=0.66
cc_62 N_VPB_c_34_p N_VPWR_c_279_n 0.0216031f $X=5.04 $Y=4.07 $X2=3.47 $Y2=0.66
cc_63 N_VPB_M1009_b N_A_316_443#_c_312_n 0.00357702f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.965
cc_64 N_VPB_M1009_b N_A_316_443#_c_313_n 0.00363242f $X=-0.33 $Y=1.885 $X2=2.665
+ $Y2=2.34
cc_65 VPB N_A_316_443#_c_313_n 0.00679947f $X=0 $Y=3.955 $X2=2.665 $Y2=2.34
cc_66 N_VPB_c_34_p N_A_316_443#_c_313_n 0.110631f $X=5.04 $Y=4.07 $X2=2.665
+ $Y2=2.34
cc_67 N_VPB_M1009_b N_A_316_443#_c_316_n 0.00196203f $X=-0.33 $Y=1.885 $X2=2.665
+ $Y2=2.34
cc_68 VPB N_A_316_443#_c_316_n 5.70856e-19 $X=0 $Y=3.955 $X2=2.665 $Y2=2.34
cc_69 N_VPB_c_34_p N_A_316_443#_c_316_n 0.0114989f $X=5.04 $Y=4.07 $X2=2.665
+ $Y2=2.34
cc_70 N_VPB_M1009_b N_A_316_443#_c_319_n 0.00107607f $X=-0.33 $Y=1.885 $X2=2.77
+ $Y2=0.63
cc_71 N_VPB_M1009_b N_A_316_443#_c_320_n 0.0075558f $X=-0.33 $Y=1.885 $X2=2.855
+ $Y2=0.545
cc_72 N_VPB_M1009_b N_A_316_443#_c_321_n 0.00535704f $X=-0.33 $Y=1.885 $X2=3.51
+ $Y2=0.63
cc_73 N_VPB_M1009_b N_A_316_443#_c_322_n 0.0574612f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_74 VPB N_A_316_443#_c_322_n 0.00101808f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_75 N_VPB_c_34_p N_A_316_443#_c_322_n 0.0158392f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_76 N_A_83_81#_c_91_p N_B2_M1000_g 0.0302314f $X=2.665 $Y=2.34 $X2=0 $Y2=0
cc_77 N_A_83_81#_c_77_n N_B2_M1002_g 0.0100937f $X=2.77 $Y=1.425 $X2=0 $Y2=0
cc_78 N_A_83_81#_c_80_n N_B2_M1002_g 0.00149484f $X=2.855 $Y=0.545 $X2=0 $Y2=0
cc_79 N_A_83_81#_c_76_n N_B2_c_143_n 0.0396107f $X=2.5 $Y=1.51 $X2=0 $Y2=0
cc_80 N_A_83_81#_c_91_p N_B2_c_143_n 0.0231573f $X=2.665 $Y=2.34 $X2=0 $Y2=0
cc_81 N_A_83_81#_c_84_n N_B2_c_143_n 0.00800965f $X=2.677 $Y=1.51 $X2=0 $Y2=0
cc_82 N_A_83_81#_c_76_n N_B2_c_148_n 0.0238596f $X=2.5 $Y=1.51 $X2=0 $Y2=0
cc_83 N_A_83_81#_c_91_p N_B2_c_148_n 0.106377f $X=2.665 $Y=2.34 $X2=0 $Y2=0
cc_84 N_A_83_81#_c_91_p B1 0.00949673f $X=2.665 $Y=2.34 $X2=0 $Y2=0
cc_85 N_A_83_81#_c_77_n B1 0.039785f $X=2.77 $Y=1.425 $X2=0 $Y2=0
cc_86 N_A_83_81#_c_78_n B1 0.0108682f $X=3.385 $Y=0.545 $X2=0 $Y2=0
cc_87 N_A_83_81#_c_82_n B1 0.0357184f $X=3.47 $Y=0.66 $X2=0 $Y2=0
cc_88 N_A_83_81#_c_84_n B1 0.0123662f $X=2.677 $Y=1.51 $X2=0 $Y2=0
cc_89 N_A_83_81#_c_91_p N_B1_M1001_g 0.0573559f $X=2.665 $Y=2.34 $X2=0 $Y2=0
cc_90 N_A_83_81#_c_77_n N_B1_M1001_g 0.0202465f $X=2.77 $Y=1.425 $X2=0 $Y2=0
cc_91 N_A_83_81#_c_78_n N_B1_M1001_g 0.0255444f $X=3.385 $Y=0.545 $X2=0 $Y2=0
cc_92 N_A_83_81#_c_80_n N_B1_M1001_g 0.00193858f $X=2.855 $Y=0.545 $X2=0 $Y2=0
cc_93 N_A_83_81#_c_82_n N_B1_M1001_g 0.00379079f $X=3.47 $Y=0.66 $X2=0 $Y2=0
cc_94 N_A_83_81#_c_84_n N_B1_M1001_g 0.00618831f $X=2.677 $Y=1.51 $X2=0 $Y2=0
cc_95 N_A_83_81#_c_78_n N_A1_M1006_g 0.00286216f $X=3.385 $Y=0.545 $X2=0 $Y2=0
cc_96 N_A_83_81#_c_82_n N_A1_M1006_g 0.0129778f $X=3.47 $Y=0.66 $X2=0 $Y2=0
cc_97 N_A_83_81#_c_82_n A1 0.0120877f $X=3.47 $Y=0.66 $X2=0.24 $Y2=0
cc_98 N_A_83_81#_c_82_n N_A1_c_207_n 7.54316e-19 $X=3.47 $Y=0.66 $X2=5.04 $Y2=0
cc_99 N_A_83_81#_c_82_n N_A2_M1007_g 2.27184e-19 $X=3.47 $Y=0.66 $X2=0 $Y2=0
cc_100 N_A_83_81#_c_115_p N_X_c_259_n 0.0223678f $X=0.75 $Y=1.51 $X2=0 $Y2=0
cc_101 N_A_83_81#_c_85_n N_X_c_259_n 0.0363348f $X=0.675 $Y=1.395 $X2=0 $Y2=0
cc_102 N_A_83_81#_c_88_n N_X_c_259_n 0.00765444f $X=0.675 $Y=2.105 $X2=0 $Y2=0
cc_103 N_A_83_81#_c_76_n N_VPWR_c_273_n 0.0193717f $X=2.5 $Y=1.51 $X2=0.24 $Y2=0
cc_104 N_A_83_81#_c_115_p N_VPWR_c_273_n 0.0126106f $X=0.75 $Y=1.51 $X2=0.24
+ $Y2=0
cc_105 N_A_83_81#_c_88_n N_VPWR_c_273_n 0.0831075f $X=0.675 $Y=2.105 $X2=0.24
+ $Y2=0
cc_106 N_A_83_81#_c_91_p N_VPWR_c_279_n 0.0230273f $X=2.665 $Y=2.34 $X2=0 $Y2=0
cc_107 N_A_83_81#_c_88_n N_VPWR_c_279_n 0.00915578f $X=0.675 $Y=2.105 $X2=0
+ $Y2=0
cc_108 N_A_83_81#_c_76_n N_A_316_443#_c_312_n 0.00603379f $X=2.5 $Y=1.51 $X2=0
+ $Y2=0
cc_109 N_A_83_81#_M1000_d N_A_316_443#_c_313_n 8.28689e-19 $X=2.525 $Y=2.215
+ $X2=5.04 $Y2=0
cc_110 N_A_83_81#_c_91_p N_A_316_443#_c_313_n 0.0178796f $X=2.665 $Y=2.34
+ $X2=5.04 $Y2=0
cc_111 N_A_83_81#_c_91_p N_A_316_443#_c_319_n 0.0450846f $X=2.665 $Y=2.34
+ $X2=2.64 $Y2=0
cc_112 N_A_83_81#_c_91_p N_A_316_443#_c_321_n 0.00614933f $X=2.665 $Y=2.34
+ $X2=2.64 $Y2=0.058
cc_113 N_A_83_81#_c_82_n N_A_316_443#_c_321_n 0.003814f $X=3.47 $Y=0.66 $X2=2.64
+ $Y2=0.058
cc_114 N_A_83_81#_c_76_n N_VGND_c_362_n 0.100023f $X=2.5 $Y=1.51 $X2=0.24 $Y2=0
cc_115 N_A_83_81#_c_77_n N_VGND_c_362_n 0.0236221f $X=2.77 $Y=1.425 $X2=0.24
+ $Y2=0
cc_116 N_A_83_81#_c_80_n N_VGND_c_362_n 0.00416061f $X=2.855 $Y=0.545 $X2=0.24
+ $Y2=0
cc_117 N_A_83_81#_c_115_p N_VGND_c_362_n 0.0251261f $X=0.75 $Y=1.51 $X2=0.24
+ $Y2=0
cc_118 N_A_83_81#_c_85_n N_VGND_c_362_n 0.054588f $X=0.675 $Y=1.395 $X2=0.24
+ $Y2=0
cc_119 N_A_83_81#_c_78_n N_VGND_c_364_n 0.010695f $X=3.385 $Y=0.545 $X2=0 $Y2=0
cc_120 N_A_83_81#_c_82_n N_VGND_c_364_n 0.0518267f $X=3.47 $Y=0.66 $X2=0 $Y2=0
cc_121 N_A_83_81#_c_78_n N_VGND_c_366_n 0.0590272f $X=3.385 $Y=0.545 $X2=0 $Y2=0
cc_122 N_A_83_81#_c_80_n N_VGND_c_366_n 0.0185205f $X=2.855 $Y=0.545 $X2=0 $Y2=0
cc_123 N_A_83_81#_c_85_n N_VGND_c_366_n 0.00925078f $X=0.675 $Y=1.395 $X2=0
+ $Y2=0
cc_124 N_A_83_81#_c_77_n A_519_107# 0.00778705f $X=2.77 $Y=1.425 $X2=0 $Y2=0
cc_125 N_A_83_81#_c_80_n A_519_107# 9.83485e-19 $X=2.855 $Y=0.545 $X2=0 $Y2=0
cc_126 N_B2_M1000_g N_B1_M1001_g 0.0196699f $X=2.275 $Y=2.965 $X2=0 $Y2=0
cc_127 N_B2_M1002_g N_B1_M1001_g 0.109469f $X=2.345 $Y=0.91 $X2=0 $Y2=0
cc_128 N_B2_c_148_n N_B1_M1001_g 4.91873e-19 $X=2.155 $Y=1.89 $X2=0 $Y2=0
cc_129 N_B2_M1000_g N_VPWR_c_273_n 7.85783e-19 $X=2.275 $Y=2.965 $X2=0.24 $Y2=0
cc_130 N_B2_M1000_g N_VPWR_c_279_n 0.0176477f $X=2.275 $Y=2.965 $X2=0 $Y2=0
cc_131 N_B2_c_148_n N_VPWR_c_279_n 0.00973411f $X=2.155 $Y=1.89 $X2=0 $Y2=0
cc_132 N_B2_M1000_g N_A_316_443#_c_312_n 0.01893f $X=2.275 $Y=2.965 $X2=0 $Y2=0
cc_133 N_B2_c_148_n N_A_316_443#_c_312_n 0.0393764f $X=2.155 $Y=1.89 $X2=0 $Y2=0
cc_134 N_B2_M1000_g N_A_316_443#_c_313_n 0.0234252f $X=2.275 $Y=2.965 $X2=5.04
+ $Y2=0
cc_135 N_B2_c_148_n N_A_316_443#_c_313_n 0.00746783f $X=2.155 $Y=1.89 $X2=5.04
+ $Y2=0
cc_136 N_B2_M1002_g N_VGND_c_362_n 0.0382459f $X=2.345 $Y=0.91 $X2=0.24 $Y2=0
cc_137 N_B2_c_143_n N_VGND_c_362_n 0.0032209f $X=2.155 $Y=1.89 $X2=0.24 $Y2=0
cc_138 N_B2_M1002_g N_VGND_c_366_n 0.021986f $X=2.345 $Y=0.91 $X2=0 $Y2=0
cc_139 B1 N_A1_M1006_g 7.49795e-19 $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_140 N_B1_M1001_g N_A1_M1006_g 0.0160006f $X=3.055 $Y=0.91 $X2=0 $Y2=0
cc_141 B1 A1 0.0135342f $X=3.035 $Y=0.84 $X2=0.24 $Y2=0
cc_142 N_B1_M1001_g A1 0.00219365f $X=3.055 $Y=0.91 $X2=0.24 $Y2=0
cc_143 B1 N_A1_c_207_n 7.70211e-19 $X=3.035 $Y=0.84 $X2=5.04 $Y2=0
cc_144 N_B1_M1001_g N_A1_c_207_n 0.0499049f $X=3.055 $Y=0.91 $X2=5.04 $Y2=0
cc_145 N_B1_M1001_g N_VPWR_c_276_n 6.22341e-19 $X=3.055 $Y=0.91 $X2=0 $Y2=0
cc_146 N_B1_M1001_g N_VPWR_c_279_n 0.0231149f $X=3.055 $Y=0.91 $X2=0 $Y2=0
cc_147 N_B1_M1001_g N_A_316_443#_c_313_n 0.022703f $X=3.055 $Y=0.91 $X2=5.04
+ $Y2=0
cc_148 N_B1_M1001_g N_A_316_443#_c_319_n 0.041302f $X=3.055 $Y=0.91 $X2=2.64
+ $Y2=0
cc_149 N_B1_M1001_g N_A_316_443#_c_321_n 0.00776846f $X=3.055 $Y=0.91 $X2=2.64
+ $Y2=0.058
cc_150 N_B1_M1001_g N_VGND_c_362_n 9.95e-19 $X=3.055 $Y=0.91 $X2=0.24 $Y2=0
cc_151 N_B1_M1001_g N_VGND_c_364_n 5.07725e-19 $X=3.055 $Y=0.91 $X2=0 $Y2=0
cc_152 B1 N_VGND_c_366_n 0.00130112f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_153 N_B1_M1001_g N_VGND_c_366_n 0.00594788f $X=3.055 $Y=0.91 $X2=0 $Y2=0
cc_154 N_A1_M1006_g N_A2_M1007_g 0.0576129f $X=3.86 $Y=0.91 $X2=0 $Y2=0
cc_155 N_A1_M1003_g N_A2_M1005_g 0.0169537f $X=3.835 $Y=2.965 $X2=0 $Y2=0
cc_156 A1 A2 0.0186148f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_157 A1 N_A2_c_239_n 0.0225955f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A1_c_207_n N_A2_c_239_n 0.0576129f $X=3.77 $Y=1.63 $X2=0 $Y2=0
cc_159 N_A1_M1003_g N_VPWR_c_276_n 0.0712157f $X=3.835 $Y=2.965 $X2=0 $Y2=0
cc_160 N_A1_M1003_g N_VPWR_c_279_n 0.00783253f $X=3.835 $Y=2.965 $X2=0 $Y2=0
cc_161 N_A1_M1003_g N_A_316_443#_c_313_n 0.00161577f $X=3.835 $Y=2.965 $X2=5.04
+ $Y2=0
cc_162 N_A1_M1003_g N_A_316_443#_c_319_n 0.00375436f $X=3.835 $Y=2.965 $X2=2.64
+ $Y2=0
cc_163 N_A1_M1003_g N_A_316_443#_c_320_n 0.0117512f $X=3.835 $Y=2.965 $X2=2.64
+ $Y2=0.058
cc_164 A1 N_A_316_443#_c_320_n 0.0762994f $X=4.475 $Y=1.58 $X2=2.64 $Y2=0.058
cc_165 N_A1_c_207_n N_A_316_443#_c_320_n 0.0186055f $X=3.77 $Y=1.63 $X2=2.64
+ $Y2=0.058
cc_166 A1 N_A_316_443#_c_321_n 0.00374296f $X=4.475 $Y=1.58 $X2=2.64 $Y2=0.058
cc_167 N_A1_M1006_g N_VGND_c_364_n 0.0549867f $X=3.86 $Y=0.91 $X2=0 $Y2=0
cc_168 A1 N_VGND_c_364_n 0.063458f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A1_M1006_g N_VGND_c_366_n 0.0106394f $X=3.86 $Y=0.91 $X2=0 $Y2=0
cc_170 N_A2_M1005_g N_VPWR_c_276_n 0.0676936f $X=4.615 $Y=2.965 $X2=0 $Y2=0
cc_171 N_A2_M1005_g N_VPWR_c_279_n 0.0108276f $X=4.615 $Y=2.965 $X2=0 $Y2=0
cc_172 N_A2_M1005_g N_A_316_443#_c_320_n 0.0131445f $X=4.615 $Y=2.965 $X2=2.64
+ $Y2=0.058
cc_173 A2 N_A_316_443#_c_320_n 0.0244725f $X=4.955 $Y=1.58 $X2=2.64 $Y2=0.058
cc_174 N_A2_c_239_n N_A_316_443#_c_320_n 0.0438482f $X=4.99 $Y=1.63 $X2=2.64
+ $Y2=0.058
cc_175 N_A2_M1005_g N_A_316_443#_c_322_n 0.0344025f $X=4.615 $Y=2.965 $X2=0
+ $Y2=0
cc_176 N_A2_M1007_g N_VGND_c_364_n 0.0745487f $X=4.57 $Y=0.91 $X2=0 $Y2=0
cc_177 A2 N_VGND_c_364_n 0.0236502f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A2_c_239_n N_VGND_c_364_n 0.00912004f $X=4.99 $Y=1.63 $X2=0 $Y2=0
cc_179 N_X_c_259_n N_VPWR_c_273_n 0.0678262f $X=0.275 $Y=0.68 $X2=0.24 $Y2=0
cc_180 N_X_M1009_s N_VPWR_c_279_n 0.00221032f $X=0.15 $Y=2.215 $X2=0 $Y2=0
cc_181 N_X_c_259_n N_VPWR_c_279_n 0.0375086f $X=0.275 $Y=0.68 $X2=0 $Y2=0
cc_182 N_X_c_259_n N_VGND_c_362_n 0.0332864f $X=0.275 $Y=0.68 $X2=0.24 $Y2=0
cc_183 N_X_M1008_s N_VGND_c_366_n 0.00137624f $X=0.15 $Y=0.535 $X2=0 $Y2=0
cc_184 N_X_c_259_n N_VGND_c_366_n 0.0283435f $X=0.275 $Y=0.68 $X2=0 $Y2=0
cc_185 N_VPWR_c_279_n N_A_316_443#_M1000_s 0.0104329f $X=4.545 $Y=3.59 $X2=0
+ $Y2=3.985
cc_186 N_VPWR_c_279_n N_A_316_443#_M1004_d 0.00221032f $X=4.545 $Y=3.59 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_273_n N_A_316_443#_c_312_n 0.113676f $X=1.075 $Y=2.34 $X2=0.24
+ $Y2=4.07
cc_188 N_VPWR_c_279_n N_A_316_443#_c_312_n 0.0209992f $X=4.545 $Y=3.59 $X2=0.24
+ $Y2=4.07
cc_189 N_VPWR_c_276_n N_A_316_443#_c_313_n 0.00650116f $X=4.225 $Y=2.365
+ $X2=5.04 $Y2=4.07
cc_190 N_VPWR_c_279_n N_A_316_443#_c_313_n 0.0617374f $X=4.545 $Y=3.59 $X2=5.04
+ $Y2=4.07
cc_191 N_VPWR_c_273_n N_A_316_443#_c_316_n 0.00827679f $X=1.075 $Y=2.34 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_279_n N_A_316_443#_c_316_n 0.00651138f $X=4.545 $Y=3.59 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_276_n N_A_316_443#_c_319_n 0.0556936f $X=4.225 $Y=2.365 $X2=2.64
+ $Y2=4.013
cc_194 N_VPWR_c_279_n N_A_316_443#_c_319_n 0.0265939f $X=4.545 $Y=3.59 $X2=2.64
+ $Y2=4.013
cc_195 N_VPWR_c_276_n N_A_316_443#_c_320_n 0.0658158f $X=4.225 $Y=2.365 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_276_n N_A_316_443#_c_322_n 0.10622f $X=4.225 $Y=2.365 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_279_n N_A_316_443#_c_322_n 0.0417129f $X=4.545 $Y=3.59 $X2=0
+ $Y2=0
cc_198 N_A_316_443#_c_320_n N_VGND_c_364_n 0.00479357f $X=4.84 $Y=2.015 $X2=0
+ $Y2=0
cc_199 N_VGND_c_366_n A_519_107# 0.00375338f $X=5.01 $Y=0.48 $X2=0 $Y2=0
