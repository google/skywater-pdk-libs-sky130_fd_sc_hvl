* File: sky130_fd_sc_hvl__nand3_1.pex.spice
* Created: Fri Aug 28 09:38:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__NAND3_1%VNB 5 7 11 25
r17 7 25 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0.058
r18 7 11 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0
r19 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r20 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND3_1%VPB 4 6 14 21
r30 10 21 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=4.07
+ $X2=1.68 $Y2=4.013
r31 10 14 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=4.07
+ $X2=3.12 $Y2=4.07
r32 9 14 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=3.12 $Y2=4.07
r33 9 10 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r34 6 21 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=4.012
+ $X2=1.68 $Y2=4.013
r35 4 14 52 $w=1.7e-07 $l=3.16221e-06 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=3.12 $Y2=4.07
r36 4 9 52 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND3_1%C 3 7 9 10 14 15
r21 14 17 39.8984 $w=5.7e-07 $l=4.15e-07 $layer=POLY_cond $X=0.93 $Y=1.67
+ $X2=0.93 $Y2=2.085
r22 14 16 24.8801 $w=5.7e-07 $l=2.55e-07 $layer=POLY_cond $X=0.93 $Y=1.67
+ $X2=0.93 $Y2=1.415
r23 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.83
+ $Y=1.67 $X2=0.83 $Y2=1.67
r24 10 15 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.67
+ $X2=0.83 $Y2=1.67
r25 9 10 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.67 $X2=0.72
+ $Y2=1.67
r26 7 16 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.965 $Y=0.91 $X2=0.965
+ $Y2=1.415
r27 3 17 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.895 $Y=2.965
+ $X2=0.895 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND3_1%B 3 6 8 9 13 15
r31 13 16 28.8219 $w=7.1e-07 $l=3.35e-07 $layer=POLY_cond $X=1.78 $Y=1.56
+ $X2=1.78 $Y2=1.895
r32 13 15 16.5107 $w=7.1e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.56
+ $X2=1.78 $Y2=1.395
r33 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.97
+ $Y=1.56 $X2=1.97 $Y2=1.56
r34 9 14 7.8307 $w=3.88e-07 $l=2.65e-07 $layer=LI1_cond $X=2.08 $Y=1.295
+ $X2=2.08 $Y2=1.56
r35 8 9 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.08 $Y=0.925 $X2=2.08
+ $Y2=1.295
r36 6 16 114.496 $w=5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.675 $Y=2.965
+ $X2=1.675 $Y2=1.895
r37 3 15 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.675 $Y=0.91 $X2=1.675
+ $Y2=1.395
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND3_1%A 3 6 8 9 13 15
r28 13 16 32.0682 $w=5.8e-07 $l=3.35e-07 $layer=POLY_cond $X=2.635 $Y=1.56
+ $X2=2.635 $Y2=1.895
r29 13 15 16.3863 $w=5.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.56
+ $X2=2.635 $Y2=1.395
r30 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.56 $X2=2.59 $Y2=1.56
r31 9 14 11.311 $w=2.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.59 $Y=1.295
+ $X2=2.59 $Y2=1.56
r32 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.59 $Y=0.925 $X2=2.59
+ $Y2=1.295
r33 6 16 114.496 $w=5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.675 $Y=2.965
+ $X2=2.675 $Y2=1.895
r34 3 15 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.595 $Y=0.91 $X2=2.595
+ $Y2=1.395
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND3_1%VPWR 1 2 7 10 20 27
r24 23 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.715 $Y=3.59
+ $X2=2.715 $Y2=3.59
r25 20 23 12.2 $w=1.248e-06 $l=1.25e-06 $layer=LI1_cond $X=2.175 $Y=2.34
+ $X2=2.175 $Y2=3.59
r26 14 17 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.195 $Y=3.63
+ $X2=0.915 $Y2=3.63
r27 13 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.915 $Y=3.59
+ $X2=0.915 $Y2=3.59
r28 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.195 $Y=3.59
+ $X2=0.195 $Y2=3.59
r29 10 13 16.3979 $w=9.28e-07 $l=1.25e-06 $layer=LI1_cond $X=0.555 $Y=2.34
+ $X2=0.555 $Y2=3.59
r30 7 27 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=1.635 $Y=3.63
+ $X2=2.715 $Y2=3.63
r31 7 17 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.635 $Y=3.63
+ $X2=0.915 $Y2=3.63
r32 7 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.635 $Y=3.59
+ $X2=1.635 $Y2=3.59
r33 2 23 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.925
+ $Y=2.215 $X2=2.065 $Y2=3.59
r34 2 20 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.925
+ $Y=2.215 $X2=2.065 $Y2=2.34
r35 1 13 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.36
+ $Y=2.215 $X2=0.505 $Y2=3.59
r36 1 10 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.36
+ $Y=2.215 $X2=0.505 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND3_1%Y 1 2 3 12 16 17 18 19 20 21 22 23 24 36 59
r40 59 60 1.67296 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=3.07 $Y=1.295 $X2=3.07
+ $Y2=1.325
r41 24 55 20.1113 $w=2.53e-07 $l=4.45e-07 $layer=LI1_cond $X=3.107 $Y=3.145
+ $X2=3.107 $Y2=3.59
r42 23 24 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.107 $Y=2.775
+ $X2=3.107 $Y2=3.145
r43 22 23 19.6593 $w=2.53e-07 $l=4.35e-07 $layer=LI1_cond $X=3.107 $Y=2.34
+ $X2=3.107 $Y2=2.775
r44 21 41 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.107 $Y=1.99
+ $X2=3.107 $Y2=1.905
r45 21 45 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.107 $Y=1.99
+ $X2=3.107 $Y2=2.075
r46 21 22 10.9821 $w=2.53e-07 $l=2.43e-07 $layer=LI1_cond $X=3.107 $Y=2.097
+ $X2=3.107 $Y2=2.34
r47 21 45 0.994265 $w=2.53e-07 $l=2.2e-08 $layer=LI1_cond $X=3.107 $Y=2.097
+ $X2=3.107 $Y2=2.075
r48 20 41 10.8465 $w=2.53e-07 $l=2.4e-07 $layer=LI1_cond $X=3.107 $Y=1.665
+ $X2=3.107 $Y2=1.905
r49 19 59 0.97783 $w=3.28e-07 $l=2.8e-08 $layer=LI1_cond $X=3.07 $Y=1.267
+ $X2=3.07 $Y2=1.295
r50 19 34 3.73671 $w=3.28e-07 $l=1.07e-07 $layer=LI1_cond $X=3.07 $Y=1.267
+ $X2=3.07 $Y2=1.16
r51 19 20 14.1457 $w=2.53e-07 $l=3.13e-07 $layer=LI1_cond $X=3.107 $Y=1.352
+ $X2=3.107 $Y2=1.665
r52 19 60 1.22023 $w=2.53e-07 $l=2.7e-08 $layer=LI1_cond $X=3.107 $Y=1.352
+ $X2=3.107 $Y2=1.325
r53 18 34 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=3.07 $Y=0.925
+ $X2=3.07 $Y2=1.16
r54 18 36 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.07 $Y=0.925
+ $X2=3.07 $Y2=0.66
r55 16 21 2.83584 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.98 $Y=1.99
+ $X2=3.107 $Y2=1.99
r56 16 17 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=2.98 $Y=1.99
+ $X2=1.37 $Y2=1.99
r57 12 14 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=1.285 $Y=2.34
+ $X2=1.285 $Y2=3.59
r58 10 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.285 $Y=2.075
+ $X2=1.37 $Y2=1.99
r59 10 12 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.285 $Y=2.075
+ $X2=1.285 $Y2=2.34
r60 3 55 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.925
+ $Y=2.215 $X2=3.065 $Y2=3.59
r61 3 22 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.925
+ $Y=2.215 $X2=3.065 $Y2=2.34
r62 2 14 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=2.215 $X2=1.285 $Y2=3.59
r63 2 12 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=2.215 $X2=1.285 $Y2=2.34
r64 1 36 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.845
+ $Y=0.535 $X2=2.99 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__NAND3_1%VGND 1 4 7
r19 7 13 1.35975 $w=1.613e-06 $l=1.8e-07 $layer=LI1_cond $X=0.897 $Y=0.48
+ $X2=0.897 $Y2=0.66
r20 7 8 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.18 $Y=0.48
+ $X2=0.18 $Y2=0.48
r21 4 8 0.552824 $w=3.7e-07 $l=1.44e-06 $layer=MET1_cond $X=1.62 $Y=0.44
+ $X2=0.18 $Y2=0.44
r22 4 7 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.62 $Y=0.48
+ $X2=1.62 $Y2=0.48
r23 1 13 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.43
+ $Y=0.535 $X2=0.575 $Y2=0.66
.ends

