* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 VGND a_1630_171# GCLK VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X1 a_1783_171# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 a_58_159# a_423_71# a_495_311# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 VPWR a_1261_133# a_1630_171# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X4 VPWR SCE a_219_457# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X5 VPWR CLK a_423_71# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X6 VPWR a_1630_171# GCLK VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X7 a_431_431# a_423_71# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR a_495_311# a_1261_133# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X9 VGND CLK a_423_71# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 a_1630_171# a_1261_133# a_1783_171# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 a_58_159# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X12 a_219_457# GATE a_58_159# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X13 a_495_311# a_423_71# a_1219_457# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 a_1219_457# a_1261_133# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_495_311# a_1261_133# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X16 a_58_159# a_431_431# a_495_311# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X17 a_1630_171# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X18 VGND GATE a_58_159# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X19 a_495_311# a_431_431# a_1219_159# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X20 a_431_431# a_423_71# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X21 a_1219_159# a_1261_133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends
