* File: sky130_fd_sc_hvl__inv_16.pxi.spice
* Created: Fri Aug 28 09:35:52 2020
* 
x_PM_SKY130_FD_SC_HVL__INV_16%VNB N_VNB_M1002_b VNB N_VNB_c_2_p
+ PM_SKY130_FD_SC_HVL__INV_16%VNB
x_PM_SKY130_FD_SC_HVL__INV_16%VPB N_VPB_M1000_b VPB N_VPB_c_69_p
+ PM_SKY130_FD_SC_HVL__INV_16%VPB
x_PM_SKY130_FD_SC_HVL__INV_16%A N_A_c_170_n N_A_M1002_g N_A_M1000_g N_A_c_172_n
+ N_A_M1003_g N_A_M1001_g N_A_c_174_n N_A_M1005_g N_A_M1004_g N_A_c_176_n
+ N_A_M1006_g N_A_M1008_g N_A_c_178_n N_A_M1007_g N_A_M1009_g N_A_c_180_n
+ N_A_M1012_g N_A_M1010_g N_A_c_182_n N_A_M1013_g N_A_M1011_g N_A_c_184_n
+ N_A_M1016_g N_A_M1014_g N_A_c_186_n N_A_M1018_g N_A_M1015_g N_A_c_188_n
+ N_A_M1020_g N_A_M1017_g N_A_c_190_n N_A_M1021_g N_A_M1019_g N_A_c_192_n
+ N_A_M1023_g N_A_M1022_g N_A_c_194_n N_A_M1025_g N_A_M1024_g N_A_c_196_n
+ N_A_M1028_g N_A_M1026_g N_A_c_198_n N_A_M1030_g N_A_M1027_g N_A_c_200_n
+ N_A_M1031_g N_A_M1029_g A N_A_c_202_n N_A_c_203_n N_A_c_204_n N_A_c_205_n
+ N_A_c_206_n N_A_c_207_n N_A_c_208_n N_A_c_209_n N_A_c_210_n N_A_c_275_p
+ N_A_c_362_p N_A_c_211_n N_A_c_283_p N_A_c_284_p N_A_c_372_p N_A_c_212_n
+ N_A_c_292_p N_A_c_293_p N_A_c_382_p N_A_c_213_n N_A_c_301_p A N_A_c_302_p
+ N_A_c_392_p N_A_c_214_n N_A_c_310_p N_A_c_311_p N_A_c_402_p N_A_c_215_n
+ N_A_c_319_p N_A_c_320_p N_A_c_412_p N_A_c_328_p PM_SKY130_FD_SC_HVL__INV_16%A
x_PM_SKY130_FD_SC_HVL__INV_16%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_M1008_d
+ N_VPWR_M1010_d N_VPWR_M1014_d N_VPWR_M1017_d N_VPWR_M1022_d N_VPWR_M1026_d
+ N_VPWR_M1029_d VPWR N_VPWR_c_534_n N_VPWR_c_537_n N_VPWR_c_540_n
+ N_VPWR_c_543_n N_VPWR_c_546_n N_VPWR_c_549_n N_VPWR_c_552_n N_VPWR_c_555_n
+ N_VPWR_c_558_n N_VPWR_c_561_n PM_SKY130_FD_SC_HVL__INV_16%VPWR
x_PM_SKY130_FD_SC_HVL__INV_16%Y N_Y_M1002_d N_Y_M1005_d N_Y_M1007_d N_Y_M1013_d
+ N_Y_M1018_d N_Y_M1021_d N_Y_M1025_d N_Y_M1030_d N_Y_M1000_s N_Y_M1004_s
+ N_Y_M1009_s N_Y_M1011_s N_Y_M1015_s N_Y_M1019_s N_Y_M1024_s N_Y_M1027_s Y
+ N_Y_c_693_n N_Y_c_696_n N_Y_c_699_n N_Y_c_702_n N_Y_c_705_n N_Y_c_708_n
+ N_Y_c_711_n N_Y_c_714_n N_Y_c_790_n N_Y_c_851_n N_Y_c_794_n N_Y_c_798_n
+ N_Y_c_799_n N_Y_c_803_n N_Y_c_804_n N_Y_c_808_n N_Y_c_809_n N_Y_c_813_n
+ N_Y_c_814_n N_Y_c_818_n N_Y_c_819_n N_Y_c_823_n PM_SKY130_FD_SC_HVL__INV_16%Y
x_PM_SKY130_FD_SC_HVL__INV_16%VGND N_VGND_M1002_s N_VGND_M1003_s N_VGND_M1006_s
+ N_VGND_M1012_s N_VGND_M1016_s N_VGND_M1020_s N_VGND_M1023_s N_VGND_M1028_s
+ N_VGND_M1031_s VGND N_VGND_c_895_n N_VGND_c_897_n N_VGND_c_899_n
+ N_VGND_c_901_n N_VGND_c_903_n N_VGND_c_905_n N_VGND_c_907_n N_VGND_c_909_n
+ N_VGND_c_911_n N_VGND_c_913_n PM_SKY130_FD_SC_HVL__INV_16%VGND
cc_1 N_VNB_M1002_b N_A_c_170_n 0.0467577f $X=-0.33 $Y=-0.265 $X2=0.675 $Y2=1.565
cc_2 N_VNB_c_2_p N_A_c_170_n 0.00114087f $X=0.24 $Y=0 $X2=0.675 $Y2=1.565
cc_3 N_VNB_M1002_b N_A_c_172_n 0.0394647f $X=-0.33 $Y=-0.265 $X2=1.455 $Y2=1.565
cc_4 N_VNB_c_2_p N_A_c_172_n 7.55443e-19 $X=0.24 $Y=0 $X2=1.455 $Y2=1.565
cc_5 N_VNB_M1002_b N_A_c_174_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=2.235 $Y2=1.565
cc_6 N_VNB_c_2_p N_A_c_174_n 7.55443e-19 $X=0.24 $Y=0 $X2=2.235 $Y2=1.565
cc_7 N_VNB_M1002_b N_A_c_176_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=3.015 $Y2=1.565
cc_8 N_VNB_c_2_p N_A_c_176_n 7.55443e-19 $X=0.24 $Y=0 $X2=3.015 $Y2=1.565
cc_9 N_VNB_M1002_b N_A_c_178_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=3.795 $Y2=1.565
cc_10 N_VNB_c_2_p N_A_c_178_n 7.55443e-19 $X=0.24 $Y=0 $X2=3.795 $Y2=1.565
cc_11 N_VNB_M1002_b N_A_c_180_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=4.575
+ $Y2=1.565
cc_12 N_VNB_c_2_p N_A_c_180_n 7.55443e-19 $X=0.24 $Y=0 $X2=4.575 $Y2=1.565
cc_13 N_VNB_M1002_b N_A_c_182_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=5.355
+ $Y2=1.565
cc_14 N_VNB_c_2_p N_A_c_182_n 7.55443e-19 $X=0.24 $Y=0 $X2=5.355 $Y2=1.565
cc_15 N_VNB_M1002_b N_A_c_184_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=6.135
+ $Y2=1.565
cc_16 N_VNB_c_2_p N_A_c_184_n 7.55443e-19 $X=0.24 $Y=0 $X2=6.135 $Y2=1.565
cc_17 N_VNB_M1002_b N_A_c_186_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=6.915
+ $Y2=1.565
cc_18 N_VNB_c_2_p N_A_c_186_n 7.55443e-19 $X=0.24 $Y=0 $X2=6.915 $Y2=1.565
cc_19 N_VNB_M1002_b N_A_c_188_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=7.695
+ $Y2=1.565
cc_20 N_VNB_c_2_p N_A_c_188_n 7.55443e-19 $X=0.24 $Y=0 $X2=7.695 $Y2=1.565
cc_21 N_VNB_M1002_b N_A_c_190_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=8.475
+ $Y2=1.565
cc_22 N_VNB_c_2_p N_A_c_190_n 7.55443e-19 $X=0.24 $Y=0 $X2=8.475 $Y2=1.565
cc_23 N_VNB_M1002_b N_A_c_192_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=9.255
+ $Y2=1.565
cc_24 N_VNB_c_2_p N_A_c_192_n 7.55443e-19 $X=0.24 $Y=0 $X2=9.255 $Y2=1.565
cc_25 N_VNB_M1002_b N_A_c_194_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=10.035
+ $Y2=1.565
cc_26 N_VNB_c_2_p N_A_c_194_n 7.55443e-19 $X=0.24 $Y=0 $X2=10.035 $Y2=1.565
cc_27 N_VNB_M1002_b N_A_c_196_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=10.815
+ $Y2=1.565
cc_28 N_VNB_c_2_p N_A_c_196_n 7.55443e-19 $X=0.24 $Y=0 $X2=10.815 $Y2=1.565
cc_29 N_VNB_M1002_b N_A_c_198_n 0.0394628f $X=-0.33 $Y=-0.265 $X2=11.595
+ $Y2=1.565
cc_30 N_VNB_c_2_p N_A_c_198_n 7.55443e-19 $X=0.24 $Y=0 $X2=11.595 $Y2=1.565
cc_31 N_VNB_M1002_b N_A_c_200_n 0.537945f $X=-0.33 $Y=-0.265 $X2=12.375
+ $Y2=1.565
cc_32 N_VNB_c_2_p N_A_c_200_n 7.55443e-19 $X=0.24 $Y=0 $X2=12.375 $Y2=1.565
cc_33 N_VNB_M1002_b N_A_c_202_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=2.04
+ $Y2=1.665
cc_34 N_VNB_M1002_b N_A_c_203_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=3.59
+ $Y2=1.665
cc_35 N_VNB_M1002_b N_A_c_204_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=5.15
+ $Y2=1.665
cc_36 N_VNB_M1002_b N_A_c_205_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=6.71
+ $Y2=1.665
cc_37 N_VNB_M1002_b N_A_c_206_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=8.27
+ $Y2=1.665
cc_38 N_VNB_M1002_b N_A_c_207_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=9.83
+ $Y2=1.665
cc_39 N_VNB_M1002_b N_A_c_208_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=11.39
+ $Y2=1.665
cc_40 N_VNB_M1002_b N_A_c_209_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=11.39
+ $Y2=1.665
cc_41 N_VNB_M1002_b N_A_c_210_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=2.07
+ $Y2=1.665
cc_42 N_VNB_M1002_b N_A_c_211_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=3.62
+ $Y2=1.665
cc_43 N_VNB_M1002_b N_A_c_212_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=5.18
+ $Y2=1.665
cc_44 N_VNB_M1002_b N_A_c_213_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=6.74
+ $Y2=1.665
cc_45 N_VNB_M1002_b N_A_c_214_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=8.3 $Y2=1.665
cc_46 N_VNB_M1002_b N_A_c_215_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=9.86
+ $Y2=1.665
cc_47 N_VNB_M1002_b N_VGND_c_895_n 0.0819067f $X=-0.33 $Y=-0.265 $X2=3.795
+ $Y2=1.08
cc_48 N_VNB_c_2_p N_VGND_c_895_n 0.00148993f $X=0.24 $Y=0 $X2=3.795 $Y2=1.08
cc_49 N_VNB_M1002_b N_VGND_c_897_n 0.0469183f $X=-0.33 $Y=-0.265 $X2=4.575
+ $Y2=1.08
cc_50 N_VNB_c_2_p N_VGND_c_897_n 0.00248228f $X=0.24 $Y=0 $X2=4.575 $Y2=1.08
cc_51 N_VNB_M1002_b N_VGND_c_899_n 0.0461879f $X=-0.33 $Y=-0.265 $X2=5.36
+ $Y2=2.965
cc_52 N_VNB_c_2_p N_VGND_c_899_n 0.00248228f $X=0.24 $Y=0 $X2=5.36 $Y2=2.965
cc_53 N_VNB_M1002_b N_VGND_c_901_n 0.0461879f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_54 N_VNB_c_2_p N_VGND_c_901_n 0.00248228f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_55 N_VNB_M1002_b N_VGND_c_903_n 0.0461879f $X=-0.33 $Y=-0.265 $X2=7.695
+ $Y2=1.08
cc_56 N_VNB_c_2_p N_VGND_c_903_n 0.00248228f $X=0.24 $Y=0 $X2=7.695 $Y2=1.08
cc_57 N_VNB_M1002_b N_VGND_c_905_n 0.0461879f $X=-0.33 $Y=-0.265 $X2=8.48
+ $Y2=2.005
cc_58 N_VNB_c_2_p N_VGND_c_905_n 0.00248228f $X=0.24 $Y=0 $X2=8.48 $Y2=2.005
cc_59 N_VNB_M1002_b N_VGND_c_907_n 0.0461879f $X=-0.33 $Y=-0.265 $X2=9.26
+ $Y2=2.965
cc_60 N_VNB_c_2_p N_VGND_c_907_n 0.00248228f $X=0.24 $Y=0 $X2=9.26 $Y2=2.965
cc_61 N_VNB_M1002_b N_VGND_c_909_n 0.0461879f $X=-0.33 $Y=-0.265 $X2=10.815
+ $Y2=1.565
cc_62 N_VNB_c_2_p N_VGND_c_909_n 0.00248228f $X=0.24 $Y=0 $X2=10.815 $Y2=1.565
cc_63 N_VNB_M1002_b N_VGND_c_911_n 0.0694401f $X=-0.33 $Y=-0.265 $X2=11.595
+ $Y2=1.08
cc_64 N_VNB_c_2_p N_VGND_c_911_n 0.00171356f $X=0.24 $Y=0 $X2=11.595 $Y2=1.08
cc_65 N_VNB_M1002_b N_VGND_c_913_n 0.214083f $X=-0.33 $Y=-0.265 $X2=11.6
+ $Y2=2.005
cc_66 N_VNB_c_2_p N_VGND_c_913_n 1.43756f $X=0.24 $Y=0 $X2=11.6 $Y2=2.005
cc_67 N_VPB_M1000_b N_A_M1000_g 0.0502865f $X=-0.33 $Y=1.885 $X2=0.68 $Y2=2.965
cc_68 VPB N_A_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.68 $Y2=2.965
cc_69 N_VPB_c_69_p N_A_M1000_g 0.0166568f $X=13.2 $Y=4.07 $X2=0.68 $Y2=2.965
cc_70 N_VPB_M1000_b N_A_M1001_g 0.040726f $X=-0.33 $Y=1.885 $X2=1.46 $Y2=2.965
cc_71 VPB N_A_M1001_g 0.00970178f $X=0 $Y=3.955 $X2=1.46 $Y2=2.965
cc_72 N_VPB_c_69_p N_A_M1001_g 0.0157621f $X=13.2 $Y=4.07 $X2=1.46 $Y2=2.965
cc_73 N_VPB_M1000_b N_A_M1004_g 0.040726f $X=-0.33 $Y=1.885 $X2=2.24 $Y2=2.965
cc_74 VPB N_A_M1004_g 0.00970178f $X=0 $Y=3.955 $X2=2.24 $Y2=2.965
cc_75 N_VPB_c_69_p N_A_M1004_g 0.0157621f $X=13.2 $Y=4.07 $X2=2.24 $Y2=2.965
cc_76 N_VPB_M1000_b N_A_M1008_g 0.040726f $X=-0.33 $Y=1.885 $X2=3.02 $Y2=2.965
cc_77 VPB N_A_M1008_g 0.00970178f $X=0 $Y=3.955 $X2=3.02 $Y2=2.965
cc_78 N_VPB_c_69_p N_A_M1008_g 0.0157621f $X=13.2 $Y=4.07 $X2=3.02 $Y2=2.965
cc_79 N_VPB_M1000_b N_A_M1009_g 0.040726f $X=-0.33 $Y=1.885 $X2=3.8 $Y2=2.965
cc_80 VPB N_A_M1009_g 0.00970178f $X=0 $Y=3.955 $X2=3.8 $Y2=2.965
cc_81 N_VPB_c_69_p N_A_M1009_g 0.0157621f $X=13.2 $Y=4.07 $X2=3.8 $Y2=2.965
cc_82 N_VPB_M1000_b N_A_M1010_g 0.040726f $X=-0.33 $Y=1.885 $X2=4.58 $Y2=2.965
cc_83 VPB N_A_M1010_g 0.00970178f $X=0 $Y=3.955 $X2=4.58 $Y2=2.965
cc_84 N_VPB_c_69_p N_A_M1010_g 0.0157621f $X=13.2 $Y=4.07 $X2=4.58 $Y2=2.965
cc_85 N_VPB_M1000_b N_A_M1011_g 0.040726f $X=-0.33 $Y=1.885 $X2=5.36 $Y2=2.965
cc_86 VPB N_A_M1011_g 0.00970178f $X=0 $Y=3.955 $X2=5.36 $Y2=2.965
cc_87 N_VPB_c_69_p N_A_M1011_g 0.0157621f $X=13.2 $Y=4.07 $X2=5.36 $Y2=2.965
cc_88 N_VPB_M1000_b N_A_M1014_g 0.040726f $X=-0.33 $Y=1.885 $X2=6.14 $Y2=2.965
cc_89 VPB N_A_M1014_g 0.00970178f $X=0 $Y=3.955 $X2=6.14 $Y2=2.965
cc_90 N_VPB_c_69_p N_A_M1014_g 0.0157621f $X=13.2 $Y=4.07 $X2=6.14 $Y2=2.965
cc_91 N_VPB_M1000_b N_A_M1015_g 0.040726f $X=-0.33 $Y=1.885 $X2=6.92 $Y2=2.965
cc_92 VPB N_A_M1015_g 0.00970178f $X=0 $Y=3.955 $X2=6.92 $Y2=2.965
cc_93 N_VPB_c_69_p N_A_M1015_g 0.0157621f $X=13.2 $Y=4.07 $X2=6.92 $Y2=2.965
cc_94 N_VPB_M1000_b N_A_M1017_g 0.040726f $X=-0.33 $Y=1.885 $X2=7.7 $Y2=2.965
cc_95 VPB N_A_M1017_g 0.00970178f $X=0 $Y=3.955 $X2=7.7 $Y2=2.965
cc_96 N_VPB_c_69_p N_A_M1017_g 0.0157621f $X=13.2 $Y=4.07 $X2=7.7 $Y2=2.965
cc_97 N_VPB_M1000_b N_A_M1019_g 0.040726f $X=-0.33 $Y=1.885 $X2=8.48 $Y2=2.965
cc_98 VPB N_A_M1019_g 0.00970178f $X=0 $Y=3.955 $X2=8.48 $Y2=2.965
cc_99 N_VPB_c_69_p N_A_M1019_g 0.0157621f $X=13.2 $Y=4.07 $X2=8.48 $Y2=2.965
cc_100 N_VPB_M1000_b N_A_M1022_g 0.040726f $X=-0.33 $Y=1.885 $X2=9.26 $Y2=2.965
cc_101 VPB N_A_M1022_g 0.00970178f $X=0 $Y=3.955 $X2=9.26 $Y2=2.965
cc_102 N_VPB_c_69_p N_A_M1022_g 0.0157621f $X=13.2 $Y=4.07 $X2=9.26 $Y2=2.965
cc_103 N_VPB_M1000_b N_A_M1024_g 0.040726f $X=-0.33 $Y=1.885 $X2=10.04 $Y2=2.965
cc_104 VPB N_A_M1024_g 0.00970178f $X=0 $Y=3.955 $X2=10.04 $Y2=2.965
cc_105 N_VPB_c_69_p N_A_M1024_g 0.0157621f $X=13.2 $Y=4.07 $X2=10.04 $Y2=2.965
cc_106 N_VPB_M1000_b N_A_M1026_g 0.040726f $X=-0.33 $Y=1.885 $X2=10.82 $Y2=2.965
cc_107 VPB N_A_M1026_g 0.00970178f $X=0 $Y=3.955 $X2=10.82 $Y2=2.965
cc_108 N_VPB_c_69_p N_A_M1026_g 0.0157621f $X=13.2 $Y=4.07 $X2=10.82 $Y2=2.965
cc_109 N_VPB_M1000_b N_A_M1027_g 0.040726f $X=-0.33 $Y=1.885 $X2=11.6 $Y2=2.965
cc_110 VPB N_A_M1027_g 0.00970178f $X=0 $Y=3.955 $X2=11.6 $Y2=2.965
cc_111 N_VPB_c_69_p N_A_M1027_g 0.0157621f $X=13.2 $Y=4.07 $X2=11.6 $Y2=2.965
cc_112 N_VPB_M1000_b N_A_c_200_n 0.209261f $X=-0.33 $Y=1.885 $X2=12.375
+ $Y2=1.565
cc_113 N_VPB_M1000_b N_A_M1029_g 0.0505482f $X=-0.33 $Y=1.885 $X2=12.38
+ $Y2=2.965
cc_114 VPB N_A_M1029_g 0.00970178f $X=0 $Y=3.955 $X2=12.38 $Y2=2.965
cc_115 N_VPB_c_69_p N_A_M1029_g 0.0159934f $X=13.2 $Y=4.07 $X2=12.38 $Y2=2.965
cc_116 N_VPB_M1000_b N_VPWR_c_534_n 0.0702832f $X=-0.33 $Y=1.885 $X2=3.795
+ $Y2=1.08
cc_117 VPB N_VPWR_c_534_n 0.00200674f $X=0 $Y=3.955 $X2=3.795 $Y2=1.08
cc_118 N_VPB_c_69_p N_VPWR_c_534_n 0.0270143f $X=13.2 $Y=4.07 $X2=3.795 $Y2=1.08
cc_119 N_VPB_M1000_b N_VPWR_c_537_n 0.00369605f $X=-0.33 $Y=1.885 $X2=4.58
+ $Y2=2.965
cc_120 VPB N_VPWR_c_537_n 0.00377602f $X=0 $Y=3.955 $X2=4.58 $Y2=2.965
cc_121 N_VPB_c_69_p N_VPWR_c_537_n 0.0445179f $X=13.2 $Y=4.07 $X2=4.58 $Y2=2.965
cc_122 N_VPB_M1000_b N_VPWR_c_540_n 0.00369605f $X=-0.33 $Y=1.885 $X2=6.135
+ $Y2=1.08
cc_123 VPB N_VPWR_c_540_n 0.00377602f $X=0 $Y=3.955 $X2=6.135 $Y2=1.08
cc_124 N_VPB_c_69_p N_VPWR_c_540_n 0.0445179f $X=13.2 $Y=4.07 $X2=6.135 $Y2=1.08
cc_125 N_VPB_M1000_b N_VPWR_c_543_n 0.00369605f $X=-0.33 $Y=1.885 $X2=6.92
+ $Y2=2.965
cc_126 VPB N_VPWR_c_543_n 0.00377602f $X=0 $Y=3.955 $X2=6.92 $Y2=2.965
cc_127 N_VPB_c_69_p N_VPWR_c_543_n 0.0445179f $X=13.2 $Y=4.07 $X2=6.92 $Y2=2.965
cc_128 N_VPB_M1000_b N_VPWR_c_546_n 0.00369605f $X=-0.33 $Y=1.885 $X2=8.475
+ $Y2=1.08
cc_129 VPB N_VPWR_c_546_n 0.00377602f $X=0 $Y=3.955 $X2=8.475 $Y2=1.08
cc_130 N_VPB_c_69_p N_VPWR_c_546_n 0.0445179f $X=13.2 $Y=4.07 $X2=8.475 $Y2=1.08
cc_131 N_VPB_M1000_b N_VPWR_c_549_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_549_n 0.00377602f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_133 N_VPB_c_69_p N_VPWR_c_549_n 0.0445179f $X=13.2 $Y=4.07 $X2=0 $Y2=0
cc_134 N_VPB_M1000_b N_VPWR_c_552_n 0.00369605f $X=-0.33 $Y=1.885 $X2=10.82
+ $Y2=2.005
cc_135 VPB N_VPWR_c_552_n 0.00377602f $X=0 $Y=3.955 $X2=10.82 $Y2=2.005
cc_136 N_VPB_c_69_p N_VPWR_c_552_n 0.0445179f $X=13.2 $Y=4.07 $X2=10.82
+ $Y2=2.005
cc_137 N_VPB_M1000_b N_VPWR_c_555_n 0.00369605f $X=-0.33 $Y=1.885 $X2=12.375
+ $Y2=1.565
cc_138 VPB N_VPWR_c_555_n 0.00377602f $X=0 $Y=3.955 $X2=12.375 $Y2=1.565
cc_139 N_VPB_c_69_p N_VPWR_c_555_n 0.0445179f $X=13.2 $Y=4.07 $X2=12.375
+ $Y2=1.565
cc_140 N_VPB_M1000_b N_VPWR_c_558_n 0.0689428f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_558_n 0.00227374f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_142 N_VPB_c_69_p N_VPWR_c_558_n 0.0216668f $X=13.2 $Y=4.07 $X2=0 $Y2=0
cc_143 N_VPB_M1000_b N_VPWR_c_561_n 0.0778476f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_561_n 1.42384f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_145 N_VPB_c_69_p N_VPWR_c_561_n 0.0594722f $X=13.2 $Y=4.07 $X2=0 $Y2=0
cc_146 N_VPB_M1000_b N_Y_c_693_n 0.00125033f $X=-0.33 $Y=1.885 $X2=7.695
+ $Y2=1.08
cc_147 VPB N_Y_c_693_n 0.00108855f $X=0 $Y=3.955 $X2=7.695 $Y2=1.08
cc_148 N_VPB_c_69_p N_Y_c_693_n 0.0171423f $X=13.2 $Y=4.07 $X2=7.695 $Y2=1.08
cc_149 N_VPB_M1000_b N_Y_c_696_n 0.00125033f $X=-0.33 $Y=1.885 $X2=8.48
+ $Y2=2.965
cc_150 VPB N_Y_c_696_n 0.00108855f $X=0 $Y=3.955 $X2=8.48 $Y2=2.965
cc_151 N_VPB_c_69_p N_Y_c_696_n 0.0171423f $X=13.2 $Y=4.07 $X2=8.48 $Y2=2.965
cc_152 N_VPB_M1000_b N_Y_c_699_n 0.00125033f $X=-0.33 $Y=1.885 $X2=10.035
+ $Y2=1.08
cc_153 VPB N_Y_c_699_n 0.00108855f $X=0 $Y=3.955 $X2=10.035 $Y2=1.08
cc_154 N_VPB_c_69_p N_Y_c_699_n 0.0171423f $X=13.2 $Y=4.07 $X2=10.035 $Y2=1.08
cc_155 N_VPB_M1000_b N_Y_c_702_n 0.00125033f $X=-0.33 $Y=1.885 $X2=10.82
+ $Y2=2.965
cc_156 VPB N_Y_c_702_n 0.00108855f $X=0 $Y=3.955 $X2=10.82 $Y2=2.965
cc_157 N_VPB_c_69_p N_Y_c_702_n 0.0171423f $X=13.2 $Y=4.07 $X2=10.82 $Y2=2.965
cc_158 N_VPB_M1000_b N_Y_c_705_n 0.00125033f $X=-0.33 $Y=1.885 $X2=12.375
+ $Y2=1.565
cc_159 VPB N_Y_c_705_n 0.00108855f $X=0 $Y=3.955 $X2=12.375 $Y2=1.565
cc_160 N_VPB_c_69_p N_Y_c_705_n 0.0171423f $X=13.2 $Y=4.07 $X2=12.375 $Y2=1.565
cc_161 N_VPB_M1000_b N_Y_c_708_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_162 VPB N_Y_c_708_n 0.00108855f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_163 N_VPB_c_69_p N_Y_c_708_n 0.0171423f $X=13.2 $Y=4.07 $X2=0 $Y2=0
cc_164 N_VPB_M1000_b N_Y_c_711_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_165 VPB N_Y_c_711_n 0.00108855f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_166 N_VPB_c_69_p N_Y_c_711_n 0.0171423f $X=13.2 $Y=4.07 $X2=0 $Y2=0
cc_167 N_VPB_M1000_b N_Y_c_714_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_168 VPB N_Y_c_714_n 0.00108855f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_169 N_VPB_c_69_p N_Y_c_714_n 0.0171423f $X=13.2 $Y=4.07 $X2=0 $Y2=0
cc_170 N_A_M1000_g N_VPWR_c_534_n 0.0746134f $X=0.68 $Y=2.965 $X2=0 $Y2=0
cc_171 N_A_M1001_g N_VPWR_c_534_n 6.26267e-19 $X=1.46 $Y=2.965 $X2=0 $Y2=0
cc_172 N_A_c_200_n N_VPWR_c_534_n 2.41927e-19 $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_173 N_A_M1000_g N_VPWR_c_537_n 6.39823e-19 $X=0.68 $Y=2.965 $X2=0 $Y2=0
cc_174 N_A_M1001_g N_VPWR_c_537_n 0.0748611f $X=1.46 $Y=2.965 $X2=0 $Y2=0
cc_175 N_A_M1004_g N_VPWR_c_537_n 0.0731299f $X=2.24 $Y=2.965 $X2=0 $Y2=0
cc_176 N_A_M1008_g N_VPWR_c_537_n 6.24063e-19 $X=3.02 $Y=2.965 $X2=0 $Y2=0
cc_177 N_A_c_200_n N_VPWR_c_537_n 0.00265364f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_178 N_A_c_202_n N_VPWR_c_537_n 0.0382003f $X=2.04 $Y=1.665 $X2=0 $Y2=0
cc_179 N_A_c_210_n N_VPWR_c_537_n 0.00287773f $X=2.07 $Y=1.665 $X2=0 $Y2=0
cc_180 N_A_c_275_p N_VPWR_c_537_n 5.94054e-19 $X=3.085 $Y=1.665 $X2=0 $Y2=0
cc_181 N_A_M1004_g N_VPWR_c_540_n 6.39823e-19 $X=2.24 $Y=2.965 $X2=0 $Y2=0
cc_182 N_A_M1008_g N_VPWR_c_540_n 0.0748208f $X=3.02 $Y=2.965 $X2=0 $Y2=0
cc_183 N_A_M1009_g N_VPWR_c_540_n 0.0731305f $X=3.8 $Y=2.965 $X2=0 $Y2=0
cc_184 N_A_M1010_g N_VPWR_c_540_n 6.24063e-19 $X=4.58 $Y=2.965 $X2=0 $Y2=0
cc_185 N_A_c_200_n N_VPWR_c_540_n 0.00265364f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_186 N_A_c_203_n N_VPWR_c_540_n 0.0373217f $X=3.59 $Y=1.665 $X2=0 $Y2=0
cc_187 N_A_c_275_p N_VPWR_c_540_n 7.08785e-19 $X=3.085 $Y=1.665 $X2=0 $Y2=0
cc_188 N_A_c_283_p N_VPWR_c_540_n 0.00287695f $X=3.2 $Y=1.665 $X2=0 $Y2=0
cc_189 N_A_c_284_p N_VPWR_c_540_n 6.5142e-19 $X=4.645 $Y=1.665 $X2=0 $Y2=0
cc_190 N_A_M1009_g N_VPWR_c_543_n 6.39823e-19 $X=3.8 $Y=2.965 $X2=0 $Y2=0
cc_191 N_A_M1010_g N_VPWR_c_543_n 0.0748208f $X=4.58 $Y=2.965 $X2=0 $Y2=0
cc_192 N_A_M1011_g N_VPWR_c_543_n 0.0731305f $X=5.36 $Y=2.965 $X2=0 $Y2=0
cc_193 N_A_M1014_g N_VPWR_c_543_n 6.24063e-19 $X=6.14 $Y=2.965 $X2=0 $Y2=0
cc_194 N_A_c_200_n N_VPWR_c_543_n 0.00265364f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_195 N_A_c_204_n N_VPWR_c_543_n 0.0373217f $X=5.15 $Y=1.665 $X2=0 $Y2=0
cc_196 N_A_c_284_p N_VPWR_c_543_n 7.08785e-19 $X=4.645 $Y=1.665 $X2=0 $Y2=0
cc_197 N_A_c_292_p N_VPWR_c_543_n 0.00287695f $X=4.76 $Y=1.665 $X2=0 $Y2=0
cc_198 N_A_c_293_p N_VPWR_c_543_n 6.5142e-19 $X=6.205 $Y=1.665 $X2=0 $Y2=0
cc_199 N_A_M1011_g N_VPWR_c_546_n 6.39823e-19 $X=5.36 $Y=2.965 $X2=0 $Y2=0
cc_200 N_A_M1014_g N_VPWR_c_546_n 0.0748208f $X=6.14 $Y=2.965 $X2=0 $Y2=0
cc_201 N_A_M1015_g N_VPWR_c_546_n 0.0731305f $X=6.92 $Y=2.965 $X2=0 $Y2=0
cc_202 N_A_M1017_g N_VPWR_c_546_n 6.24063e-19 $X=7.7 $Y=2.965 $X2=0 $Y2=0
cc_203 N_A_c_200_n N_VPWR_c_546_n 0.00265364f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_204 N_A_c_205_n N_VPWR_c_546_n 0.0373217f $X=6.71 $Y=1.665 $X2=0 $Y2=0
cc_205 N_A_c_293_p N_VPWR_c_546_n 7.08785e-19 $X=6.205 $Y=1.665 $X2=0 $Y2=0
cc_206 N_A_c_301_p N_VPWR_c_546_n 0.00287695f $X=6.32 $Y=1.665 $X2=0 $Y2=0
cc_207 N_A_c_302_p N_VPWR_c_546_n 6.5142e-19 $X=7.765 $Y=1.665 $X2=0 $Y2=0
cc_208 N_A_M1015_g N_VPWR_c_549_n 6.39823e-19 $X=6.92 $Y=2.965 $X2=0 $Y2=0
cc_209 N_A_M1017_g N_VPWR_c_549_n 0.0748208f $X=7.7 $Y=2.965 $X2=0 $Y2=0
cc_210 N_A_M1019_g N_VPWR_c_549_n 0.0731305f $X=8.48 $Y=2.965 $X2=0 $Y2=0
cc_211 N_A_M1022_g N_VPWR_c_549_n 6.24063e-19 $X=9.26 $Y=2.965 $X2=0 $Y2=0
cc_212 N_A_c_200_n N_VPWR_c_549_n 0.00265364f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_213 N_A_c_206_n N_VPWR_c_549_n 0.0373217f $X=8.27 $Y=1.665 $X2=0 $Y2=0
cc_214 N_A_c_302_p N_VPWR_c_549_n 7.08785e-19 $X=7.765 $Y=1.665 $X2=0 $Y2=0
cc_215 N_A_c_310_p N_VPWR_c_549_n 0.00287695f $X=7.88 $Y=1.665 $X2=0 $Y2=0
cc_216 N_A_c_311_p N_VPWR_c_549_n 6.5142e-19 $X=9.325 $Y=1.665 $X2=0 $Y2=0
cc_217 N_A_M1019_g N_VPWR_c_552_n 6.39823e-19 $X=8.48 $Y=2.965 $X2=0 $Y2=0
cc_218 N_A_M1022_g N_VPWR_c_552_n 0.0748208f $X=9.26 $Y=2.965 $X2=0 $Y2=0
cc_219 N_A_M1024_g N_VPWR_c_552_n 0.0731305f $X=10.04 $Y=2.965 $X2=0 $Y2=0
cc_220 N_A_M1026_g N_VPWR_c_552_n 6.24063e-19 $X=10.82 $Y=2.965 $X2=0 $Y2=0
cc_221 N_A_c_200_n N_VPWR_c_552_n 0.00265364f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_222 N_A_c_207_n N_VPWR_c_552_n 0.0373217f $X=9.83 $Y=1.665 $X2=0 $Y2=0
cc_223 N_A_c_311_p N_VPWR_c_552_n 7.08785e-19 $X=9.325 $Y=1.665 $X2=0 $Y2=0
cc_224 N_A_c_319_p N_VPWR_c_552_n 0.00287695f $X=9.44 $Y=1.665 $X2=0 $Y2=0
cc_225 N_A_c_320_p N_VPWR_c_552_n 6.5142e-19 $X=10.885 $Y=1.665 $X2=0 $Y2=0
cc_226 N_A_M1024_g N_VPWR_c_555_n 6.39823e-19 $X=10.04 $Y=2.965 $X2=0 $Y2=0
cc_227 N_A_M1026_g N_VPWR_c_555_n 0.0748208f $X=10.82 $Y=2.965 $X2=0 $Y2=0
cc_228 N_A_M1027_g N_VPWR_c_555_n 0.0731643f $X=11.6 $Y=2.965 $X2=0 $Y2=0
cc_229 N_A_c_200_n N_VPWR_c_555_n 0.00265364f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_230 N_A_M1029_g N_VPWR_c_555_n 6.24063e-19 $X=12.38 $Y=2.965 $X2=0 $Y2=0
cc_231 N_A_c_208_n N_VPWR_c_555_n 0.0380692f $X=11.39 $Y=1.665 $X2=0 $Y2=0
cc_232 N_A_c_320_p N_VPWR_c_555_n 7.08785e-19 $X=10.885 $Y=1.665 $X2=0 $Y2=0
cc_233 N_A_c_328_p N_VPWR_c_555_n 0.00287773f $X=11 $Y=1.665 $X2=0 $Y2=0
cc_234 N_A_M1027_g N_VPWR_c_558_n 5.15209e-19 $X=11.6 $Y=2.965 $X2=0 $Y2=0
cc_235 N_A_M1029_g N_VPWR_c_558_n 0.0847648f $X=12.38 $Y=2.965 $X2=0 $Y2=0
cc_236 N_A_M1000_g N_VPWR_c_561_n 0.0142508f $X=0.68 $Y=2.965 $X2=0 $Y2=0
cc_237 N_A_M1001_g N_VPWR_c_561_n 0.00965647f $X=1.46 $Y=2.965 $X2=0 $Y2=0
cc_238 N_A_M1004_g N_VPWR_c_561_n 0.00965647f $X=2.24 $Y=2.965 $X2=0 $Y2=0
cc_239 N_A_M1008_g N_VPWR_c_561_n 0.00965647f $X=3.02 $Y=2.965 $X2=0 $Y2=0
cc_240 N_A_M1009_g N_VPWR_c_561_n 0.00965647f $X=3.8 $Y=2.965 $X2=0 $Y2=0
cc_241 N_A_M1010_g N_VPWR_c_561_n 0.00965647f $X=4.58 $Y=2.965 $X2=0 $Y2=0
cc_242 N_A_M1011_g N_VPWR_c_561_n 0.00965647f $X=5.36 $Y=2.965 $X2=0 $Y2=0
cc_243 N_A_M1014_g N_VPWR_c_561_n 0.00965647f $X=6.14 $Y=2.965 $X2=0 $Y2=0
cc_244 N_A_M1015_g N_VPWR_c_561_n 0.00965647f $X=6.92 $Y=2.965 $X2=0 $Y2=0
cc_245 N_A_M1017_g N_VPWR_c_561_n 0.00965647f $X=7.7 $Y=2.965 $X2=0 $Y2=0
cc_246 N_A_M1019_g N_VPWR_c_561_n 0.00965647f $X=8.48 $Y=2.965 $X2=0 $Y2=0
cc_247 N_A_M1022_g N_VPWR_c_561_n 0.00965647f $X=9.26 $Y=2.965 $X2=0 $Y2=0
cc_248 N_A_M1024_g N_VPWR_c_561_n 0.00965647f $X=10.04 $Y=2.965 $X2=0 $Y2=0
cc_249 N_A_M1026_g N_VPWR_c_561_n 0.00965647f $X=10.82 $Y=2.965 $X2=0 $Y2=0
cc_250 N_A_M1027_g N_VPWR_c_561_n 0.00965647f $X=11.6 $Y=2.965 $X2=0 $Y2=0
cc_251 N_A_M1029_g N_VPWR_c_561_n 0.0116277f $X=12.38 $Y=2.965 $X2=0 $Y2=0
cc_252 N_A_c_170_n N_Y_c_693_n 0.0196155f $X=0.675 $Y=1.565 $X2=0 $Y2=0
cc_253 N_A_M1000_g N_Y_c_693_n 0.0425154f $X=0.68 $Y=2.965 $X2=0 $Y2=0
cc_254 N_A_c_172_n N_Y_c_693_n 0.0189908f $X=1.455 $Y=1.565 $X2=0 $Y2=0
cc_255 N_A_M1001_g N_Y_c_693_n 0.0348822f $X=1.46 $Y=2.965 $X2=0 $Y2=0
cc_256 N_A_c_200_n N_Y_c_693_n 0.0481037f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_257 N_A_c_202_n N_Y_c_693_n 0.0251266f $X=2.04 $Y=1.665 $X2=0 $Y2=0
cc_258 N_A_c_210_n N_Y_c_693_n 0.00168021f $X=2.07 $Y=1.665 $X2=0 $Y2=0
cc_259 N_A_c_174_n N_Y_c_696_n 0.0189824f $X=2.235 $Y=1.565 $X2=0 $Y2=0
cc_260 N_A_M1004_g N_Y_c_696_n 0.0365608f $X=2.24 $Y=2.965 $X2=0 $Y2=0
cc_261 N_A_c_176_n N_Y_c_696_n 0.018988f $X=3.015 $Y=1.565 $X2=0 $Y2=0
cc_262 N_A_M1008_g N_Y_c_696_n 0.0348822f $X=3.02 $Y=2.965 $X2=0 $Y2=0
cc_263 N_A_c_200_n N_Y_c_696_n 0.0361022f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_264 N_A_c_202_n N_Y_c_696_n 0.0235891f $X=2.04 $Y=1.665 $X2=0 $Y2=0
cc_265 N_A_c_203_n N_Y_c_696_n 0.0236027f $X=3.59 $Y=1.665 $X2=0 $Y2=0
cc_266 N_A_c_275_p N_Y_c_696_n 0.0375764f $X=3.085 $Y=1.665 $X2=0 $Y2=0
cc_267 N_A_c_362_p N_Y_c_696_n 8.46898e-19 $X=2.185 $Y=1.665 $X2=0 $Y2=0
cc_268 N_A_c_283_p N_Y_c_696_n 8.22499e-19 $X=3.2 $Y=1.665 $X2=0 $Y2=0
cc_269 N_A_c_178_n N_Y_c_699_n 0.0189852f $X=3.795 $Y=1.565 $X2=0 $Y2=0
cc_270 N_A_M1009_g N_Y_c_699_n 0.0365608f $X=3.8 $Y=2.965 $X2=0 $Y2=0
cc_271 N_A_c_180_n N_Y_c_699_n 0.018988f $X=4.575 $Y=1.565 $X2=0 $Y2=0
cc_272 N_A_M1010_g N_Y_c_699_n 0.0348822f $X=4.58 $Y=2.965 $X2=0 $Y2=0
cc_273 N_A_c_200_n N_Y_c_699_n 0.036103f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_274 N_A_c_203_n N_Y_c_699_n 0.0235959f $X=3.59 $Y=1.665 $X2=0 $Y2=0
cc_275 N_A_c_204_n N_Y_c_699_n 0.0236027f $X=5.15 $Y=1.665 $X2=0 $Y2=0
cc_276 N_A_c_284_p N_Y_c_699_n 0.0375764f $X=4.645 $Y=1.665 $X2=0 $Y2=0
cc_277 N_A_c_372_p N_Y_c_699_n 8.34534e-19 $X=3.735 $Y=1.665 $X2=0 $Y2=0
cc_278 N_A_c_292_p N_Y_c_699_n 8.22499e-19 $X=4.76 $Y=1.665 $X2=0 $Y2=0
cc_279 N_A_c_182_n N_Y_c_702_n 0.0189852f $X=5.355 $Y=1.565 $X2=0 $Y2=0
cc_280 N_A_M1011_g N_Y_c_702_n 0.0365608f $X=5.36 $Y=2.965 $X2=0 $Y2=0
cc_281 N_A_c_184_n N_Y_c_702_n 0.018988f $X=6.135 $Y=1.565 $X2=0 $Y2=0
cc_282 N_A_M1014_g N_Y_c_702_n 0.0348822f $X=6.14 $Y=2.965 $X2=0 $Y2=0
cc_283 N_A_c_200_n N_Y_c_702_n 0.036103f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_284 N_A_c_204_n N_Y_c_702_n 0.0235959f $X=5.15 $Y=1.665 $X2=0 $Y2=0
cc_285 N_A_c_205_n N_Y_c_702_n 0.0236027f $X=6.71 $Y=1.665 $X2=0 $Y2=0
cc_286 N_A_c_293_p N_Y_c_702_n 0.0375764f $X=6.205 $Y=1.665 $X2=0 $Y2=0
cc_287 N_A_c_382_p N_Y_c_702_n 8.34534e-19 $X=5.295 $Y=1.665 $X2=0 $Y2=0
cc_288 N_A_c_301_p N_Y_c_702_n 8.22499e-19 $X=6.32 $Y=1.665 $X2=0 $Y2=0
cc_289 N_A_c_186_n N_Y_c_705_n 0.0189852f $X=6.915 $Y=1.565 $X2=0 $Y2=0
cc_290 N_A_M1015_g N_Y_c_705_n 0.0365608f $X=6.92 $Y=2.965 $X2=0 $Y2=0
cc_291 N_A_c_188_n N_Y_c_705_n 0.018988f $X=7.695 $Y=1.565 $X2=0 $Y2=0
cc_292 N_A_M1017_g N_Y_c_705_n 0.0348822f $X=7.7 $Y=2.965 $X2=0 $Y2=0
cc_293 N_A_c_200_n N_Y_c_705_n 0.036103f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_294 N_A_c_205_n N_Y_c_705_n 0.0235959f $X=6.71 $Y=1.665 $X2=0 $Y2=0
cc_295 N_A_c_206_n N_Y_c_705_n 0.0236027f $X=8.27 $Y=1.665 $X2=0 $Y2=0
cc_296 N_A_c_302_p N_Y_c_705_n 0.0375764f $X=7.765 $Y=1.665 $X2=0 $Y2=0
cc_297 N_A_c_392_p N_Y_c_705_n 8.34534e-19 $X=6.855 $Y=1.665 $X2=0 $Y2=0
cc_298 N_A_c_310_p N_Y_c_705_n 8.22499e-19 $X=7.88 $Y=1.665 $X2=0 $Y2=0
cc_299 N_A_c_190_n N_Y_c_708_n 0.0189852f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_300 N_A_M1019_g N_Y_c_708_n 0.0365608f $X=8.48 $Y=2.965 $X2=0 $Y2=0
cc_301 N_A_c_192_n N_Y_c_708_n 0.018988f $X=9.255 $Y=1.565 $X2=0 $Y2=0
cc_302 N_A_M1022_g N_Y_c_708_n 0.0348822f $X=9.26 $Y=2.965 $X2=0 $Y2=0
cc_303 N_A_c_200_n N_Y_c_708_n 0.036103f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_304 N_A_c_206_n N_Y_c_708_n 0.0235959f $X=8.27 $Y=1.665 $X2=0 $Y2=0
cc_305 N_A_c_207_n N_Y_c_708_n 0.0236027f $X=9.83 $Y=1.665 $X2=0 $Y2=0
cc_306 N_A_c_311_p N_Y_c_708_n 0.0375764f $X=9.325 $Y=1.665 $X2=0 $Y2=0
cc_307 N_A_c_402_p N_Y_c_708_n 8.34534e-19 $X=8.415 $Y=1.665 $X2=0 $Y2=0
cc_308 N_A_c_319_p N_Y_c_708_n 8.22499e-19 $X=9.44 $Y=1.665 $X2=0 $Y2=0
cc_309 N_A_c_194_n N_Y_c_711_n 0.0189852f $X=10.035 $Y=1.565 $X2=0 $Y2=0
cc_310 N_A_M1024_g N_Y_c_711_n 0.0365608f $X=10.04 $Y=2.965 $X2=0 $Y2=0
cc_311 N_A_c_196_n N_Y_c_711_n 0.018988f $X=10.815 $Y=1.565 $X2=0 $Y2=0
cc_312 N_A_M1026_g N_Y_c_711_n 0.0348822f $X=10.82 $Y=2.965 $X2=0 $Y2=0
cc_313 N_A_c_200_n N_Y_c_711_n 0.036103f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_314 N_A_c_207_n N_Y_c_711_n 0.0235959f $X=9.83 $Y=1.665 $X2=0 $Y2=0
cc_315 N_A_c_208_n N_Y_c_711_n 0.0236027f $X=11.39 $Y=1.665 $X2=0 $Y2=0
cc_316 N_A_c_320_p N_Y_c_711_n 0.0375764f $X=10.885 $Y=1.665 $X2=0 $Y2=0
cc_317 N_A_c_412_p N_Y_c_711_n 8.34534e-19 $X=9.975 $Y=1.665 $X2=0 $Y2=0
cc_318 N_A_c_328_p N_Y_c_711_n 8.22499e-19 $X=11 $Y=1.665 $X2=0 $Y2=0
cc_319 N_A_c_198_n N_Y_c_714_n 0.0189852f $X=11.595 $Y=1.565 $X2=0 $Y2=0
cc_320 N_A_M1027_g N_Y_c_714_n 0.0365608f $X=11.6 $Y=2.965 $X2=0 $Y2=0
cc_321 N_A_c_200_n N_Y_c_714_n 0.067459f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_322 N_A_M1029_g N_Y_c_714_n 0.0372205f $X=12.38 $Y=2.965 $X2=0 $Y2=0
cc_323 N_A_c_208_n N_Y_c_714_n 0.0250621f $X=11.39 $Y=1.665 $X2=0 $Y2=0
cc_324 N_A_c_209_n N_Y_c_714_n 0.00174341f $X=11.39 $Y=1.665 $X2=0 $Y2=0
cc_325 N_A_M1001_g N_Y_c_790_n 0.014391f $X=1.46 $Y=2.965 $X2=0 $Y2=0
cc_326 N_A_M1004_g N_Y_c_790_n 0.014391f $X=2.24 $Y=2.965 $X2=0 $Y2=0
cc_327 N_A_c_202_n N_Y_c_790_n 0.00350242f $X=2.04 $Y=1.665 $X2=0 $Y2=0
cc_328 N_A_c_210_n N_Y_c_790_n 0.0256867f $X=2.07 $Y=1.665 $X2=0 $Y2=0
cc_329 N_A_M1008_g N_Y_c_794_n 0.014391f $X=3.02 $Y=2.965 $X2=0 $Y2=0
cc_330 N_A_M1009_g N_Y_c_794_n 0.014391f $X=3.8 $Y=2.965 $X2=0 $Y2=0
cc_331 N_A_c_203_n N_Y_c_794_n 0.00350242f $X=3.59 $Y=1.665 $X2=0 $Y2=0
cc_332 N_A_c_283_p N_Y_c_794_n 0.0256666f $X=3.2 $Y=1.665 $X2=0 $Y2=0
cc_333 N_A_c_275_p N_Y_c_798_n 0.0114767f $X=3.085 $Y=1.665 $X2=0 $Y2=0
cc_334 N_A_M1010_g N_Y_c_799_n 0.014391f $X=4.58 $Y=2.965 $X2=0 $Y2=0
cc_335 N_A_M1011_g N_Y_c_799_n 0.014391f $X=5.36 $Y=2.965 $X2=0 $Y2=0
cc_336 N_A_c_204_n N_Y_c_799_n 0.00350242f $X=5.15 $Y=1.665 $X2=0 $Y2=0
cc_337 N_A_c_292_p N_Y_c_799_n 0.0256666f $X=4.76 $Y=1.665 $X2=0 $Y2=0
cc_338 N_A_c_284_p N_Y_c_803_n 0.0114767f $X=4.645 $Y=1.665 $X2=0 $Y2=0
cc_339 N_A_M1014_g N_Y_c_804_n 0.014391f $X=6.14 $Y=2.965 $X2=0 $Y2=0
cc_340 N_A_M1015_g N_Y_c_804_n 0.014391f $X=6.92 $Y=2.965 $X2=0 $Y2=0
cc_341 N_A_c_205_n N_Y_c_804_n 0.00350242f $X=6.71 $Y=1.665 $X2=0 $Y2=0
cc_342 N_A_c_301_p N_Y_c_804_n 0.0256666f $X=6.32 $Y=1.665 $X2=0 $Y2=0
cc_343 N_A_c_293_p N_Y_c_808_n 0.0114767f $X=6.205 $Y=1.665 $X2=0 $Y2=0
cc_344 N_A_M1017_g N_Y_c_809_n 0.014391f $X=7.7 $Y=2.965 $X2=0 $Y2=0
cc_345 N_A_M1019_g N_Y_c_809_n 0.014391f $X=8.48 $Y=2.965 $X2=0 $Y2=0
cc_346 N_A_c_206_n N_Y_c_809_n 0.00350242f $X=8.27 $Y=1.665 $X2=0 $Y2=0
cc_347 N_A_c_310_p N_Y_c_809_n 0.0256666f $X=7.88 $Y=1.665 $X2=0 $Y2=0
cc_348 N_A_c_302_p N_Y_c_813_n 0.0114767f $X=7.765 $Y=1.665 $X2=0 $Y2=0
cc_349 N_A_M1022_g N_Y_c_814_n 0.014391f $X=9.26 $Y=2.965 $X2=0 $Y2=0
cc_350 N_A_M1024_g N_Y_c_814_n 0.014391f $X=10.04 $Y=2.965 $X2=0 $Y2=0
cc_351 N_A_c_207_n N_Y_c_814_n 0.00350242f $X=9.83 $Y=1.665 $X2=0 $Y2=0
cc_352 N_A_c_319_p N_Y_c_814_n 0.0256666f $X=9.44 $Y=1.665 $X2=0 $Y2=0
cc_353 N_A_c_311_p N_Y_c_818_n 0.0114767f $X=9.325 $Y=1.665 $X2=0 $Y2=0
cc_354 N_A_M1026_g N_Y_c_819_n 0.014391f $X=10.82 $Y=2.965 $X2=0 $Y2=0
cc_355 N_A_M1027_g N_Y_c_819_n 0.014391f $X=11.6 $Y=2.965 $X2=0 $Y2=0
cc_356 N_A_c_208_n N_Y_c_819_n 0.00350242f $X=11.39 $Y=1.665 $X2=0 $Y2=0
cc_357 N_A_c_328_p N_Y_c_819_n 0.0256867f $X=11 $Y=1.665 $X2=0 $Y2=0
cc_358 N_A_c_320_p N_Y_c_823_n 0.0114767f $X=10.885 $Y=1.665 $X2=0 $Y2=0
cc_359 N_A_c_170_n N_VGND_c_895_n 0.0521092f $X=0.675 $Y=1.565 $X2=0 $Y2=0
cc_360 N_A_c_172_n N_VGND_c_895_n 0.00113076f $X=1.455 $Y=1.565 $X2=0 $Y2=0
cc_361 N_A_c_170_n N_VGND_c_897_n 0.00111754f $X=0.675 $Y=1.565 $X2=0 $Y2=0
cc_362 N_A_c_172_n N_VGND_c_897_n 0.0479045f $X=1.455 $Y=1.565 $X2=0 $Y2=0
cc_363 N_A_c_174_n N_VGND_c_897_n 0.0475415f $X=2.235 $Y=1.565 $X2=0 $Y2=0
cc_364 N_A_c_176_n N_VGND_c_897_n 6.55742e-19 $X=3.015 $Y=1.565 $X2=0 $Y2=0
cc_365 N_A_c_200_n N_VGND_c_897_n 7.87671e-19 $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_366 N_A_c_202_n N_VGND_c_897_n 0.0584447f $X=2.04 $Y=1.665 $X2=0 $Y2=0
cc_367 N_A_c_210_n N_VGND_c_897_n 0.0171266f $X=2.07 $Y=1.665 $X2=0 $Y2=0
cc_368 N_A_c_275_p N_VGND_c_897_n 8.06456e-19 $X=3.085 $Y=1.665 $X2=0 $Y2=0
cc_369 N_A_c_174_n N_VGND_c_899_n 6.55742e-19 $X=2.235 $Y=1.565 $X2=0 $Y2=0
cc_370 N_A_c_176_n N_VGND_c_899_n 0.0475428f $X=3.015 $Y=1.565 $X2=0 $Y2=0
cc_371 N_A_c_178_n N_VGND_c_899_n 0.0475421f $X=3.795 $Y=1.565 $X2=0 $Y2=0
cc_372 N_A_c_180_n N_VGND_c_899_n 6.55742e-19 $X=4.575 $Y=1.565 $X2=0 $Y2=0
cc_373 N_A_c_200_n N_VGND_c_899_n 7.87671e-19 $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_374 N_A_c_203_n N_VGND_c_899_n 0.0574267f $X=3.59 $Y=1.665 $X2=0 $Y2=0
cc_375 N_A_c_275_p N_VGND_c_899_n 9.6243e-19 $X=3.085 $Y=1.665 $X2=0 $Y2=0
cc_376 N_A_c_283_p N_VGND_c_899_n 0.0171054f $X=3.2 $Y=1.665 $X2=0 $Y2=0
cc_377 N_A_c_284_p N_VGND_c_899_n 8.84443e-19 $X=4.645 $Y=1.665 $X2=0 $Y2=0
cc_378 N_A_c_178_n N_VGND_c_901_n 6.55742e-19 $X=3.795 $Y=1.565 $X2=0 $Y2=0
cc_379 N_A_c_180_n N_VGND_c_901_n 0.0475428f $X=4.575 $Y=1.565 $X2=0 $Y2=0
cc_380 N_A_c_182_n N_VGND_c_901_n 0.0475421f $X=5.355 $Y=1.565 $X2=0 $Y2=0
cc_381 N_A_c_184_n N_VGND_c_901_n 6.55742e-19 $X=6.135 $Y=1.565 $X2=0 $Y2=0
cc_382 N_A_c_200_n N_VGND_c_901_n 7.87671e-19 $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_383 N_A_c_204_n N_VGND_c_901_n 0.0574267f $X=5.15 $Y=1.665 $X2=0 $Y2=0
cc_384 N_A_c_284_p N_VGND_c_901_n 9.6243e-19 $X=4.645 $Y=1.665 $X2=0 $Y2=0
cc_385 N_A_c_292_p N_VGND_c_901_n 0.0171054f $X=4.76 $Y=1.665 $X2=0 $Y2=0
cc_386 N_A_c_293_p N_VGND_c_901_n 8.84443e-19 $X=6.205 $Y=1.665 $X2=0 $Y2=0
cc_387 N_A_c_182_n N_VGND_c_903_n 6.55742e-19 $X=5.355 $Y=1.565 $X2=0 $Y2=0
cc_388 N_A_c_184_n N_VGND_c_903_n 0.0475428f $X=6.135 $Y=1.565 $X2=0 $Y2=0
cc_389 N_A_c_186_n N_VGND_c_903_n 0.0475421f $X=6.915 $Y=1.565 $X2=0 $Y2=0
cc_390 N_A_c_188_n N_VGND_c_903_n 6.55742e-19 $X=7.695 $Y=1.565 $X2=0 $Y2=0
cc_391 N_A_c_200_n N_VGND_c_903_n 7.87671e-19 $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_392 N_A_c_205_n N_VGND_c_903_n 0.0574267f $X=6.71 $Y=1.665 $X2=0 $Y2=0
cc_393 N_A_c_293_p N_VGND_c_903_n 9.6243e-19 $X=6.205 $Y=1.665 $X2=0 $Y2=0
cc_394 N_A_c_301_p N_VGND_c_903_n 0.0171054f $X=6.32 $Y=1.665 $X2=0 $Y2=0
cc_395 N_A_c_302_p N_VGND_c_903_n 8.84443e-19 $X=7.765 $Y=1.665 $X2=0 $Y2=0
cc_396 N_A_c_186_n N_VGND_c_905_n 6.55742e-19 $X=6.915 $Y=1.565 $X2=0 $Y2=0
cc_397 N_A_c_188_n N_VGND_c_905_n 0.0475428f $X=7.695 $Y=1.565 $X2=0 $Y2=0
cc_398 N_A_c_190_n N_VGND_c_905_n 0.0475421f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_399 N_A_c_192_n N_VGND_c_905_n 6.55742e-19 $X=9.255 $Y=1.565 $X2=0 $Y2=0
cc_400 N_A_c_200_n N_VGND_c_905_n 7.87671e-19 $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_401 N_A_c_206_n N_VGND_c_905_n 0.0574267f $X=8.27 $Y=1.665 $X2=0 $Y2=0
cc_402 N_A_c_302_p N_VGND_c_905_n 9.6243e-19 $X=7.765 $Y=1.665 $X2=0 $Y2=0
cc_403 N_A_c_310_p N_VGND_c_905_n 0.0171054f $X=7.88 $Y=1.665 $X2=0 $Y2=0
cc_404 N_A_c_311_p N_VGND_c_905_n 8.84443e-19 $X=9.325 $Y=1.665 $X2=0 $Y2=0
cc_405 N_A_c_190_n N_VGND_c_907_n 6.55742e-19 $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_406 N_A_c_192_n N_VGND_c_907_n 0.0475428f $X=9.255 $Y=1.565 $X2=0 $Y2=0
cc_407 N_A_c_194_n N_VGND_c_907_n 0.0475421f $X=10.035 $Y=1.565 $X2=0 $Y2=0
cc_408 N_A_c_196_n N_VGND_c_907_n 6.55742e-19 $X=10.815 $Y=1.565 $X2=0 $Y2=0
cc_409 N_A_c_200_n N_VGND_c_907_n 7.87671e-19 $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_410 N_A_c_207_n N_VGND_c_907_n 0.0574267f $X=9.83 $Y=1.665 $X2=0 $Y2=0
cc_411 N_A_c_311_p N_VGND_c_907_n 9.6243e-19 $X=9.325 $Y=1.665 $X2=0 $Y2=0
cc_412 N_A_c_319_p N_VGND_c_907_n 0.0171054f $X=9.44 $Y=1.665 $X2=0 $Y2=0
cc_413 N_A_c_320_p N_VGND_c_907_n 8.84443e-19 $X=10.885 $Y=1.665 $X2=0 $Y2=0
cc_414 N_A_c_194_n N_VGND_c_909_n 6.55742e-19 $X=10.035 $Y=1.565 $X2=0 $Y2=0
cc_415 N_A_c_196_n N_VGND_c_909_n 0.0475428f $X=10.815 $Y=1.565 $X2=0 $Y2=0
cc_416 N_A_c_198_n N_VGND_c_909_n 0.0476016f $X=11.595 $Y=1.565 $X2=0 $Y2=0
cc_417 N_A_c_200_n N_VGND_c_909_n 0.00144341f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_418 N_A_c_208_n N_VGND_c_909_n 0.058292f $X=11.39 $Y=1.665 $X2=0 $Y2=0
cc_419 N_A_c_320_p N_VGND_c_909_n 9.6243e-19 $X=10.885 $Y=1.665 $X2=0 $Y2=0
cc_420 N_A_c_328_p N_VGND_c_909_n 0.0171266f $X=11 $Y=1.665 $X2=0 $Y2=0
cc_421 N_A_c_198_n N_VGND_c_911_n 6.54796e-19 $X=11.595 $Y=1.565 $X2=0 $Y2=0
cc_422 N_A_c_200_n N_VGND_c_911_n 0.0604827f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_423 N_A_c_170_n N_VGND_c_913_n 0.0169491f $X=0.675 $Y=1.565 $X2=0 $Y2=0
cc_424 N_A_c_172_n N_VGND_c_913_n 0.0109655f $X=1.455 $Y=1.565 $X2=0 $Y2=0
cc_425 N_A_c_174_n N_VGND_c_913_n 0.0109655f $X=2.235 $Y=1.565 $X2=0 $Y2=0
cc_426 N_A_c_176_n N_VGND_c_913_n 0.0109655f $X=3.015 $Y=1.565 $X2=0 $Y2=0
cc_427 N_A_c_178_n N_VGND_c_913_n 0.0109655f $X=3.795 $Y=1.565 $X2=0 $Y2=0
cc_428 N_A_c_180_n N_VGND_c_913_n 0.0109655f $X=4.575 $Y=1.565 $X2=0 $Y2=0
cc_429 N_A_c_182_n N_VGND_c_913_n 0.0109655f $X=5.355 $Y=1.565 $X2=0 $Y2=0
cc_430 N_A_c_184_n N_VGND_c_913_n 0.0109655f $X=6.135 $Y=1.565 $X2=0 $Y2=0
cc_431 N_A_c_186_n N_VGND_c_913_n 0.0109655f $X=6.915 $Y=1.565 $X2=0 $Y2=0
cc_432 N_A_c_188_n N_VGND_c_913_n 0.0109655f $X=7.695 $Y=1.565 $X2=0 $Y2=0
cc_433 N_A_c_190_n N_VGND_c_913_n 0.0109655f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_434 N_A_c_192_n N_VGND_c_913_n 0.0109655f $X=9.255 $Y=1.565 $X2=0 $Y2=0
cc_435 N_A_c_194_n N_VGND_c_913_n 0.0109655f $X=10.035 $Y=1.565 $X2=0 $Y2=0
cc_436 N_A_c_196_n N_VGND_c_913_n 0.0109655f $X=10.815 $Y=1.565 $X2=0 $Y2=0
cc_437 N_A_c_198_n N_VGND_c_913_n 0.0109655f $X=11.595 $Y=1.565 $X2=0 $Y2=0
cc_438 N_A_c_200_n N_VGND_c_913_n 0.0109655f $X=12.375 $Y=1.565 $X2=0 $Y2=0
cc_439 N_VPWR_c_555_n Y 4.454e-19 $X=11.21 $Y=2.34 $X2=0 $Y2=0
cc_440 N_VPWR_c_558_n Y 0.00169694f $X=12.77 $Y=2.36 $X2=0 $Y2=0
cc_441 N_VPWR_c_534_n N_Y_c_693_n 0.0854647f $X=0.29 $Y=2.36 $X2=0 $Y2=0
cc_442 N_VPWR_c_537_n N_Y_c_693_n 0.118346f $X=1.85 $Y=2.34 $X2=0 $Y2=0
cc_443 N_VPWR_c_561_n N_Y_c_693_n 0.0389073f $X=12.81 $Y=3.56 $X2=0 $Y2=0
cc_444 N_VPWR_c_537_n N_Y_c_696_n 0.118355f $X=1.85 $Y=2.34 $X2=0 $Y2=0
cc_445 N_VPWR_c_540_n N_Y_c_696_n 0.118346f $X=3.41 $Y=2.34 $X2=0 $Y2=0
cc_446 N_VPWR_c_561_n N_Y_c_696_n 0.037804f $X=12.81 $Y=3.56 $X2=0 $Y2=0
cc_447 N_VPWR_c_540_n N_Y_c_699_n 0.118355f $X=3.41 $Y=2.34 $X2=0 $Y2=0
cc_448 N_VPWR_c_543_n N_Y_c_699_n 0.118346f $X=4.97 $Y=2.34 $X2=0 $Y2=0
cc_449 N_VPWR_c_561_n N_Y_c_699_n 0.037804f $X=12.81 $Y=3.56 $X2=0 $Y2=0
cc_450 N_VPWR_c_543_n N_Y_c_702_n 0.118355f $X=4.97 $Y=2.34 $X2=0 $Y2=0
cc_451 N_VPWR_c_546_n N_Y_c_702_n 0.118346f $X=6.53 $Y=2.34 $X2=0 $Y2=0
cc_452 N_VPWR_c_561_n N_Y_c_702_n 0.037804f $X=12.81 $Y=3.56 $X2=0 $Y2=0
cc_453 N_VPWR_c_546_n N_Y_c_705_n 0.118355f $X=6.53 $Y=2.34 $X2=0 $Y2=0
cc_454 N_VPWR_c_549_n N_Y_c_705_n 0.118346f $X=8.09 $Y=2.34 $X2=0 $Y2=0
cc_455 N_VPWR_c_561_n N_Y_c_705_n 0.037804f $X=12.81 $Y=3.56 $X2=0 $Y2=0
cc_456 N_VPWR_c_549_n N_Y_c_708_n 0.118355f $X=8.09 $Y=2.34 $X2=0 $Y2=0
cc_457 N_VPWR_c_552_n N_Y_c_708_n 0.118346f $X=9.65 $Y=2.34 $X2=0 $Y2=0
cc_458 N_VPWR_c_561_n N_Y_c_708_n 0.037804f $X=12.81 $Y=3.56 $X2=0 $Y2=0
cc_459 N_VPWR_c_552_n N_Y_c_711_n 0.118355f $X=9.65 $Y=2.34 $X2=0 $Y2=0
cc_460 N_VPWR_c_555_n N_Y_c_711_n 0.118346f $X=11.21 $Y=2.34 $X2=0 $Y2=0
cc_461 N_VPWR_c_561_n N_Y_c_711_n 0.037804f $X=12.81 $Y=3.56 $X2=0 $Y2=0
cc_462 N_VPWR_c_555_n N_Y_c_714_n 0.118355f $X=11.21 $Y=2.34 $X2=0 $Y2=0
cc_463 N_VPWR_c_558_n N_Y_c_714_n 0.113368f $X=12.77 $Y=2.36 $X2=0 $Y2=0
cc_464 N_VPWR_c_561_n N_Y_c_714_n 0.0392154f $X=12.81 $Y=3.56 $X2=0 $Y2=0
cc_465 N_VPWR_c_537_n N_Y_c_790_n 0.0838262f $X=1.85 $Y=2.34 $X2=0 $Y2=0
cc_466 N_VPWR_c_534_n N_Y_c_851_n 0.00157834f $X=0.29 $Y=2.36 $X2=0 $Y2=0
cc_467 N_VPWR_c_537_n N_Y_c_851_n 4.58442e-19 $X=1.85 $Y=2.34 $X2=0 $Y2=0
cc_468 N_VPWR_c_540_n N_Y_c_794_n 0.0838262f $X=3.41 $Y=2.34 $X2=0 $Y2=0
cc_469 N_VPWR_c_537_n N_Y_c_798_n 4.454e-19 $X=1.85 $Y=2.34 $X2=0 $Y2=0
cc_470 N_VPWR_c_540_n N_Y_c_798_n 4.58442e-19 $X=3.41 $Y=2.34 $X2=0 $Y2=0
cc_471 N_VPWR_c_543_n N_Y_c_799_n 0.0838262f $X=4.97 $Y=2.34 $X2=0 $Y2=0
cc_472 N_VPWR_c_540_n N_Y_c_803_n 4.454e-19 $X=3.41 $Y=2.34 $X2=0 $Y2=0
cc_473 N_VPWR_c_543_n N_Y_c_803_n 4.58442e-19 $X=4.97 $Y=2.34 $X2=0 $Y2=0
cc_474 N_VPWR_c_546_n N_Y_c_804_n 0.0838262f $X=6.53 $Y=2.34 $X2=0 $Y2=0
cc_475 N_VPWR_c_543_n N_Y_c_808_n 4.454e-19 $X=4.97 $Y=2.34 $X2=0 $Y2=0
cc_476 N_VPWR_c_546_n N_Y_c_808_n 4.58442e-19 $X=6.53 $Y=2.34 $X2=0 $Y2=0
cc_477 N_VPWR_c_549_n N_Y_c_809_n 0.0838262f $X=8.09 $Y=2.34 $X2=0 $Y2=0
cc_478 N_VPWR_c_546_n N_Y_c_813_n 4.454e-19 $X=6.53 $Y=2.34 $X2=0 $Y2=0
cc_479 N_VPWR_c_549_n N_Y_c_813_n 4.58442e-19 $X=8.09 $Y=2.34 $X2=0 $Y2=0
cc_480 N_VPWR_c_552_n N_Y_c_814_n 0.0838262f $X=9.65 $Y=2.34 $X2=0 $Y2=0
cc_481 N_VPWR_c_549_n N_Y_c_818_n 4.454e-19 $X=8.09 $Y=2.34 $X2=0 $Y2=0
cc_482 N_VPWR_c_552_n N_Y_c_818_n 4.58442e-19 $X=9.65 $Y=2.34 $X2=0 $Y2=0
cc_483 N_VPWR_c_555_n N_Y_c_819_n 0.0838262f $X=11.21 $Y=2.34 $X2=0 $Y2=0
cc_484 N_VPWR_c_552_n N_Y_c_823_n 4.454e-19 $X=9.65 $Y=2.34 $X2=0 $Y2=0
cc_485 N_VPWR_c_555_n N_Y_c_823_n 4.58442e-19 $X=11.21 $Y=2.34 $X2=0 $Y2=0
cc_486 N_Y_c_693_n N_VGND_c_895_n 0.0366134f $X=1.065 $Y=0.96 $X2=0 $Y2=0
cc_487 N_Y_c_693_n N_VGND_c_897_n 0.0476685f $X=1.065 $Y=0.96 $X2=0 $Y2=0
cc_488 N_Y_c_696_n N_VGND_c_897_n 0.0476685f $X=2.625 $Y=0.96 $X2=0 $Y2=0
cc_489 N_Y_c_696_n N_VGND_c_899_n 0.0476685f $X=2.625 $Y=0.96 $X2=0 $Y2=0
cc_490 N_Y_c_699_n N_VGND_c_899_n 0.0476685f $X=4.185 $Y=0.96 $X2=0 $Y2=0
cc_491 N_Y_c_699_n N_VGND_c_901_n 0.0476685f $X=4.185 $Y=0.96 $X2=0 $Y2=0
cc_492 N_Y_c_702_n N_VGND_c_901_n 0.0476685f $X=5.745 $Y=0.96 $X2=0 $Y2=0
cc_493 N_Y_c_702_n N_VGND_c_903_n 0.0476685f $X=5.745 $Y=0.96 $X2=0 $Y2=0
cc_494 N_Y_c_705_n N_VGND_c_903_n 0.0476685f $X=7.305 $Y=0.96 $X2=0 $Y2=0
cc_495 N_Y_c_705_n N_VGND_c_905_n 0.0476685f $X=7.305 $Y=0.96 $X2=0 $Y2=0
cc_496 N_Y_c_708_n N_VGND_c_905_n 0.0476685f $X=8.865 $Y=0.96 $X2=0 $Y2=0
cc_497 N_Y_c_708_n N_VGND_c_907_n 0.0476685f $X=8.865 $Y=0.96 $X2=0 $Y2=0
cc_498 N_Y_c_711_n N_VGND_c_907_n 0.0476685f $X=10.425 $Y=0.96 $X2=0 $Y2=0
cc_499 N_Y_c_711_n N_VGND_c_909_n 0.0476685f $X=10.425 $Y=0.96 $X2=0 $Y2=0
cc_500 N_Y_c_714_n N_VGND_c_909_n 0.0476685f $X=11.985 $Y=0.96 $X2=0 $Y2=0
cc_501 N_Y_c_714_n N_VGND_c_911_n 0.0472745f $X=11.985 $Y=0.96 $X2=0 $Y2=0
cc_502 N_Y_c_693_n N_VGND_c_913_n 0.0183067f $X=1.065 $Y=0.96 $X2=0 $Y2=0
cc_503 N_Y_c_696_n N_VGND_c_913_n 0.0183067f $X=2.625 $Y=0.96 $X2=0 $Y2=0
cc_504 N_Y_c_699_n N_VGND_c_913_n 0.0183067f $X=4.185 $Y=0.96 $X2=0 $Y2=0
cc_505 N_Y_c_702_n N_VGND_c_913_n 0.0183067f $X=5.745 $Y=0.96 $X2=0 $Y2=0
cc_506 N_Y_c_705_n N_VGND_c_913_n 0.0183067f $X=7.305 $Y=0.96 $X2=0 $Y2=0
cc_507 N_Y_c_708_n N_VGND_c_913_n 0.0183067f $X=8.865 $Y=0.96 $X2=0 $Y2=0
cc_508 N_Y_c_711_n N_VGND_c_913_n 0.0183067f $X=10.425 $Y=0.96 $X2=0 $Y2=0
cc_509 N_Y_c_714_n N_VGND_c_913_n 0.0183067f $X=11.985 $Y=0.96 $X2=0 $Y2=0
