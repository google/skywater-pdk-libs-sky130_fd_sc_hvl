* File: sky130_fd_sc_hvl__sdlclkp_1.spice
* Created: Wed Sep  2 09:10:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__sdlclkp_1.pex.spice"
.subckt sky130_fd_sc_hvl__sdlclkp_1  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_SCE_M1002_g N_A_58_159#_M1002_s N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1281 PD=0.7 PS=1.45 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1018 N_A_58_159#_M1018_d N_GATE_M1018_g N_VGND_M1002_d N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250001
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1008 N_A_495_311#_M1008_d N_A_423_71#_M1008_g N_A_58_159#_M1018_d
+ N_VNB_M1002_b NHV L=0.5 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0
+ M=1 R=0.84 SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1013 N_VGND_M1013_d N_A_423_71#_M1013_g N_A_431_431#_M1013_s N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1004 N_A_423_71#_M1004_d N_CLK_M1004_g N_VGND_M1013_d N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250001
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1005 A_1219_159# N_A_431_431#_M1005_g N_A_495_311#_M1005_s N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1006 N_VGND_M1006_d N_A_1261_133#_M1006_g A_1219_159# N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1000 N_A_1261_133#_M1000_d N_A_495_311#_M1000_g N_VGND_M1006_d N_VNB_M1002_b
+ NHV L=0.5 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1017 A_1783_171# N_A_1261_133#_M1017_g N_A_1630_171#_M1017_s N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=23.0622 NRS=0 M=1 R=0.84
+ SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1010 N_VGND_M1010_d N_CLK_M1010_g A_1783_171# N_VNB_M1002_b NHV L=0.5 W=0.42
+ AD=0.0826538 AS=0.0588 PD=0.782564 PS=0.7 NRD=16.2792 NRS=23.0622 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1001 N_GCLK_M1001_d N_A_1630_171#_M1001_g N_VGND_M1010_d N_VNB_M1002_b NHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.147596 PD=2.03 PS=1.39744 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1011 A_219_457# N_SCE_M1011_g N_VPWR_M1011_s N_VPB_M1011_b PHV L=0.5 W=0.75
+ AD=0.105 AS=0.22875 PD=1.03 PS=2.11 NRD=21.6403 NRS=0 M=1 R=1.5 SA=250000
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1020 N_A_58_159#_M1020_d N_GATE_M1020_g A_219_457# N_VPB_M1011_b PHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=21.6403 M=1 R=1.5 SA=250001
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1019 N_A_495_311#_M1019_d N_A_431_431#_M1019_g N_A_58_159#_M1020_d
+ N_VPB_M1011_b PHV L=0.5 W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0
+ M=1 R=1.5 SA=250002 SB=250000 A=0.375 P=2.5 MULT=1
MM1014 N_VPWR_M1014_d N_A_423_71#_M1014_g N_A_431_431#_M1014_s N_VPB_M1011_b PHV
+ L=0.5 W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1007 N_A_423_71#_M1007_d N_CLK_M1007_g N_VPWR_M1014_d N_VPB_M1011_b PHV L=0.5
+ W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250001
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1015 A_1219_457# N_A_423_71#_M1015_g N_A_495_311#_M1015_s N_VPB_M1011_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1016 N_VPWR_M1016_d N_A_1261_133#_M1016_g A_1219_457# N_VPB_M1011_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1009 N_A_1261_133#_M1009_d N_A_495_311#_M1009_g N_VPWR_M1016_d N_VPB_M1011_b
+ PHV L=0.5 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1003 N_A_1630_171#_M1003_d N_A_1261_133#_M1003_g N_VPWR_M1003_s N_VPB_M1011_b
+ PHV L=0.5 W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250002 A=0.375 P=2.5 MULT=1
MM1021 N_VPWR_M1021_d N_CLK_M1021_g N_A_1630_171#_M1003_d N_VPB_M1011_b PHV
+ L=0.5 W=0.75 AD=0.15125 AS=0.105 PD=1.22667 PS=1.03 NRD=15.2609 NRS=0 M=1
+ R=1.5 SA=250001 SB=250001 A=0.375 P=2.5 MULT=1
MM1012 N_GCLK_M1012_d N_A_1630_171#_M1012_g N_VPWR_M1021_d N_VPB_M1011_b PHV
+ L=0.5 W=1.5 AD=0.3975 AS=0.3025 PD=3.53 PS=2.45333 NRD=0 NRS=0 M=1 R=3
+ SA=250001 SB=250000 A=0.75 P=4 MULT=1
DX22_noxref N_VNB_M1002_b N_VPB_M1011_b NWDIODE A=30.42 P=28.6
*
.include "sky130_fd_sc_hvl__sdlclkp_1.pxi.spice"
*
.ends
*
*
