* NGSPICE file created from sky130_fd_sc_hvl__o21ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_205_443# A1 VPWR VPB phv w=1.5e+06u l=500000u
+  ad=3.15e+11p pd=3.42e+06u as=8.55e+11p ps=7.14e+06u
M1001 Y A2 a_205_443# VPB phv w=1.5e+06u l=500000u
+  ad=4.2e+11p pd=3.56e+06u as=0p ps=0u
M1002 Y B1 a_30_107# VNB nhv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=4.2375e+11p ps=4.13e+06u
M1003 VGND A1 a_30_107# VNB nhv w=750000u l=500000u
+  ad=2.25e+11p pd=2.1e+06u as=0p ps=0u
M1004 a_30_107# A2 VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B1 Y VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends

