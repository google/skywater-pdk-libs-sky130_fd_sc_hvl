* File: sky130_fd_sc_hvl__o21a_1.spice
* Created: Fri Aug 28 09:38:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__o21a_1.pex.spice"
.subckt sky130_fd_sc_hvl__o21a_1  VNB VPB B1 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_83_87#_M1000_g N_X_M1000_s N_VNB_M1000_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.19875 PD=2.07 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1005 N_A_460_107#_M1005_d N_B1_M1005_g N_A_83_87#_M1005_s N_VNB_M1000_b NHV
+ L=0.5 W=0.75 AD=0.105 AS=0.21375 PD=1.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250002 A=0.375 P=2.5 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g N_A_460_107#_M1005_d N_VNB_M1000_b NHV L=0.5
+ W=0.75 AD=0.1125 AS=0.105 PD=1.05 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250001
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1004 N_A_460_107#_M1004_d N_A1_M1004_g N_VGND_M1003_d N_VNB_M1000_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.1125 PD=2.07 PS=1.05 NRD=0 NRS=3.0324 M=1 R=1.5
+ SA=250002 SB=250000 A=0.375 P=2.5 MULT=1
MM1002 N_VPWR_M1002_d N_A_83_87#_M1002_g N_X_M1002_s N_VPB_M1002_b PHV L=0.5
+ W=1.5 AD=0.375 AS=0.4275 PD=2 PS=3.57 NRD=0 NRS=0 M=1 R=3 SA=250000 SB=250003
+ A=0.75 P=4 MULT=1
MM1006 N_A_83_87#_M1006_d N_B1_M1006_g N_VPWR_M1002_d N_VPB_M1002_b PHV L=0.5
+ W=1.5 AD=0.27 AS=0.375 PD=1.86 PS=2 NRD=0 NRS=28.0006 M=1 R=3 SA=250001
+ SB=250002 A=0.75 P=4 MULT=1
MM1001 A_602_443# N_A2_M1001_g N_A_83_87#_M1006_d N_VPB_M1002_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.27 PD=1.78 PS=1.86 NRD=10.8106 NRS=10.1803 M=1 R=3 SA=250002
+ SB=250001 A=0.75 P=4 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g A_602_443# N_VPB_M1002_b PHV L=0.5 W=1.5
+ AD=0.4275 AS=0.21 PD=3.57 PS=1.78 NRD=0 NRS=10.8106 M=1 R=3 SA=250003
+ SB=250000 A=0.75 P=4 MULT=1
DX8_noxref N_VNB_M1000_b N_VPB_M1002_b NWDIODE A=12.948 P=15.16
*
.include "sky130_fd_sc_hvl__o21a_1.pxi.spice"
*
.ends
*
*
