# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__conb_1
  CLASS CORE TIEHIGH ;
  FOREIGN sky130_fd_sc_hvl__conb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.290000 0.430000 0.865000 1.070000 ;
        RECT 0.615000 1.070000 0.865000 1.935000 ;
        RECT 0.615000 1.935000 1.325000 2.185000 ;
        RECT 1.075000 2.185000 1.325000 3.530000 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 0.500000 1.365000 1.500000 ;
        RECT 1.035000 1.500000 1.795000 1.765000 ;
        RECT 1.530000 1.765000 1.795000 3.175000 ;
        RECT 1.530000 3.175000 2.110000 3.815000 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 2.400000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 2.400000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 2.400000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 2.400000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.985000 2.400000 4.155000 ;
      RECT 0.215000  3.175000 0.620000 3.445000 ;
      RECT 0.215000  3.445000 0.865000 3.785000 ;
      RECT 1.535000  0.285000 2.185000 0.625000 ;
      RECT 1.780000  0.625000 2.185000 1.070000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.275000  3.505000 0.445000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.505000 0.805000 3.675000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  0.395000 1.765000 0.565000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.955000  0.395000 2.125000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
  END
END sky130_fd_sc_hvl__conb_1
END LIBRARY
