* File: sky130_fd_sc_hvl__dfxbp_1.pxi.spice
* Created: Fri Aug 28 09:34:35 2020
* 
x_PM_SKY130_FD_SC_HVL__DFXBP_1%VNB N_VNB_M1025_b VNB N_VNB_c_2_p
+ PM_SKY130_FD_SC_HVL__DFXBP_1%VNB
x_PM_SKY130_FD_SC_HVL__DFXBP_1%VPB N_VPB_M1012_b VPB N_VPB_c_101_p
+ PM_SKY130_FD_SC_HVL__DFXBP_1%VPB
x_PM_SKY130_FD_SC_HVL__DFXBP_1%CLK N_CLK_M1025_g N_CLK_M1012_g CLK CLK
+ N_CLK_c_236_n PM_SKY130_FD_SC_HVL__DFXBP_1%CLK
x_PM_SKY130_FD_SC_HVL__DFXBP_1%A_30_112# N_A_30_112#_M1025_s N_A_30_112#_M1012_s
+ N_A_30_112#_M1004_g N_A_30_112#_M1022_g N_A_30_112#_c_266_n
+ N_A_30_112#_M1026_g N_A_30_112#_c_281_n N_A_30_112#_M1011_g
+ N_A_30_112#_M1007_g N_A_30_112#_c_267_n N_A_30_112#_c_269_n
+ N_A_30_112#_c_270_n N_A_30_112#_c_384_p N_A_30_112#_c_334_n
+ N_A_30_112#_c_283_n N_A_30_112#_c_284_n N_A_30_112#_c_287_n
+ N_A_30_112#_c_290_n N_A_30_112#_c_291_n N_A_30_112#_c_292_n
+ N_A_30_112#_c_293_n N_A_30_112#_c_294_n N_A_30_112#_c_297_n
+ N_A_30_112#_c_348_p N_A_30_112#_c_271_n N_A_30_112#_c_301_n
+ N_A_30_112#_c_357_p N_A_30_112#_c_304_n N_A_30_112#_c_305_n
+ N_A_30_112#_c_402_p N_A_30_112#_c_306_n N_A_30_112#_c_309_n
+ N_A_30_112#_c_404_p N_A_30_112#_c_311_n N_A_30_112#_c_272_n
+ N_A_30_112#_c_273_n N_A_30_112#_c_274_n N_A_30_112#_c_275_n
+ N_A_30_112#_c_276_n N_A_30_112#_c_316_n N_A_30_112#_c_424_p
+ N_A_30_112#_c_371_p N_A_30_112#_c_319_n N_A_30_112#_c_322_n
+ N_A_30_112#_M1000_g N_A_30_112#_c_277_n PM_SKY130_FD_SC_HVL__DFXBP_1%A_30_112#
x_PM_SKY130_FD_SC_HVL__DFXBP_1%D N_D_M1013_g N_D_M1006_g N_D_c_517_n N_D_c_521_n
+ D N_D_c_518_n N_D_c_519_n PM_SKY130_FD_SC_HVL__DFXBP_1%D
x_PM_SKY130_FD_SC_HVL__DFXBP_1%A_339_112# N_A_339_112#_M1004_d
+ N_A_339_112#_M1022_d N_A_339_112#_c_558_n N_A_339_112#_M1019_g
+ N_A_339_112#_M1002_g N_A_339_112#_c_559_n N_A_339_112#_c_582_n
+ N_A_339_112#_c_583_n N_A_339_112#_c_560_n N_A_339_112#_c_562_n
+ N_A_339_112#_c_611_n N_A_339_112#_c_563_n N_A_339_112#_c_565_n
+ N_A_339_112#_c_567_n N_A_339_112#_c_637_p N_A_339_112#_c_568_n
+ N_A_339_112#_c_570_n N_A_339_112#_c_642_p N_A_339_112#_c_613_n
+ N_A_339_112#_c_572_n N_A_339_112#_c_573_n N_A_339_112#_c_622_n
+ N_A_339_112#_c_623_n N_A_339_112#_c_624_n N_A_339_112#_M1018_g
+ N_A_339_112#_M1024_g PM_SKY130_FD_SC_HVL__DFXBP_1%A_339_112#
x_PM_SKY130_FD_SC_HVL__DFXBP_1%A_1063_85# N_A_1063_85#_M1023_d
+ N_A_1063_85#_M1017_d N_A_1063_85#_c_729_n N_A_1063_85#_c_725_n
+ N_A_1063_85#_c_726_n N_A_1063_85#_c_727_n N_A_1063_85#_c_731_n
+ N_A_1063_85#_c_744_n N_A_1063_85#_c_732_n N_A_1063_85#_M1021_g
+ N_A_1063_85#_M1015_g PM_SKY130_FD_SC_HVL__DFXBP_1%A_1063_85#
x_PM_SKY130_FD_SC_HVL__DFXBP_1%A_865_111# N_A_865_111#_M1026_d
+ N_A_865_111#_M1019_d N_A_865_111#_c_786_n N_A_865_111#_c_790_n
+ N_A_865_111#_c_791_n N_A_865_111#_c_787_n N_A_865_111#_c_792_n
+ N_A_865_111#_c_829_n N_A_865_111#_M1023_g N_A_865_111#_M1017_g
+ PM_SKY130_FD_SC_HVL__DFXBP_1%A_865_111#
x_PM_SKY130_FD_SC_HVL__DFXBP_1%A_1711_85# N_A_1711_85#_M1009_d
+ N_A_1711_85#_M1003_d N_A_1711_85#_M1016_g N_A_1711_85#_M1008_g
+ N_A_1711_85#_M1010_g N_A_1711_85#_M1001_g N_A_1711_85#_c_860_n
+ N_A_1711_85#_M1005_g N_A_1711_85#_M1014_g N_A_1711_85#_c_862_n
+ N_A_1711_85#_c_863_n N_A_1711_85#_c_864_n N_A_1711_85#_c_865_n
+ N_A_1711_85#_c_866_n N_A_1711_85#_c_879_n N_A_1711_85#_c_893_p
+ N_A_1711_85#_c_868_n N_A_1711_85#_c_869_n
+ PM_SKY130_FD_SC_HVL__DFXBP_1%A_1711_85#
x_PM_SKY130_FD_SC_HVL__DFXBP_1%A_1494_539# N_A_1494_539#_M1024_d
+ N_A_1494_539#_M1000_d N_A_1494_539#_M1009_g N_A_1494_539#_M1003_g
+ N_A_1494_539#_c_990_n N_A_1494_539#_c_1013_n N_A_1494_539#_c_979_n
+ N_A_1494_539#_c_981_n N_A_1494_539#_c_983_n N_A_1494_539#_c_992_n
+ N_A_1494_539#_c_993_n N_A_1494_539#_c_1047_n N_A_1494_539#_c_984_n
+ N_A_1494_539#_c_995_n N_A_1494_539#_c_985_n N_A_1494_539#_c_986_n
+ PM_SKY130_FD_SC_HVL__DFXBP_1%A_1494_539#
x_PM_SKY130_FD_SC_HVL__DFXBP_1%A_2365_443# N_A_2365_443#_M1014_s
+ N_A_2365_443#_M1005_s N_A_2365_443#_M1020_g N_A_2365_443#_M1027_g
+ N_A_2365_443#_c_1084_n N_A_2365_443#_c_1078_n N_A_2365_443#_c_1079_n
+ N_A_2365_443#_c_1080_n N_A_2365_443#_c_1087_n N_A_2365_443#_c_1103_n
+ PM_SKY130_FD_SC_HVL__DFXBP_1%A_2365_443#
x_PM_SKY130_FD_SC_HVL__DFXBP_1%VPWR N_VPWR_M1012_d N_VPWR_M1006_s N_VPWR_M1015_d
+ N_VPWR_M1008_d N_VPWR_M1001_d N_VPWR_M1005_d VPWR N_VPWR_c_1125_n
+ N_VPWR_c_1128_n N_VPWR_c_1131_n N_VPWR_c_1134_n N_VPWR_c_1137_n
+ N_VPWR_c_1140_n N_VPWR_c_1143_n PM_SKY130_FD_SC_HVL__DFXBP_1%VPWR
x_PM_SKY130_FD_SC_HVL__DFXBP_1%A_709_111# N_A_709_111#_M1013_d
+ N_A_709_111#_M1006_d N_A_709_111#_c_1224_n N_A_709_111#_c_1225_n
+ N_A_709_111#_c_1229_n N_A_709_111#_c_1223_n
+ PM_SKY130_FD_SC_HVL__DFXBP_1%A_709_111#
x_PM_SKY130_FD_SC_HVL__DFXBP_1%Q N_Q_M1010_s N_Q_M1001_s Q Q Q Q Q Q Q
+ N_Q_c_1256_n Q N_Q_c_1262_n Q PM_SKY130_FD_SC_HVL__DFXBP_1%Q
x_PM_SKY130_FD_SC_HVL__DFXBP_1%Q_N N_Q_N_M1027_d N_Q_N_M1020_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N Q_N PM_SKY130_FD_SC_HVL__DFXBP_1%Q_N
x_PM_SKY130_FD_SC_HVL__DFXBP_1%VGND N_VGND_M1025_d N_VGND_M1013_s N_VGND_M1021_d
+ N_VGND_M1016_d N_VGND_M1010_d N_VGND_M1014_d VGND N_VGND_c_1302_n
+ N_VGND_c_1304_n N_VGND_c_1306_n N_VGND_c_1308_n N_VGND_c_1310_n
+ N_VGND_c_1312_n N_VGND_c_1314_n PM_SKY130_FD_SC_HVL__DFXBP_1%VGND
cc_1 N_VNB_M1025_b N_CLK_M1025_g 0.0874785f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=0.77
cc_2 N_VNB_c_2_p N_CLK_M1025_g 9.31318e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=0.77
cc_3 N_VNB_M1025_b N_CLK_c_236_n 0.0353715f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=1.715
cc_4 N_VNB_M1025_b N_A_30_112#_M1004_g 0.0446898f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.58
cc_5 N_VNB_c_2_p N_A_30_112#_M1004_g 5.69641e-19 $X=0.24 $Y=0 $X2=0.635 $Y2=1.58
cc_6 N_VNB_M1025_b N_A_30_112#_c_266_n 0.110108f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=1.715
cc_7 N_VNB_M1025_b N_A_30_112#_c_267_n 0.0344242f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_8 N_VNB_c_2_p N_A_30_112#_c_267_n 7.73497e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_9 N_VNB_M1025_b N_A_30_112#_c_269_n 0.0265284f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_10 N_VNB_M1025_b N_A_30_112#_c_270_n 0.0115986f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1025_b N_A_30_112#_c_271_n 0.00138672f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1025_b N_A_30_112#_c_272_n 0.00286616f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1025_b N_A_30_112#_c_273_n 0.0421975f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_M1025_b N_A_30_112#_c_274_n 0.0091351f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_15 N_VNB_M1025_b N_A_30_112#_c_275_n 0.0762164f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_16 N_VNB_M1025_b N_A_30_112#_c_276_n 8.06181e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_17 N_VNB_M1025_b N_A_30_112#_c_277_n 0.0440429f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_c_2_p N_A_30_112#_c_277_n 0.00227358f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_19 N_VNB_M1025_b N_D_M1013_g 0.0465542f $X=-0.33 $Y=-0.265 $X2=0.665 $Y2=0.77
cc_20 N_VNB_c_2_p N_D_M1013_g 5.84397e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=0.77
cc_21 N_VNB_M1025_b N_D_c_517_n 0.0307406f $X=-0.33 $Y=-0.265 $X2=0.635 $Y2=1.58
cc_22 N_VNB_M1025_b N_D_c_518_n 0.0550216f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=1.665
cc_23 N_VNB_M1025_b N_D_c_519_n 0.0137238f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_24 N_VNB_M1025_b N_A_339_112#_c_558_n 0.0361874f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.815
cc_25 N_VNB_M1025_b N_A_339_112#_c_559_n 0.0528328f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_26 N_VNB_M1025_b N_A_339_112#_c_560_n 0.0157449f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_27 N_VNB_c_2_p N_A_339_112#_c_560_n 3.80008e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_28 N_VNB_M1025_b N_A_339_112#_c_562_n 0.040699f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_29 N_VNB_M1025_b N_A_339_112#_c_563_n 0.117555f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_30 N_VNB_c_2_p N_A_339_112#_c_563_n 0.00552846f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_31 N_VNB_M1025_b N_A_339_112#_c_565_n 0.013621f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_32 N_VNB_c_2_p N_A_339_112#_c_565_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_33 N_VNB_M1025_b N_A_339_112#_c_567_n 0.013451f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_M1025_b N_A_339_112#_c_568_n 0.0640612f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_35 N_VNB_c_2_p N_A_339_112#_c_568_n 0.00289338f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_36 N_VNB_M1025_b N_A_339_112#_c_570_n 0.0136293f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_37 N_VNB_c_2_p N_A_339_112#_c_570_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_38 N_VNB_M1025_b N_A_339_112#_c_572_n 0.0183611f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_39 N_VNB_M1025_b N_A_339_112#_c_573_n 0.00267798f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_M1025_b N_A_339_112#_M1018_g 0.089141f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_41 N_VNB_c_2_p N_A_339_112#_M1018_g 5.84397e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_42 N_VNB_M1025_b N_A_339_112#_M1024_g 0.0981681f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_c_2_p N_A_339_112#_M1024_g 0.00101638f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_44 N_VNB_M1025_b N_A_1063_85#_c_725_n 0.00136456f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_45 N_VNB_M1025_b N_A_1063_85#_c_726_n 0.00677277f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=1.715
cc_46 N_VNB_M1025_b N_A_1063_85#_c_727_n 0.0105307f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=1.715
cc_47 N_VNB_M1025_b N_A_1063_85#_M1021_g 0.108324f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_M1025_b N_A_865_111#_c_786_n 0.00712802f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_49 N_VNB_M1025_b N_A_865_111#_c_787_n 0.00215102f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=1.53
cc_50 N_VNB_M1025_b N_A_865_111#_M1023_g 0.0872879f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_51 N_VNB_c_2_p N_A_865_111#_M1023_g 5.84397e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_52 N_VNB_M1025_b N_A_1711_85#_M1016_g 0.0724861f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.58
cc_53 N_VNB_c_2_p N_A_1711_85#_M1016_g 0.00100492f $X=0.24 $Y=0 $X2=0.635
+ $Y2=1.58
cc_54 N_VNB_M1025_b N_A_1711_85#_M1010_g 0.0505647f $X=-0.33 $Y=-0.265 $X2=0.675
+ $Y2=2.31
cc_55 N_VNB_c_2_p N_A_1711_85#_M1010_g 0.00121146f $X=0.24 $Y=0 $X2=0.675
+ $Y2=2.31
cc_56 N_VNB_M1025_b N_A_1711_85#_c_860_n 0.0497326f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_57 N_VNB_M1025_b N_A_1711_85#_M1014_g 0.0429716f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_58 N_VNB_M1025_b N_A_1711_85#_c_862_n 0.0450201f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_59 N_VNB_M1025_b N_A_1711_85#_c_863_n 0.01645f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_60 N_VNB_M1025_b N_A_1711_85#_c_864_n 0.0225559f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_61 N_VNB_M1025_b N_A_1711_85#_c_865_n 0.00738444f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_62 N_VNB_M1025_b N_A_1711_85#_c_866_n 0.0206553f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_63 N_VNB_c_2_p N_A_1711_85#_c_866_n 7.78491e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_64 N_VNB_M1025_b N_A_1711_85#_c_868_n 0.0424423f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_65 N_VNB_M1025_b N_A_1711_85#_c_869_n 7.96456e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_66 N_VNB_M1025_b N_A_1494_539#_M1009_g 0.0818995f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=1.58
cc_67 N_VNB_c_2_p N_A_1494_539#_M1009_g 9.36715e-19 $X=0.24 $Y=0 $X2=0.635
+ $Y2=1.58
cc_68 N_VNB_M1025_b N_A_1494_539#_c_979_n 0.0206539f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_69 N_VNB_c_2_p N_A_1494_539#_c_979_n 0.00268535f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_70 N_VNB_M1025_b N_A_1494_539#_c_981_n 0.00829488f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_71 N_VNB_c_2_p N_A_1494_539#_c_981_n 6.31888e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_72 N_VNB_M1025_b N_A_1494_539#_c_983_n 0.00644207f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_73 N_VNB_M1025_b N_A_1494_539#_c_984_n 0.00716132f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_74 N_VNB_M1025_b N_A_1494_539#_c_985_n 0.0108774f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_75 N_VNB_M1025_b N_A_1494_539#_c_986_n 0.00139559f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_76 N_VNB_M1025_b N_A_2365_443#_M1027_g 0.0496474f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=1.715
cc_77 N_VNB_c_2_p N_A_2365_443#_M1027_g 9.38781e-19 $X=0.24 $Y=0 $X2=0.675
+ $Y2=1.715
cc_78 N_VNB_M1025_b N_A_2365_443#_c_1078_n 0.0105503f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=2.035
cc_79 N_VNB_M1025_b N_A_2365_443#_c_1079_n 0.00321504f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_80 N_VNB_M1025_b N_A_2365_443#_c_1080_n 0.0339026f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_81 N_VNB_M1025_b N_A_709_111#_c_1223_n 0.00611033f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=2.31
cc_82 N_VNB_M1025_b Q 8.282e-19 $X=-0.33 $Y=-0.265 $X2=0.635 $Y2=1.58
cc_83 N_VNB_M1025_b N_Q_c_1256_n 0.0149895f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_84 N_VNB_M1025_b Q 0.00433696f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_85 N_VNB_M1025_b Q_N 0.0564553f $X=-0.33 $Y=-0.265 $X2=0.685 $Y2=2.815
cc_86 N_VNB_M1025_b N_VGND_c_1302_n 0.0499581f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_87 N_VNB_c_2_p N_VGND_c_1302_n 0.00269208f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_88 N_VNB_M1025_b N_VGND_c_1304_n 0.0734131f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_89 N_VNB_c_2_p N_VGND_c_1304_n 0.002522f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_90 N_VNB_M1025_b N_VGND_c_1306_n 0.0512348f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_91 N_VNB_c_2_p N_VGND_c_1306_n 0.00269097f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_92 N_VNB_M1025_b N_VGND_c_1308_n 0.0508811f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_93 N_VNB_c_2_p N_VGND_c_1308_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_94 N_VNB_M1025_b N_VGND_c_1310_n 0.0602757f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_95 N_VNB_c_2_p N_VGND_c_1310_n 0.00156945f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_96 N_VNB_M1025_b N_VGND_c_1312_n 0.0734054f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_97 N_VNB_c_2_p N_VGND_c_1312_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_98 N_VNB_M1025_b N_VGND_c_1314_n 0.201857f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_99 N_VNB_c_2_p N_VGND_c_1314_n 1.48807f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_100 N_VPB_M1012_b N_CLK_M1012_g 0.041921f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.815
cc_101 N_VPB_c_101_p N_CLK_M1012_g 0.00365752f $X=13.68 $Y=4.07 $X2=0.685
+ $Y2=2.815
cc_102 N_VPB_M1012_b N_CLK_c_236_n 0.0431928f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=1.715
cc_103 N_VPB_M1012_b N_A_30_112#_M1022_g 0.0810772f $X=-0.33 $Y=1.885 $X2=0.675
+ $Y2=1.715
cc_104 N_VPB_c_101_p N_A_30_112#_M1022_g 0.0032569f $X=13.68 $Y=4.07 $X2=0.675
+ $Y2=1.715
cc_105 N_VPB_M1012_b N_A_30_112#_c_281_n 0.0763066f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=1.665
cc_106 N_VPB_M1012_b N_A_30_112#_c_269_n 0.0637276f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_107 N_VPB_M1012_b N_A_30_112#_c_283_n 0.00210798f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_108 N_VPB_M1012_b N_A_30_112#_c_284_n 0.020517f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_109 VPB N_A_30_112#_c_284_n 0.00187532f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_110 N_VPB_c_101_p N_A_30_112#_c_284_n 0.0217805f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_111 N_VPB_M1012_b N_A_30_112#_c_287_n 0.00250055f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_112 VPB N_A_30_112#_c_287_n 4.01254e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_113 N_VPB_c_101_p N_A_30_112#_c_287_n 0.00485128f $X=13.68 $Y=4.07 $X2=0
+ $Y2=0
cc_114 N_VPB_M1012_b N_A_30_112#_c_290_n 0.0264006f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_115 N_VPB_M1012_b N_A_30_112#_c_291_n 0.0290225f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_116 N_VPB_M1012_b N_A_30_112#_c_292_n 0.00919848f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_117 N_VPB_M1012_b N_A_30_112#_c_293_n 0.00209454f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_118 N_VPB_M1012_b N_A_30_112#_c_294_n 0.0140415f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_119 VPB N_A_30_112#_c_294_n 0.00130714f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_120 N_VPB_c_101_p N_A_30_112#_c_294_n 0.0133181f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_121 N_VPB_M1012_b N_A_30_112#_c_297_n 0.00308907f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_122 VPB N_A_30_112#_c_297_n 3.61175e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_123 N_VPB_c_101_p N_A_30_112#_c_297_n 0.00388086f $X=13.68 $Y=4.07 $X2=0
+ $Y2=0
cc_124 N_VPB_M1012_b N_A_30_112#_c_271_n 0.00410851f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_125 N_VPB_M1012_b N_A_30_112#_c_301_n 0.019616f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_126 VPB N_A_30_112#_c_301_n 0.00208457f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_127 N_VPB_c_101_p N_A_30_112#_c_301_n 0.0216298f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_128 N_VPB_M1012_b N_A_30_112#_c_304_n 0.00214923f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_129 N_VPB_M1012_b N_A_30_112#_c_305_n 0.00676553f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_130 N_VPB_M1012_b N_A_30_112#_c_306_n 0.00100701f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_131 VPB N_A_30_112#_c_306_n 0.00203434f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_132 N_VPB_c_101_p N_A_30_112#_c_306_n 0.03408f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_133 VPB N_A_30_112#_c_309_n 8.21022e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_134 N_VPB_c_101_p N_A_30_112#_c_309_n 0.0108189f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_135 N_VPB_M1012_b N_A_30_112#_c_311_n 0.0103797f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_136 VPB N_A_30_112#_c_311_n 0.00350141f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_137 N_VPB_c_101_p N_A_30_112#_c_311_n 0.0643075f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_138 N_VPB_M1012_b N_A_30_112#_c_272_n 0.00898533f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_139 N_VPB_M1012_b N_A_30_112#_c_275_n 0.00159637f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_140 N_VPB_M1012_b N_A_30_112#_c_316_n 0.00180427f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_141 VPB N_A_30_112#_c_316_n 3.61175e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_142 N_VPB_c_101_p N_A_30_112#_c_316_n 0.00388086f $X=13.68 $Y=4.07 $X2=0
+ $Y2=0
cc_143 N_VPB_M1012_b N_A_30_112#_c_319_n 0.0859255f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_144 VPB N_A_30_112#_c_319_n 0.00957431f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_145 N_VPB_c_101_p N_A_30_112#_c_319_n 0.0131476f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_146 VPB N_A_30_112#_c_322_n 8.21022e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_147 N_VPB_c_101_p N_A_30_112#_c_322_n 0.0108189f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_148 N_VPB_M1012_b N_D_M1006_g 0.0822763f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.815
cc_149 N_VPB_M1012_b N_D_c_521_n 0.0311014f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_150 N_VPB_M1012_b N_D_c_518_n 0.00367852f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=1.665
cc_151 N_VPB_M1012_b N_D_c_519_n 0.0110064f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_152 N_VPB_M1012_b N_A_339_112#_c_558_n 0.0611067f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.815
cc_153 N_VPB_M1012_b N_A_339_112#_M1019_g 0.0698011f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_154 N_VPB_M1012_b N_A_339_112#_M1002_g 0.0395284f $X=-0.33 $Y=1.885 $X2=0.675
+ $Y2=1.715
cc_155 N_VPB_M1012_b N_A_339_112#_c_559_n 0.0929467f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_156 N_VPB_M1012_b N_A_339_112#_c_582_n 0.00186698f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=2.035
cc_157 N_VPB_M1012_b N_A_339_112#_c_583_n 0.00221638f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_158 N_VPB_M1012_b N_A_339_112#_c_572_n 0.0168755f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_159 N_VPB_M1012_b N_A_1063_85#_c_729_n 0.011026f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.815
cc_160 N_VPB_M1012_b N_A_1063_85#_c_727_n 0.0133535f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=1.715
cc_161 N_VPB_M1012_b N_A_1063_85#_c_731_n 0.00403608f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=2.31
cc_162 N_VPB_M1012_b N_A_1063_85#_c_732_n 0.00130462f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_163 N_VPB_M1012_b N_A_1063_85#_M1021_g 0.10214f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_164 N_VPB_M1012_b N_A_865_111#_c_790_n 0.0106031f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_165 N_VPB_M1012_b N_A_865_111#_c_791_n 0.0210532f $X=-0.33 $Y=1.885 $X2=0.675
+ $Y2=1.715
cc_166 N_VPB_M1012_b N_A_865_111#_c_792_n 8.61801e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_167 N_VPB_M1012_b N_A_865_111#_M1023_g 0.101318f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_168 VPB N_A_865_111#_M1023_g 0.00957431f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_169 N_VPB_c_101_p N_A_865_111#_M1023_g 0.0153316f $X=13.68 $Y=4.07 $X2=0
+ $Y2=0
cc_170 N_VPB_M1012_b N_A_1711_85#_M1008_g 0.0681845f $X=-0.33 $Y=1.885 $X2=0.675
+ $Y2=1.715
cc_171 N_VPB_M1012_b N_A_1711_85#_M1001_g 0.0440283f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=2.035
cc_172 VPB N_A_1711_85#_M1001_g 0.00970178f $X=0 $Y=3.955 $X2=0.725 $Y2=2.035
cc_173 N_VPB_c_101_p N_A_1711_85#_M1001_g 0.0159423f $X=13.68 $Y=4.07 $X2=0.725
+ $Y2=2.035
cc_174 N_VPB_M1012_b N_A_1711_85#_c_860_n 0.0395208f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_175 N_VPB_M1012_b N_A_1711_85#_M1005_g 0.0430607f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_176 N_VPB_M1012_b N_A_1711_85#_c_862_n 0.0367864f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_177 N_VPB_M1012_b N_A_1711_85#_c_863_n 0.0106129f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_178 N_VPB_M1012_b N_A_1711_85#_c_864_n 0.015276f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_179 N_VPB_M1012_b N_A_1711_85#_c_879_n 0.0175381f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_180 VPB N_A_1711_85#_c_879_n 9.90209e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_181 N_VPB_c_101_p N_A_1711_85#_c_879_n 0.0146337f $X=13.68 $Y=4.07 $X2=0
+ $Y2=0
cc_182 N_VPB_M1012_b N_A_1711_85#_c_868_n 0.0282485f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_183 N_VPB_M1012_b N_A_1494_539#_M1003_g 0.0422146f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=1.715
cc_184 VPB N_A_1494_539#_M1003_g 0.00957431f $X=0 $Y=3.955 $X2=0.675 $Y2=1.715
cc_185 N_VPB_c_101_p N_A_1494_539#_M1003_g 0.0186208f $X=13.68 $Y=4.07 $X2=0.675
+ $Y2=1.715
cc_186 N_VPB_M1012_b N_A_1494_539#_c_990_n 0.00365543f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=2.31
cc_187 N_VPB_M1012_b N_A_1494_539#_c_983_n 0.00260295f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_188 N_VPB_M1012_b N_A_1494_539#_c_992_n 0.0076152f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_189 N_VPB_M1012_b N_A_1494_539#_c_993_n 0.00475525f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_190 N_VPB_M1012_b N_A_1494_539#_c_984_n 0.0699515f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_191 N_VPB_M1012_b N_A_1494_539#_c_995_n 0.00300391f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_192 N_VPB_M1012_b N_A_1494_539#_c_985_n 0.0177673f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_193 N_VPB_M1012_b N_A_2365_443#_M1020_g 0.04251f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_194 VPB N_A_2365_443#_M1020_g 0.00970178f $X=0 $Y=3.955 $X2=0.635 $Y2=1.58
cc_195 N_VPB_c_101_p N_A_2365_443#_M1020_g 0.0162989f $X=13.68 $Y=4.07 $X2=0.635
+ $Y2=1.58
cc_196 N_VPB_M1012_b N_A_2365_443#_c_1084_n 0.0126545f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=2.31
cc_197 N_VPB_M1012_b N_A_2365_443#_c_1079_n 0.00321504f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_198 N_VPB_M1012_b N_A_2365_443#_c_1080_n 0.0226342f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_199 N_VPB_M1012_b N_A_2365_443#_c_1087_n 0.00156688f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_200 N_VPB_M1012_b N_VPWR_c_1125_n 0.0299117f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1125_n 0.00166879f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_202 N_VPB_c_101_p N_VPWR_c_1125_n 0.0254284f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_203 N_VPB_M1012_b N_VPWR_c_1128_n 0.0399828f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1128_n 0.0014985f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_205 N_VPB_c_101_p N_VPWR_c_1128_n 0.0228337f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_206 N_VPB_M1012_b N_VPWR_c_1131_n 0.0174832f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1131_n 0.00278037f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_208 N_VPB_c_101_p N_VPWR_c_1131_n 0.0423987f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_209 N_VPB_M1012_b N_VPWR_c_1134_n 0.0201614f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1134_n 0.00277683f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_211 N_VPB_c_101_p N_VPWR_c_1134_n 0.0424752f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_212 N_VPB_M1012_b N_VPWR_c_1137_n 0.0377499f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1137_n 0.00192587f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_214 N_VPB_c_101_p N_VPWR_c_1137_n 0.0251442f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_215 N_VPB_M1012_b N_VPWR_c_1140_n 0.0323138f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1140_n 0.00335473f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_217 N_VPB_c_101_p N_VPWR_c_1140_n 0.0490696f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_218 N_VPB_M1012_b N_VPWR_c_1143_n 0.165787f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1143_n 1.48432f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_220 N_VPB_c_101_p N_VPWR_c_1143_n 0.0660327f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_221 N_VPB_M1012_b N_A_709_111#_c_1224_n 0.00300301f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=1.58
cc_222 N_VPB_M1012_b N_A_709_111#_c_1225_n 0.00212457f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_223 N_VPB_M1012_b N_A_709_111#_c_1223_n 0.00535647f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=2.31
cc_224 N_VPB_M1012_b Q 8.29097e-19 $X=-0.33 $Y=1.885 $X2=0.635 $Y2=1.58
cc_225 N_VPB_M1012_b Q 0.0131234f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_226 VPB Q 0.00152012f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_227 N_VPB_c_101_p Q 0.020524f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_228 N_VPB_M1012_b N_Q_c_1262_n 0.00435692f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_229 N_VPB_M1012_b Q_N 0.0120961f $X=-0.33 $Y=1.885 $X2=0.685 $Y2=2.815
cc_230 N_VPB_M1012_b Q_N 0.00694735f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_231 N_VPB_M1012_b Q_N 0.0486863f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_232 VPB Q_N 0.00110823f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_233 N_VPB_c_101_p Q_N 0.0182942f $X=13.68 $Y=4.07 $X2=0 $Y2=0
cc_234 N_CLK_M1025_g N_A_30_112#_M1004_g 0.03642f $X=0.665 $Y=0.77 $X2=0 $Y2=0
cc_235 CLK N_A_30_112#_M1022_g 0.0013606f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_236 N_CLK_c_236_n N_A_30_112#_M1022_g 0.0378138f $X=0.725 $Y=1.715 $X2=0
+ $Y2=0
cc_237 N_CLK_M1025_g N_A_30_112#_c_267_n 0.0215326f $X=0.665 $Y=0.77 $X2=0 $Y2=0
cc_238 N_CLK_M1025_g N_A_30_112#_c_269_n 0.0326698f $X=0.665 $Y=0.77 $X2=0 $Y2=0
cc_239 N_CLK_M1012_g N_A_30_112#_c_269_n 0.00926821f $X=0.685 $Y=2.815 $X2=0
+ $Y2=0
cc_240 CLK N_A_30_112#_c_269_n 0.0499846f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_241 N_CLK_M1025_g N_A_30_112#_c_270_n 0.0289405f $X=0.665 $Y=0.77 $X2=0 $Y2=0
cc_242 CLK N_A_30_112#_c_270_n 0.0238298f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_243 N_CLK_c_236_n N_A_30_112#_c_270_n 8.3915e-19 $X=0.725 $Y=1.715 $X2=0
+ $Y2=0
cc_244 N_CLK_M1025_g N_A_30_112#_c_334_n 0.00108574f $X=0.665 $Y=0.77 $X2=0
+ $Y2=0
cc_245 CLK N_A_30_112#_c_334_n 0.0142697f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_246 N_CLK_c_236_n N_A_30_112#_c_334_n 0.00144974f $X=0.725 $Y=1.715 $X2=0
+ $Y2=0
cc_247 N_CLK_M1012_g N_A_30_112#_c_283_n 4.02551e-19 $X=0.685 $Y=2.815 $X2=0
+ $Y2=0
cc_248 CLK N_A_30_112#_c_283_n 0.0113249f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_249 N_CLK_c_236_n N_A_30_112#_c_283_n 0.00225003f $X=0.725 $Y=1.715 $X2=0
+ $Y2=0
cc_250 N_CLK_M1025_g N_A_30_112#_c_274_n 0.00513266f $X=0.665 $Y=0.77 $X2=0
+ $Y2=0
cc_251 CLK N_A_30_112#_c_275_n 0.0013278f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_252 N_CLK_c_236_n N_A_30_112#_c_275_n 0.0185399f $X=0.725 $Y=1.715 $X2=0
+ $Y2=0
cc_253 N_CLK_M1012_g N_VPWR_c_1125_n 0.0605327f $X=0.685 $Y=2.815 $X2=0 $Y2=0
cc_254 CLK N_VPWR_c_1125_n 0.0256698f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_255 N_CLK_M1012_g N_VPWR_c_1143_n 0.00440303f $X=0.685 $Y=2.815 $X2=0 $Y2=0
cc_256 N_CLK_M1025_g N_VGND_c_1302_n 0.0364365f $X=0.665 $Y=0.77 $X2=0 $Y2=0
cc_257 N_CLK_M1025_g N_VGND_c_1314_n 0.00662845f $X=0.665 $Y=0.77 $X2=0 $Y2=0
cc_258 N_A_30_112#_c_266_n N_D_M1013_g 0.0574353f $X=4.075 $Y=1.085 $X2=0 $Y2=0
cc_259 N_A_30_112#_c_291_n N_D_M1006_g 0.0217824f $X=3.18 $Y=2.39 $X2=0 $Y2=0
cc_260 N_A_30_112#_c_293_n N_D_M1006_g 0.0382915f $X=3.265 $Y=3.335 $X2=0 $Y2=0
cc_261 N_A_30_112#_c_294_n N_D_M1006_g 0.00858364f $X=3.95 $Y=3.42 $X2=0 $Y2=0
cc_262 N_A_30_112#_c_271_n N_D_M1006_g 3.35339e-19 $X=4.035 $Y=3.335 $X2=0 $Y2=0
cc_263 N_A_30_112#_c_348_p N_D_c_517_n 2.59988e-19 $X=3.965 $Y=1.28 $X2=0 $Y2=0
cc_264 N_A_30_112#_c_291_n N_D_c_521_n 0.00127067f $X=3.18 $Y=2.39 $X2=0 $Y2=0
cc_265 N_A_30_112#_c_271_n N_D_c_521_n 7.63678e-19 $X=4.035 $Y=3.335 $X2=0 $Y2=0
cc_266 N_A_30_112#_c_271_n N_D_c_518_n 9.81101e-19 $X=4.035 $Y=3.335 $X2=0 $Y2=0
cc_267 N_A_30_112#_c_276_n N_D_c_518_n 2.59988e-19 $X=4 $Y=1.785 $X2=0 $Y2=0
cc_268 N_A_30_112#_c_291_n N_D_c_519_n 0.0643689f $X=3.18 $Y=2.39 $X2=0 $Y2=0
cc_269 N_A_30_112#_c_266_n N_A_339_112#_c_558_n 0.0363646f $X=4.075 $Y=1.085
+ $X2=0 $Y2=0
cc_270 N_A_30_112#_c_281_n N_A_339_112#_c_558_n 0.0274836f $X=4.855 $Y=2.645
+ $X2=0 $Y2=0
cc_271 N_A_30_112#_c_271_n N_A_339_112#_c_558_n 0.0103931f $X=4.035 $Y=3.335
+ $X2=0 $Y2=0
cc_272 N_A_30_112#_c_357_p N_A_339_112#_c_558_n 3.18044e-19 $X=4.92 $Y=2.37
+ $X2=0 $Y2=0
cc_273 N_A_30_112#_c_276_n N_A_339_112#_c_558_n 5.26688e-19 $X=4 $Y=1.785 $X2=0
+ $Y2=0
cc_274 N_A_30_112#_c_281_n N_A_339_112#_M1019_g 0.025122f $X=4.855 $Y=2.645
+ $X2=0 $Y2=0
cc_275 N_A_30_112#_c_293_n N_A_339_112#_M1019_g 4.65037e-19 $X=3.265 $Y=3.335
+ $X2=0 $Y2=0
cc_276 N_A_30_112#_c_294_n N_A_339_112#_M1019_g 0.00564101f $X=3.95 $Y=3.42
+ $X2=0 $Y2=0
cc_277 N_A_30_112#_c_271_n N_A_339_112#_M1019_g 0.0449057f $X=4.035 $Y=3.335
+ $X2=0 $Y2=0
cc_278 N_A_30_112#_c_301_n N_A_339_112#_M1019_g 0.00887434f $X=4.755 $Y=3.42
+ $X2=0 $Y2=0
cc_279 N_A_30_112#_c_357_p N_A_339_112#_M1019_g 3.0317e-19 $X=4.92 $Y=2.37 $X2=0
+ $Y2=0
cc_280 N_A_30_112#_c_304_n N_A_339_112#_M1019_g 4.54326e-19 $X=4.92 $Y=3.335
+ $X2=0 $Y2=0
cc_281 N_A_30_112#_c_311_n N_A_339_112#_M1002_g 0.00368291f $X=7.975 $Y=3.72
+ $X2=0 $Y2=0
cc_282 N_A_30_112#_c_272_n N_A_339_112#_M1002_g 0.0358196f $X=8.11 $Y=1.27 $X2=0
+ $Y2=0
cc_283 N_A_30_112#_c_319_n N_A_339_112#_M1002_g 0.0132295f $X=7.26 $Y=2.37 $X2=0
+ $Y2=0
cc_284 N_A_30_112#_c_272_n N_A_339_112#_c_559_n 0.0420127f $X=8.11 $Y=1.27 $X2=0
+ $Y2=0
cc_285 N_A_30_112#_c_273_n N_A_339_112#_c_559_n 0.0379051f $X=8.11 $Y=1.27 $X2=0
+ $Y2=0
cc_286 N_A_30_112#_c_371_p N_A_339_112#_c_559_n 0.00163564f $X=7.26 $Y=2.37
+ $X2=0 $Y2=0
cc_287 N_A_30_112#_c_319_n N_A_339_112#_c_559_n 0.0417054f $X=7.26 $Y=2.37 $X2=0
+ $Y2=0
cc_288 N_A_30_112#_M1022_g N_A_339_112#_c_582_n 0.00404718f $X=1.465 $Y=2.815
+ $X2=6.96 $Y2=0
cc_289 N_A_30_112#_c_283_n N_A_339_112#_c_582_n 0.0553435f $X=1.425 $Y=3.41
+ $X2=6.96 $Y2=0
cc_290 N_A_30_112#_c_290_n N_A_339_112#_c_582_n 0.0551288f $X=2.205 $Y=3.41
+ $X2=6.96 $Y2=0
cc_291 N_A_30_112#_M1022_g N_A_339_112#_c_583_n 0.0146186f $X=1.465 $Y=2.815
+ $X2=6.96 $Y2=0.057
cc_292 N_A_30_112#_c_284_n N_A_339_112#_c_583_n 0.0179369f $X=2.12 $Y=3.495
+ $X2=6.96 $Y2=0.057
cc_293 N_A_30_112#_M1004_g N_A_339_112#_c_560_n 0.00674345f $X=1.445 $Y=0.77
+ $X2=0 $Y2=0
cc_294 N_A_30_112#_c_275_n N_A_339_112#_c_560_n 0.00389821f $X=1.38 $Y=1.365
+ $X2=0 $Y2=0
cc_295 N_A_30_112#_c_266_n N_A_339_112#_c_611_n 0.0011153f $X=4.075 $Y=1.085
+ $X2=0 $Y2=0
cc_296 N_A_30_112#_c_266_n N_A_339_112#_c_563_n 0.0206675f $X=4.075 $Y=1.085
+ $X2=0 $Y2=0
cc_297 N_A_30_112#_c_371_p N_A_339_112#_c_613_n 0.0112667f $X=7.26 $Y=2.37 $X2=0
+ $Y2=0
cc_298 N_A_30_112#_c_319_n N_A_339_112#_c_613_n 9.68092e-19 $X=7.26 $Y=2.37
+ $X2=0 $Y2=0
cc_299 N_A_30_112#_c_384_p N_A_339_112#_c_572_n 3.15803e-19 $X=1.38 $Y=1.37
+ $X2=0 $Y2=0
cc_300 N_A_30_112#_c_334_n N_A_339_112#_c_572_n 0.0328584f $X=1.38 $Y=1.705
+ $X2=0 $Y2=0
cc_301 N_A_30_112#_c_283_n N_A_339_112#_c_572_n 0.0294849f $X=1.425 $Y=3.41
+ $X2=0 $Y2=0
cc_302 N_A_30_112#_c_292_n N_A_339_112#_c_572_n 0.0139222f $X=2.29 $Y=2.39 $X2=0
+ $Y2=0
cc_303 N_A_30_112#_c_275_n N_A_339_112#_c_572_n 0.0306932f $X=1.38 $Y=1.365
+ $X2=0 $Y2=0
cc_304 N_A_30_112#_c_384_p N_A_339_112#_c_573_n 0.0127633f $X=1.38 $Y=1.37 $X2=0
+ $Y2=0
cc_305 N_A_30_112#_c_275_n N_A_339_112#_c_573_n 0.00535051f $X=1.38 $Y=1.365
+ $X2=0 $Y2=0
cc_306 N_A_30_112#_c_266_n N_A_339_112#_c_622_n 2.22051e-19 $X=4.075 $Y=1.085
+ $X2=0 $Y2=0
cc_307 N_A_30_112#_c_266_n N_A_339_112#_c_623_n 0.00137837f $X=4.075 $Y=1.085
+ $X2=0 $Y2=0
cc_308 N_A_30_112#_c_277_n N_A_339_112#_c_624_n 5.95172e-19 $X=8.08 $Y=1.085
+ $X2=0 $Y2=0
cc_309 N_A_30_112#_c_266_n N_A_339_112#_M1018_g 0.0326122f $X=4.075 $Y=1.085
+ $X2=0 $Y2=0
cc_310 N_A_30_112#_c_273_n N_A_339_112#_M1024_g 0.0182621f $X=8.11 $Y=1.27 $X2=0
+ $Y2=0
cc_311 N_A_30_112#_c_277_n N_A_339_112#_M1024_g 0.0125297f $X=8.08 $Y=1.085
+ $X2=0 $Y2=0
cc_312 N_A_30_112#_c_306_n N_A_1063_85#_M1017_d 8.28689e-19 $X=7.095 $Y=3.72
+ $X2=0 $Y2=0
cc_313 N_A_30_112#_c_305_n N_A_1063_85#_c_729_n 0.0123662f $X=6.395 $Y=2.72
+ $X2=0 $Y2=0
cc_314 N_A_30_112#_c_371_p N_A_1063_85#_c_727_n 0.00567639f $X=7.26 $Y=2.37
+ $X2=0 $Y2=0
cc_315 N_A_30_112#_c_319_n N_A_1063_85#_c_727_n 0.00119386f $X=7.26 $Y=2.37
+ $X2=0 $Y2=0
cc_316 N_A_30_112#_c_305_n N_A_1063_85#_c_731_n 0.00897876f $X=6.395 $Y=2.72
+ $X2=13.68 $Y2=0
cc_317 N_A_30_112#_c_402_p N_A_1063_85#_c_731_n 0.0211567f $X=6.48 $Y=3.635
+ $X2=13.68 $Y2=0
cc_318 N_A_30_112#_c_306_n N_A_1063_85#_c_731_n 0.0110776f $X=7.095 $Y=3.72
+ $X2=13.68 $Y2=0
cc_319 N_A_30_112#_c_404_p N_A_1063_85#_c_731_n 0.0384152f $X=7.18 $Y=3.635
+ $X2=13.68 $Y2=0
cc_320 N_A_30_112#_c_371_p N_A_1063_85#_c_731_n 0.0027839f $X=7.26 $Y=2.37
+ $X2=13.68 $Y2=0
cc_321 N_A_30_112#_c_319_n N_A_1063_85#_c_731_n 0.00249778f $X=7.26 $Y=2.37
+ $X2=13.68 $Y2=0
cc_322 N_A_30_112#_c_281_n N_A_1063_85#_c_744_n 5.99429e-19 $X=4.855 $Y=2.645
+ $X2=6.96 $Y2=0.057
cc_323 N_A_30_112#_c_357_p N_A_1063_85#_c_744_n 0.00876288f $X=4.92 $Y=2.37
+ $X2=6.96 $Y2=0.057
cc_324 N_A_30_112#_c_305_n N_A_1063_85#_c_744_n 0.0652037f $X=6.395 $Y=2.72
+ $X2=6.96 $Y2=0.057
cc_325 N_A_30_112#_c_371_p N_A_1063_85#_c_732_n 0.0137935f $X=7.26 $Y=2.37 $X2=0
+ $Y2=0
cc_326 N_A_30_112#_c_319_n N_A_1063_85#_c_732_n 0.0016316f $X=7.26 $Y=2.37 $X2=0
+ $Y2=0
cc_327 N_A_30_112#_c_281_n N_A_1063_85#_M1021_g 0.0707818f $X=4.855 $Y=2.645
+ $X2=0 $Y2=0
cc_328 N_A_30_112#_c_357_p N_A_1063_85#_M1021_g 0.00206163f $X=4.92 $Y=2.37
+ $X2=0 $Y2=0
cc_329 N_A_30_112#_c_304_n N_A_1063_85#_M1021_g 0.00155612f $X=4.92 $Y=3.335
+ $X2=0 $Y2=0
cc_330 N_A_30_112#_c_305_n N_A_1063_85#_M1021_g 0.0275132f $X=6.395 $Y=2.72
+ $X2=0 $Y2=0
cc_331 N_A_30_112#_c_402_p N_A_1063_85#_M1021_g 0.00101104f $X=6.48 $Y=3.635
+ $X2=0 $Y2=0
cc_332 N_A_30_112#_c_266_n N_A_865_111#_c_786_n 0.013981f $X=4.075 $Y=1.085
+ $X2=0 $Y2=0
cc_333 N_A_30_112#_c_348_p N_A_865_111#_c_786_n 0.0544512f $X=3.965 $Y=1.28
+ $X2=0 $Y2=0
cc_334 N_A_30_112#_c_281_n N_A_865_111#_c_790_n 0.00559049f $X=4.855 $Y=2.645
+ $X2=0.24 $Y2=0
cc_335 N_A_30_112#_c_271_n N_A_865_111#_c_790_n 0.0719568f $X=4.035 $Y=3.335
+ $X2=0.24 $Y2=0
cc_336 N_A_30_112#_c_301_n N_A_865_111#_c_790_n 0.0182867f $X=4.755 $Y=3.42
+ $X2=0.24 $Y2=0
cc_337 N_A_30_112#_c_357_p N_A_865_111#_c_790_n 0.0255344f $X=4.92 $Y=2.37
+ $X2=0.24 $Y2=0
cc_338 N_A_30_112#_c_304_n N_A_865_111#_c_790_n 0.0126374f $X=4.92 $Y=3.335
+ $X2=0.24 $Y2=0
cc_339 N_A_30_112#_c_424_p N_A_865_111#_c_790_n 0.00819387f $X=4.92 $Y=2.72
+ $X2=0.24 $Y2=0
cc_340 N_A_30_112#_c_281_n N_A_865_111#_c_791_n 0.00534014f $X=4.855 $Y=2.645
+ $X2=0 $Y2=0
cc_341 N_A_30_112#_c_357_p N_A_865_111#_c_791_n 0.0250952f $X=4.92 $Y=2.37 $X2=0
+ $Y2=0
cc_342 N_A_30_112#_c_305_n N_A_865_111#_c_791_n 0.0105357f $X=6.395 $Y=2.72
+ $X2=0 $Y2=0
cc_343 N_A_30_112#_c_266_n N_A_865_111#_c_787_n 0.0111722f $X=4.075 $Y=1.085
+ $X2=13.68 $Y2=0
cc_344 N_A_30_112#_c_271_n N_A_865_111#_c_792_n 0.0131177f $X=4.035 $Y=3.335
+ $X2=0 $Y2=0
cc_345 N_A_30_112#_c_305_n N_A_865_111#_M1023_g 0.023505f $X=6.395 $Y=2.72 $X2=0
+ $Y2=0
cc_346 N_A_30_112#_c_402_p N_A_865_111#_M1023_g 0.0313291f $X=6.48 $Y=3.635
+ $X2=0 $Y2=0
cc_347 N_A_30_112#_c_306_n N_A_865_111#_M1023_g 0.0071006f $X=7.095 $Y=3.72
+ $X2=0 $Y2=0
cc_348 N_A_30_112#_c_309_n N_A_865_111#_M1023_g 0.00541751f $X=6.565 $Y=3.72
+ $X2=0 $Y2=0
cc_349 N_A_30_112#_c_404_p N_A_865_111#_M1023_g 8.52474e-19 $X=7.18 $Y=3.635
+ $X2=0 $Y2=0
cc_350 N_A_30_112#_c_319_n N_A_865_111#_M1023_g 0.0417779f $X=7.26 $Y=2.37 $X2=0
+ $Y2=0
cc_351 N_A_30_112#_c_272_n N_A_1711_85#_M1016_g 0.00138972f $X=8.11 $Y=1.27
+ $X2=0 $Y2=0
cc_352 N_A_30_112#_c_277_n N_A_1711_85#_M1016_g 0.0668216f $X=8.08 $Y=1.085
+ $X2=0 $Y2=0
cc_353 N_A_30_112#_c_272_n N_A_1711_85#_M1008_g 0.0016306f $X=8.11 $Y=1.27 $X2=0
+ $Y2=0
cc_354 N_A_30_112#_c_272_n N_A_1711_85#_c_868_n 7.14182e-19 $X=8.11 $Y=1.27
+ $X2=0 $Y2=0
cc_355 N_A_30_112#_c_311_n N_A_1494_539#_M1000_d 0.00131594f $X=7.975 $Y=3.72
+ $X2=0 $Y2=0
cc_356 N_A_30_112#_c_311_n N_A_1494_539#_c_990_n 0.0212448f $X=7.975 $Y=3.72
+ $X2=13.68 $Y2=0
cc_357 N_A_30_112#_c_319_n N_A_1494_539#_c_990_n 0.012018f $X=7.26 $Y=2.37
+ $X2=13.68 $Y2=0
cc_358 N_A_30_112#_c_272_n N_A_1494_539#_c_979_n 0.00791264f $X=8.11 $Y=1.27
+ $X2=0 $Y2=0
cc_359 N_A_30_112#_c_277_n N_A_1494_539#_c_979_n 0.0304298f $X=8.08 $Y=1.085
+ $X2=0 $Y2=0
cc_360 N_A_30_112#_c_272_n N_A_1494_539#_c_983_n 0.0873067f $X=8.11 $Y=1.27
+ $X2=0 $Y2=0
cc_361 N_A_30_112#_c_277_n N_A_1494_539#_c_983_n 0.00748307f $X=8.08 $Y=1.085
+ $X2=0 $Y2=0
cc_362 N_A_30_112#_c_272_n N_A_1494_539#_c_993_n 0.0135452f $X=8.11 $Y=1.27
+ $X2=0 $Y2=0
cc_363 N_A_30_112#_c_404_p N_A_1494_539#_c_995_n 0.0533485f $X=7.18 $Y=3.635
+ $X2=0 $Y2=0
cc_364 N_A_30_112#_c_319_n N_A_1494_539#_c_995_n 0.00375255f $X=7.26 $Y=2.37
+ $X2=0 $Y2=0
cc_365 N_A_30_112#_c_404_p N_A_1494_539#_c_985_n 0.00733919f $X=7.18 $Y=3.635
+ $X2=0 $Y2=0
cc_366 N_A_30_112#_c_272_n N_A_1494_539#_c_985_n 0.153199f $X=8.11 $Y=1.27 $X2=0
+ $Y2=0
cc_367 N_A_30_112#_c_273_n N_A_1494_539#_c_985_n 0.00330621f $X=8.11 $Y=1.27
+ $X2=0 $Y2=0
cc_368 N_A_30_112#_c_371_p N_A_1494_539#_c_985_n 0.0192366f $X=7.26 $Y=2.37
+ $X2=0 $Y2=0
cc_369 N_A_30_112#_c_319_n N_A_1494_539#_c_985_n 0.00464212f $X=7.26 $Y=2.37
+ $X2=0 $Y2=0
cc_370 N_A_30_112#_c_277_n N_A_1494_539#_c_986_n 0.00164554f $X=8.08 $Y=1.085
+ $X2=0 $Y2=0
cc_371 N_A_30_112#_c_305_n N_VPWR_M1015_d 0.00293905f $X=6.395 $Y=2.72 $X2=0
+ $Y2=0
cc_372 N_A_30_112#_M1022_g N_VPWR_c_1125_n 0.00220539f $X=1.465 $Y=2.815 $X2=0
+ $Y2=0
cc_373 N_A_30_112#_c_269_n N_VPWR_c_1125_n 0.0340456f $X=0.295 $Y=2.565 $X2=0
+ $Y2=0
cc_374 N_A_30_112#_c_283_n N_VPWR_c_1125_n 0.044259f $X=1.425 $Y=3.41 $X2=0
+ $Y2=0
cc_375 N_A_30_112#_c_287_n N_VPWR_c_1125_n 0.0125296f $X=1.51 $Y=3.495 $X2=0
+ $Y2=0
cc_376 N_A_30_112#_c_284_n N_VPWR_c_1128_n 0.0124892f $X=2.12 $Y=3.495 $X2=0
+ $Y2=0
cc_377 N_A_30_112#_c_290_n N_VPWR_c_1128_n 0.0597013f $X=2.205 $Y=3.41 $X2=0
+ $Y2=0
cc_378 N_A_30_112#_c_291_n N_VPWR_c_1128_n 0.0428236f $X=3.18 $Y=2.39 $X2=0
+ $Y2=0
cc_379 N_A_30_112#_c_293_n N_VPWR_c_1128_n 0.0333954f $X=3.265 $Y=3.335 $X2=0
+ $Y2=0
cc_380 N_A_30_112#_c_297_n N_VPWR_c_1128_n 0.013855f $X=3.35 $Y=3.42 $X2=0 $Y2=0
cc_381 N_A_30_112#_c_281_n N_VPWR_c_1131_n 0.00131903f $X=4.855 $Y=2.645 $X2=0
+ $Y2=0
cc_382 N_A_30_112#_c_301_n N_VPWR_c_1131_n 0.0141178f $X=4.755 $Y=3.42 $X2=0
+ $Y2=0
cc_383 N_A_30_112#_c_304_n N_VPWR_c_1131_n 0.0227056f $X=4.92 $Y=3.335 $X2=0
+ $Y2=0
cc_384 N_A_30_112#_c_305_n N_VPWR_c_1131_n 0.0582416f $X=6.395 $Y=2.72 $X2=0
+ $Y2=0
cc_385 N_A_30_112#_c_402_p N_VPWR_c_1131_n 0.0450675f $X=6.48 $Y=3.635 $X2=0
+ $Y2=0
cc_386 N_A_30_112#_c_309_n N_VPWR_c_1131_n 0.00492718f $X=6.565 $Y=3.72 $X2=0
+ $Y2=0
cc_387 N_A_30_112#_c_311_n N_VPWR_c_1134_n 0.0039033f $X=7.975 $Y=3.72 $X2=0
+ $Y2=0
cc_388 N_A_30_112#_c_272_n N_VPWR_c_1134_n 0.0418828f $X=8.11 $Y=1.27 $X2=0
+ $Y2=0
cc_389 N_A_30_112#_M1022_g N_VPWR_c_1143_n 0.0040826f $X=1.465 $Y=2.815 $X2=0
+ $Y2=0
cc_390 N_A_30_112#_c_281_n N_VPWR_c_1143_n 6.53579e-19 $X=4.855 $Y=2.645 $X2=0
+ $Y2=0
cc_391 N_A_30_112#_c_269_n N_VPWR_c_1143_n 0.0146884f $X=0.295 $Y=2.565 $X2=0
+ $Y2=0
cc_392 N_A_30_112#_c_284_n N_VPWR_c_1143_n 0.0499525f $X=2.12 $Y=3.495 $X2=0
+ $Y2=0
cc_393 N_A_30_112#_c_287_n N_VPWR_c_1143_n 0.0113249f $X=1.51 $Y=3.495 $X2=0
+ $Y2=0
cc_394 N_A_30_112#_c_294_n N_VPWR_c_1143_n 0.0278131f $X=3.95 $Y=3.42 $X2=0
+ $Y2=0
cc_395 N_A_30_112#_c_297_n N_VPWR_c_1143_n 0.00968423f $X=3.35 $Y=3.42 $X2=0
+ $Y2=0
cc_396 N_A_30_112#_c_301_n N_VPWR_c_1143_n 0.0476017f $X=4.755 $Y=3.42 $X2=0
+ $Y2=0
cc_397 N_A_30_112#_c_402_p N_VPWR_c_1143_n 0.0190049f $X=6.48 $Y=3.635 $X2=0
+ $Y2=0
cc_398 N_A_30_112#_c_306_n N_VPWR_c_1143_n 0.0199613f $X=7.095 $Y=3.72 $X2=0
+ $Y2=0
cc_399 N_A_30_112#_c_309_n N_VPWR_c_1143_n 0.00674178f $X=6.565 $Y=3.72 $X2=0
+ $Y2=0
cc_400 N_A_30_112#_c_404_p N_VPWR_c_1143_n 0.0220458f $X=7.18 $Y=3.635 $X2=0
+ $Y2=0
cc_401 N_A_30_112#_c_311_n N_VPWR_c_1143_n 0.0361699f $X=7.975 $Y=3.72 $X2=0
+ $Y2=0
cc_402 N_A_30_112#_c_272_n N_VPWR_c_1143_n 0.0222621f $X=8.11 $Y=1.27 $X2=0
+ $Y2=0
cc_403 N_A_30_112#_c_316_n N_VPWR_c_1143_n 0.00901673f $X=4.035 $Y=3.42 $X2=0
+ $Y2=0
cc_404 N_A_30_112#_c_319_n N_VPWR_c_1143_n 0.0172808f $X=7.26 $Y=2.37 $X2=0
+ $Y2=0
cc_405 N_A_30_112#_c_322_n N_VPWR_c_1143_n 0.00353126f $X=7.18 $Y=3.72 $X2=0
+ $Y2=0
cc_406 N_A_30_112#_c_271_n N_A_709_111#_c_1224_n 0.019156f $X=4.035 $Y=3.335
+ $X2=0 $Y2=0
cc_407 N_A_30_112#_c_294_n N_A_709_111#_c_1225_n 0.0174665f $X=3.95 $Y=3.42
+ $X2=0.24 $Y2=0
cc_408 N_A_30_112#_c_266_n N_A_709_111#_c_1229_n 0.011591f $X=4.075 $Y=1.085
+ $X2=0 $Y2=0
cc_409 N_A_30_112#_c_266_n N_A_709_111#_c_1223_n 0.00675884f $X=4.075 $Y=1.085
+ $X2=13.68 $Y2=0
cc_410 N_A_30_112#_c_291_n N_A_709_111#_c_1223_n 0.0123662f $X=3.18 $Y=2.39
+ $X2=13.68 $Y2=0
cc_411 N_A_30_112#_c_293_n N_A_709_111#_c_1223_n 0.0448079f $X=3.265 $Y=3.335
+ $X2=13.68 $Y2=0
cc_412 N_A_30_112#_c_348_p N_A_709_111#_c_1223_n 0.0470461f $X=3.965 $Y=1.28
+ $X2=13.68 $Y2=0
cc_413 N_A_30_112#_c_271_n N_A_709_111#_c_1223_n 0.0474085f $X=4.035 $Y=3.335
+ $X2=13.68 $Y2=0
cc_414 N_A_30_112#_c_305_n A_1021_539# 0.00366293f $X=6.395 $Y=2.72 $X2=0 $Y2=0
cc_415 N_A_30_112#_M1004_g N_VGND_c_1302_n 0.0402642f $X=1.445 $Y=0.77 $X2=0
+ $Y2=0
cc_416 N_A_30_112#_c_267_n N_VGND_c_1302_n 0.0351962f $X=0.275 $Y=0.77 $X2=0
+ $Y2=0
cc_417 N_A_30_112#_c_270_n N_VGND_c_1302_n 0.0441137f $X=1.215 $Y=1.285 $X2=0
+ $Y2=0
cc_418 N_A_30_112#_c_384_p N_VGND_c_1302_n 0.0257617f $X=1.38 $Y=1.37 $X2=0
+ $Y2=0
cc_419 N_A_30_112#_M1004_g N_VGND_c_1304_n 0.00214016f $X=1.445 $Y=0.77 $X2=0
+ $Y2=0
cc_420 N_A_30_112#_c_277_n N_VGND_c_1308_n 0.00101203f $X=8.08 $Y=1.085 $X2=0
+ $Y2=0
cc_421 N_A_30_112#_M1004_g N_VGND_c_1314_n 0.00940063f $X=1.445 $Y=0.77 $X2=0
+ $Y2=0
cc_422 N_A_30_112#_c_266_n N_VGND_c_1314_n 0.0159214f $X=4.075 $Y=1.085 $X2=0
+ $Y2=0
cc_423 N_A_30_112#_c_267_n N_VGND_c_1314_n 0.0305594f $X=0.275 $Y=0.77 $X2=0
+ $Y2=0
cc_424 N_A_30_112#_c_270_n N_VGND_c_1314_n 0.00680911f $X=1.215 $Y=1.285 $X2=0
+ $Y2=0
cc_425 N_A_30_112#_c_384_p N_VGND_c_1314_n 0.00115862f $X=1.38 $Y=1.37 $X2=0
+ $Y2=0
cc_426 N_A_30_112#_c_348_p N_VGND_c_1314_n 0.0081908f $X=3.965 $Y=1.28 $X2=0
+ $Y2=0
cc_427 N_A_30_112#_c_272_n N_VGND_c_1314_n 0.00170486f $X=8.11 $Y=1.27 $X2=0
+ $Y2=0
cc_428 N_A_30_112#_c_275_n N_VGND_c_1314_n 5.12378e-19 $X=1.38 $Y=1.365 $X2=0
+ $Y2=0
cc_429 N_A_30_112#_c_277_n N_VGND_c_1314_n 0.00647473f $X=8.08 $Y=1.085 $X2=0
+ $Y2=0
cc_430 N_D_c_521_n N_A_339_112#_c_558_n 0.0192786f $X=3.272 $Y=2.19 $X2=0 $Y2=0
cc_431 N_D_M1006_g N_A_339_112#_M1019_g 0.0192786f $X=3.295 $Y=2.905 $X2=0 $Y2=0
cc_432 N_D_c_517_n N_A_339_112#_c_562_n 0.0207418f $X=3.272 $Y=1.377 $X2=0 $Y2=0
cc_433 N_D_c_519_n N_A_339_112#_c_562_n 0.0634044f $X=3.185 $Y=1.665 $X2=0 $Y2=0
cc_434 N_D_M1013_g N_A_339_112#_c_611_n 0.0285066f $X=3.295 $Y=0.765 $X2=0 $Y2=0
cc_435 N_D_c_517_n N_A_339_112#_c_611_n 0.00605373f $X=3.272 $Y=1.377 $X2=0
+ $Y2=0
cc_436 N_D_M1013_g N_A_339_112#_c_563_n 0.00838107f $X=3.295 $Y=0.765 $X2=0
+ $Y2=0
cc_437 N_D_M1013_g N_A_339_112#_c_565_n 0.00319605f $X=3.295 $Y=0.765 $X2=0
+ $Y2=0
cc_438 N_D_c_519_n N_A_339_112#_c_572_n 0.020788f $X=3.185 $Y=1.665 $X2=0 $Y2=0
cc_439 N_D_M1006_g N_VPWR_c_1128_n 0.00575003f $X=3.295 $Y=2.905 $X2=0 $Y2=0
cc_440 N_D_M1006_g N_VPWR_c_1143_n 0.00421533f $X=3.295 $Y=2.905 $X2=0 $Y2=0
cc_441 N_D_M1006_g N_A_709_111#_c_1224_n 0.00236737f $X=3.295 $Y=2.905 $X2=0
+ $Y2=0
cc_442 N_D_M1006_g N_A_709_111#_c_1225_n 0.00649712f $X=3.295 $Y=2.905 $X2=0.24
+ $Y2=0
cc_443 N_D_M1013_g N_A_709_111#_c_1229_n 0.00588258f $X=3.295 $Y=0.765 $X2=0
+ $Y2=0
cc_444 N_D_M1013_g N_A_709_111#_c_1223_n 0.00362844f $X=3.295 $Y=0.765 $X2=13.68
+ $Y2=0
cc_445 N_D_M1006_g N_A_709_111#_c_1223_n 0.0137258f $X=3.295 $Y=2.905 $X2=13.68
+ $Y2=0
cc_446 N_D_c_517_n N_A_709_111#_c_1223_n 0.0061619f $X=3.272 $Y=1.377 $X2=13.68
+ $Y2=0
cc_447 N_D_c_521_n N_A_709_111#_c_1223_n 0.00883535f $X=3.272 $Y=2.19 $X2=13.68
+ $Y2=0
cc_448 N_D_c_518_n N_A_709_111#_c_1223_n 0.0176248f $X=3.185 $Y=1.665 $X2=13.68
+ $Y2=0
cc_449 N_D_c_519_n N_A_709_111#_c_1223_n 0.0419725f $X=3.185 $Y=1.665 $X2=13.68
+ $Y2=0
cc_450 N_D_M1013_g N_VGND_c_1304_n 0.0143015f $X=3.295 $Y=0.765 $X2=0 $Y2=0
cc_451 N_D_M1013_g N_VGND_c_1314_n 0.0157471f $X=3.295 $Y=0.765 $X2=0 $Y2=0
cc_452 N_D_c_517_n N_VGND_c_1314_n 0.00118275f $X=3.272 $Y=1.377 $X2=0 $Y2=0
cc_453 N_A_339_112#_c_637_p N_A_1063_85#_c_725_n 0.0428346f $X=6.4 $Y=1.245
+ $X2=0.24 $Y2=0
cc_454 N_A_339_112#_c_568_n N_A_1063_85#_c_725_n 0.0209527f $X=7.175 $Y=0.35
+ $X2=0.24 $Y2=0
cc_455 N_A_339_112#_c_624_n N_A_1063_85#_c_725_n 0.0254843f $X=7.31 $Y=1.195
+ $X2=0.24 $Y2=0
cc_456 N_A_339_112#_M1024_g N_A_1063_85#_c_725_n 0.00722721f $X=7.315 $Y=0.765
+ $X2=0.24 $Y2=0
cc_457 N_A_339_112#_c_567_n N_A_1063_85#_c_726_n 0.0060982f $X=6.315 $Y=1.33
+ $X2=0 $Y2=0
cc_458 N_A_339_112#_c_642_p N_A_1063_85#_c_726_n 0.0254843f $X=7.31 $Y=1.33
+ $X2=0 $Y2=0
cc_459 N_A_339_112#_c_567_n N_A_1063_85#_c_727_n 0.00519058f $X=6.315 $Y=1.33
+ $X2=0 $Y2=0
cc_460 N_A_339_112#_c_642_p N_A_1063_85#_c_727_n 0.0290197f $X=7.31 $Y=1.33
+ $X2=0 $Y2=0
cc_461 N_A_339_112#_M1024_g N_A_1063_85#_c_727_n 0.00774939f $X=7.315 $Y=0.765
+ $X2=0 $Y2=0
cc_462 N_A_339_112#_c_567_n N_A_1063_85#_M1021_g 0.0312441f $X=6.315 $Y=1.33
+ $X2=0 $Y2=0
cc_463 N_A_339_112#_c_637_p N_A_1063_85#_M1021_g 0.00146975f $X=6.4 $Y=1.245
+ $X2=0 $Y2=0
cc_464 N_A_339_112#_c_622_n N_A_1063_85#_M1021_g 0.00181092f $X=4.815 $Y=1.295
+ $X2=0 $Y2=0
cc_465 N_A_339_112#_c_623_n N_A_1063_85#_M1021_g 0.00163063f $X=4.815 $Y=1.195
+ $X2=0 $Y2=0
cc_466 N_A_339_112#_M1018_g N_A_1063_85#_M1021_g 0.109616f $X=4.855 $Y=0.765
+ $X2=0 $Y2=0
cc_467 N_A_339_112#_c_558_n N_A_865_111#_c_786_n 0.0172305f $X=4.075 $Y=2.185
+ $X2=0 $Y2=0
cc_468 N_A_339_112#_c_622_n N_A_865_111#_c_786_n 0.0378138f $X=4.815 $Y=1.295
+ $X2=0 $Y2=0
cc_469 N_A_339_112#_c_623_n N_A_865_111#_c_786_n 0.00764027f $X=4.815 $Y=1.195
+ $X2=0 $Y2=0
cc_470 N_A_339_112#_M1018_g N_A_865_111#_c_786_n 0.00542639f $X=4.855 $Y=0.765
+ $X2=0 $Y2=0
cc_471 N_A_339_112#_c_558_n N_A_865_111#_c_790_n 0.0110512f $X=4.075 $Y=2.185
+ $X2=0.24 $Y2=0
cc_472 N_A_339_112#_M1019_g N_A_865_111#_c_790_n 0.0222283f $X=4.075 $Y=2.905
+ $X2=0.24 $Y2=0
cc_473 N_A_339_112#_c_558_n N_A_865_111#_c_791_n 0.0206522f $X=4.075 $Y=2.185
+ $X2=0 $Y2=0
cc_474 N_A_339_112#_c_567_n N_A_865_111#_c_791_n 0.0396457f $X=6.315 $Y=1.33
+ $X2=0 $Y2=0
cc_475 N_A_339_112#_c_622_n N_A_865_111#_c_791_n 0.0236215f $X=4.815 $Y=1.295
+ $X2=0 $Y2=0
cc_476 N_A_339_112#_c_558_n N_A_865_111#_c_787_n 0.00359469f $X=4.075 $Y=2.185
+ $X2=13.68 $Y2=0
cc_477 N_A_339_112#_c_563_n N_A_865_111#_c_787_n 0.0198871f $X=4.81 $Y=0.35
+ $X2=13.68 $Y2=0
cc_478 N_A_339_112#_c_623_n N_A_865_111#_c_787_n 0.0272138f $X=4.815 $Y=1.195
+ $X2=13.68 $Y2=0
cc_479 N_A_339_112#_M1018_g N_A_865_111#_c_787_n 0.00836329f $X=4.855 $Y=0.765
+ $X2=13.68 $Y2=0
cc_480 N_A_339_112#_c_558_n N_A_865_111#_c_792_n 0.0128473f $X=4.075 $Y=2.185
+ $X2=0 $Y2=0
cc_481 N_A_339_112#_c_567_n N_A_865_111#_c_829_n 0.0207976f $X=6.315 $Y=1.33
+ $X2=6.96 $Y2=0
cc_482 N_A_339_112#_c_567_n N_A_865_111#_M1023_g 0.0193817f $X=6.315 $Y=1.33
+ $X2=0 $Y2=0
cc_483 N_A_339_112#_c_637_p N_A_865_111#_M1023_g 0.0324204f $X=6.4 $Y=1.245
+ $X2=0 $Y2=0
cc_484 N_A_339_112#_c_568_n N_A_865_111#_M1023_g 0.00840832f $X=7.175 $Y=0.35
+ $X2=0 $Y2=0
cc_485 N_A_339_112#_c_570_n N_A_865_111#_M1023_g 0.00319589f $X=6.485 $Y=0.35
+ $X2=0 $Y2=0
cc_486 N_A_339_112#_c_624_n N_A_865_111#_M1023_g 0.00135049f $X=7.31 $Y=1.195
+ $X2=0 $Y2=0
cc_487 N_A_339_112#_M1024_g N_A_865_111#_M1023_g 0.0352403f $X=7.315 $Y=0.765
+ $X2=0 $Y2=0
cc_488 N_A_339_112#_M1002_g N_A_1711_85#_M1008_g 0.041637f $X=8.095 $Y=2.905
+ $X2=0 $Y2=0
cc_489 N_A_339_112#_c_559_n N_A_1711_85#_c_868_n 0.058834f $X=7.315 $Y=1.665
+ $X2=0 $Y2=0
cc_490 N_A_339_112#_c_624_n N_A_1494_539#_c_1013_n 0.0206198f $X=7.31 $Y=1.195
+ $X2=0 $Y2=0
cc_491 N_A_339_112#_M1024_g N_A_1494_539#_c_1013_n 0.00344306f $X=7.315 $Y=0.765
+ $X2=0 $Y2=0
cc_492 N_A_339_112#_c_624_n N_A_1494_539#_c_981_n 0.0102933f $X=7.31 $Y=1.195
+ $X2=0 $Y2=0
cc_493 N_A_339_112#_M1024_g N_A_1494_539#_c_981_n 0.00312065f $X=7.315 $Y=0.765
+ $X2=0 $Y2=0
cc_494 N_A_339_112#_c_559_n N_A_1494_539#_c_983_n 0.00467238f $X=7.315 $Y=1.665
+ $X2=0 $Y2=0
cc_495 N_A_339_112#_c_559_n N_A_1494_539#_c_993_n 0.00135748f $X=7.315 $Y=1.665
+ $X2=0 $Y2=0
cc_496 N_A_339_112#_c_559_n N_A_1494_539#_c_995_n 0.00427724f $X=7.315 $Y=1.665
+ $X2=0 $Y2=0
cc_497 N_A_339_112#_M1002_g N_A_1494_539#_c_985_n 0.00572804f $X=8.095 $Y=2.905
+ $X2=0 $Y2=0
cc_498 N_A_339_112#_c_559_n N_A_1494_539#_c_985_n 0.0351763f $X=7.315 $Y=1.665
+ $X2=0 $Y2=0
cc_499 N_A_339_112#_c_642_p N_A_1494_539#_c_985_n 0.0466752f $X=7.31 $Y=1.33
+ $X2=0 $Y2=0
cc_500 N_A_339_112#_c_624_n N_A_1494_539#_c_985_n 0.00882626f $X=7.31 $Y=1.195
+ $X2=0 $Y2=0
cc_501 N_A_339_112#_M1024_g N_A_1494_539#_c_985_n 0.00958912f $X=7.315 $Y=0.765
+ $X2=0 $Y2=0
cc_502 N_A_339_112#_c_559_n N_A_1494_539#_c_986_n 0.00154311f $X=7.315 $Y=1.665
+ $X2=0 $Y2=0
cc_503 N_A_339_112#_M1024_g N_A_1494_539#_c_986_n 0.00388684f $X=7.315 $Y=0.765
+ $X2=0 $Y2=0
cc_504 N_A_339_112#_M1002_g N_VPWR_c_1134_n 0.00264766f $X=8.095 $Y=2.905 $X2=0
+ $Y2=0
cc_505 N_A_339_112#_M1002_g N_VPWR_c_1143_n 0.00718544f $X=8.095 $Y=2.905 $X2=0
+ $Y2=0
cc_506 N_A_339_112#_c_583_n N_VPWR_c_1143_n 0.0018836f $X=1.855 $Y=2.565 $X2=0
+ $Y2=0
cc_507 N_A_339_112#_M1019_g N_A_709_111#_c_1224_n 8.56501e-19 $X=4.075 $Y=2.905
+ $X2=0 $Y2=0
cc_508 N_A_339_112#_c_611_n N_A_709_111#_c_1229_n 0.0217567f $X=3.255 $Y=1.195
+ $X2=0 $Y2=0
cc_509 N_A_339_112#_c_563_n N_A_709_111#_c_1229_n 0.0198711f $X=4.81 $Y=0.35
+ $X2=0 $Y2=0
cc_510 N_A_339_112#_c_558_n N_A_709_111#_c_1223_n 0.00549146f $X=4.075 $Y=2.185
+ $X2=13.68 $Y2=0
cc_511 N_A_339_112#_c_562_n N_A_709_111#_c_1223_n 0.0118397f $X=3.17 $Y=1.28
+ $X2=13.68 $Y2=0
cc_512 N_A_339_112#_c_611_n N_A_709_111#_c_1223_n 0.0159966f $X=3.255 $Y=1.195
+ $X2=13.68 $Y2=0
cc_513 N_A_339_112#_c_567_n N_VGND_M1021_d 0.00231909f $X=6.315 $Y=1.33 $X2=0
+ $Y2=0
cc_514 N_A_339_112#_c_560_n N_VGND_c_1302_n 0.0228606f $X=1.835 $Y=0.77 $X2=0
+ $Y2=0
cc_515 N_A_339_112#_c_560_n N_VGND_c_1304_n 0.0381207f $X=1.835 $Y=0.77 $X2=0
+ $Y2=0
cc_516 N_A_339_112#_c_562_n N_VGND_c_1304_n 0.0697162f $X=3.17 $Y=1.28 $X2=0
+ $Y2=0
cc_517 N_A_339_112#_c_611_n N_VGND_c_1304_n 0.0254957f $X=3.255 $Y=1.195 $X2=0
+ $Y2=0
cc_518 N_A_339_112#_c_565_n N_VGND_c_1304_n 0.00485941f $X=3.34 $Y=0.35 $X2=0
+ $Y2=0
cc_519 N_A_339_112#_c_563_n N_VGND_c_1306_n 0.00422833f $X=4.81 $Y=0.35 $X2=0
+ $Y2=0
cc_520 N_A_339_112#_c_567_n N_VGND_c_1306_n 0.0719024f $X=6.315 $Y=1.33 $X2=0
+ $Y2=0
cc_521 N_A_339_112#_c_637_p N_VGND_c_1306_n 0.025472f $X=6.4 $Y=1.245 $X2=0
+ $Y2=0
cc_522 N_A_339_112#_c_570_n N_VGND_c_1306_n 0.00481634f $X=6.485 $Y=0.35 $X2=0
+ $Y2=0
cc_523 N_A_339_112#_c_623_n N_VGND_c_1306_n 0.0409055f $X=4.815 $Y=1.195 $X2=0
+ $Y2=0
cc_524 N_A_339_112#_M1018_g N_VGND_c_1306_n 0.00492682f $X=4.855 $Y=0.765 $X2=0
+ $Y2=0
cc_525 N_A_339_112#_M1004_d N_VGND_c_1314_n 0.00261451f $X=1.695 $Y=0.56 $X2=0
+ $Y2=0
cc_526 N_A_339_112#_c_560_n N_VGND_c_1314_n 0.0165746f $X=1.835 $Y=0.77 $X2=0
+ $Y2=0
cc_527 N_A_339_112#_c_562_n N_VGND_c_1314_n 0.0136799f $X=3.17 $Y=1.28 $X2=0
+ $Y2=0
cc_528 N_A_339_112#_c_611_n N_VGND_c_1314_n 0.0199629f $X=3.255 $Y=1.195 $X2=0
+ $Y2=0
cc_529 N_A_339_112#_c_563_n N_VGND_c_1314_n 0.059123f $X=4.81 $Y=0.35 $X2=0
+ $Y2=0
cc_530 N_A_339_112#_c_565_n N_VGND_c_1314_n 0.00776317f $X=3.34 $Y=0.35 $X2=0
+ $Y2=0
cc_531 N_A_339_112#_c_637_p N_VGND_c_1314_n 0.0199533f $X=6.4 $Y=1.245 $X2=0
+ $Y2=0
cc_532 N_A_339_112#_c_568_n N_VGND_c_1314_n 0.0340299f $X=7.175 $Y=0.35 $X2=0
+ $Y2=0
cc_533 N_A_339_112#_c_570_n N_VGND_c_1314_n 0.00778401f $X=6.485 $Y=0.35 $X2=0
+ $Y2=0
cc_534 N_A_339_112#_c_642_p N_VGND_c_1314_n 0.00312631f $X=7.31 $Y=1.33 $X2=0
+ $Y2=0
cc_535 N_A_339_112#_c_573_n N_VGND_c_1314_n 7.85374e-19 $X=1.845 $Y=1.28 $X2=0
+ $Y2=0
cc_536 N_A_339_112#_c_622_n N_VGND_c_1314_n 0.00488823f $X=4.815 $Y=1.295 $X2=0
+ $Y2=0
cc_537 N_A_339_112#_c_623_n N_VGND_c_1314_n 0.0201864f $X=4.815 $Y=1.195 $X2=0
+ $Y2=0
cc_538 N_A_339_112#_c_624_n N_VGND_c_1314_n 0.0213675f $X=7.31 $Y=1.195 $X2=0
+ $Y2=0
cc_539 N_A_339_112#_M1018_g N_VGND_c_1314_n 0.0124829f $X=4.855 $Y=0.765 $X2=0
+ $Y2=0
cc_540 N_A_339_112#_M1024_g N_VGND_c_1314_n 0.0153564f $X=7.315 $Y=0.765 $X2=0
+ $Y2=0
cc_541 N_A_1063_85#_c_729_n N_A_865_111#_c_791_n 0.0283298f $X=6.745 $Y=2.37
+ $X2=0 $Y2=0
cc_542 N_A_1063_85#_c_744_n N_A_865_111#_c_791_n 0.0216359f $X=5.765 $Y=2.355
+ $X2=0 $Y2=0
cc_543 N_A_1063_85#_M1021_g N_A_865_111#_c_791_n 0.034016f $X=5.565 $Y=0.765
+ $X2=0 $Y2=0
cc_544 N_A_1063_85#_c_729_n N_A_865_111#_c_829_n 0.0232944f $X=6.745 $Y=2.37
+ $X2=6.96 $Y2=0
cc_545 N_A_1063_85#_c_727_n N_A_865_111#_c_829_n 0.0332953f $X=6.83 $Y=2.285
+ $X2=6.96 $Y2=0
cc_546 N_A_1063_85#_M1021_g N_A_865_111#_c_829_n 0.00233339f $X=5.565 $Y=0.765
+ $X2=6.96 $Y2=0
cc_547 N_A_1063_85#_c_729_n N_A_865_111#_M1023_g 0.0343437f $X=6.745 $Y=2.37
+ $X2=0 $Y2=0
cc_548 N_A_1063_85#_c_725_n N_A_865_111#_M1023_g 0.0100708f $X=6.83 $Y=0.7 $X2=0
+ $Y2=0
cc_549 N_A_1063_85#_c_726_n N_A_865_111#_M1023_g 0.00422531f $X=6.83 $Y=1.325
+ $X2=0 $Y2=0
cc_550 N_A_1063_85#_c_727_n N_A_865_111#_M1023_g 0.0195782f $X=6.83 $Y=2.285
+ $X2=0 $Y2=0
cc_551 N_A_1063_85#_c_731_n N_A_865_111#_M1023_g 0.00547527f $X=6.83 $Y=2.82
+ $X2=0 $Y2=0
cc_552 N_A_1063_85#_M1021_g N_A_865_111#_M1023_g 0.0899344f $X=5.565 $Y=0.765
+ $X2=0 $Y2=0
cc_553 N_A_1063_85#_M1021_g N_VPWR_c_1131_n 0.0353945f $X=5.565 $Y=0.765 $X2=0
+ $Y2=0
cc_554 N_A_1063_85#_M1017_d N_VPWR_c_1143_n 0.00442064f $X=6.69 $Y=2.695 $X2=0
+ $Y2=0
cc_555 N_A_1063_85#_c_731_n N_VPWR_c_1143_n 0.0117439f $X=6.83 $Y=2.82 $X2=0
+ $Y2=0
cc_556 N_A_1063_85#_M1021_g N_VGND_c_1306_n 0.0566471f $X=5.565 $Y=0.765 $X2=0
+ $Y2=0
cc_557 N_A_1063_85#_M1023_d N_VGND_c_1314_n 0.002961f $X=6.69 $Y=0.555 $X2=0
+ $Y2=0
cc_558 N_A_1063_85#_c_725_n N_VGND_c_1314_n 0.0227392f $X=6.83 $Y=0.7 $X2=0
+ $Y2=0
cc_559 N_A_865_111#_M1023_g N_VPWR_c_1131_n 0.0138266f $X=6.44 $Y=0.93 $X2=0
+ $Y2=0
cc_560 N_A_865_111#_c_790_n N_VPWR_c_1143_n 0.00158339f $X=4.465 $Y=2.905 $X2=0
+ $Y2=0
cc_561 N_A_865_111#_M1023_g N_VPWR_c_1143_n 0.0175835f $X=6.44 $Y=0.93 $X2=0
+ $Y2=0
cc_562 N_A_865_111#_c_787_n N_A_709_111#_c_1229_n 0.0107595f $X=4.465 $Y=0.775
+ $X2=0 $Y2=0
cc_563 N_A_865_111#_c_787_n N_A_709_111#_c_1223_n 0.00493683f $X=4.465 $Y=0.775
+ $X2=13.68 $Y2=0
cc_564 N_A_865_111#_M1023_g N_VGND_c_1306_n 0.00195592f $X=6.44 $Y=0.93 $X2=0
+ $Y2=0
cc_565 N_A_865_111#_c_787_n N_VGND_c_1314_n 0.0219009f $X=4.465 $Y=0.775 $X2=0
+ $Y2=0
cc_566 N_A_865_111#_M1023_g N_VGND_c_1314_n 0.0175795f $X=6.44 $Y=0.93 $X2=0
+ $Y2=0
cc_567 N_A_1711_85#_M1016_g N_A_1494_539#_M1009_g 0.0240079f $X=8.805 $Y=0.765
+ $X2=0 $Y2=0
cc_568 N_A_1711_85#_c_862_n N_A_1494_539#_M1009_g 0.0305575f $X=10.76 $Y=1.83
+ $X2=0 $Y2=0
cc_569 N_A_1711_85#_c_865_n N_A_1494_539#_M1009_g 0.0338301f $X=9.905 $Y=1.59
+ $X2=0 $Y2=0
cc_570 N_A_1711_85#_c_866_n N_A_1494_539#_M1009_g 0.027033f $X=10.07 $Y=0.7
+ $X2=0 $Y2=0
cc_571 N_A_1711_85#_c_893_p N_A_1494_539#_M1009_g 9.72163e-19 $X=8.94 $Y=1.655
+ $X2=0 $Y2=0
cc_572 N_A_1711_85#_c_868_n N_A_1494_539#_M1009_g 0.0161348f $X=8.94 $Y=1.655
+ $X2=0 $Y2=0
cc_573 N_A_1711_85#_c_869_n N_A_1494_539#_M1009_g 0.0114365f $X=10.07 $Y=1.74
+ $X2=0 $Y2=0
cc_574 N_A_1711_85#_M1008_g N_A_1494_539#_M1003_g 0.0142089f $X=8.805 $Y=2.905
+ $X2=0 $Y2=0
cc_575 N_A_1711_85#_c_879_n N_A_1494_539#_M1003_g 0.0335315f $X=10.07 $Y=2.84
+ $X2=0 $Y2=0
cc_576 N_A_1711_85#_M1016_g N_A_1494_539#_c_979_n 0.00428769f $X=8.805 $Y=0.765
+ $X2=0 $Y2=0
cc_577 N_A_1711_85#_M1016_g N_A_1494_539#_c_983_n 0.0220359f $X=8.805 $Y=0.765
+ $X2=0 $Y2=0
cc_578 N_A_1711_85#_M1008_g N_A_1494_539#_c_983_n 0.00718821f $X=8.805 $Y=2.905
+ $X2=0 $Y2=0
cc_579 N_A_1711_85#_c_893_p N_A_1494_539#_c_983_n 0.0443906f $X=8.94 $Y=1.655
+ $X2=0 $Y2=0
cc_580 N_A_1711_85#_c_868_n N_A_1494_539#_c_983_n 0.0207158f $X=8.94 $Y=1.655
+ $X2=0 $Y2=0
cc_581 N_A_1711_85#_M1008_g N_A_1494_539#_c_992_n 0.0278233f $X=8.805 $Y=2.905
+ $X2=0 $Y2=0
cc_582 N_A_1711_85#_c_865_n N_A_1494_539#_c_992_n 0.00838914f $X=9.905 $Y=1.59
+ $X2=0 $Y2=0
cc_583 N_A_1711_85#_c_879_n N_A_1494_539#_c_992_n 0.0129587f $X=10.07 $Y=2.84
+ $X2=0 $Y2=0
cc_584 N_A_1711_85#_c_893_p N_A_1494_539#_c_992_n 0.0239231f $X=8.94 $Y=1.655
+ $X2=0 $Y2=0
cc_585 N_A_1711_85#_c_868_n N_A_1494_539#_c_992_n 0.00201454f $X=8.94 $Y=1.655
+ $X2=0 $Y2=0
cc_586 N_A_1711_85#_M1008_g N_A_1494_539#_c_993_n 0.00209745f $X=8.805 $Y=2.905
+ $X2=0 $Y2=0
cc_587 N_A_1711_85#_M1008_g N_A_1494_539#_c_1047_n 9.65496e-19 $X=8.805 $Y=2.905
+ $X2=0 $Y2=0
cc_588 N_A_1711_85#_c_865_n N_A_1494_539#_c_1047_n 0.0238665f $X=9.905 $Y=1.59
+ $X2=0 $Y2=0
cc_589 N_A_1711_85#_c_879_n N_A_1494_539#_c_1047_n 0.0250172f $X=10.07 $Y=2.84
+ $X2=0 $Y2=0
cc_590 N_A_1711_85#_c_893_p N_A_1494_539#_c_1047_n 0.0141999f $X=8.94 $Y=1.655
+ $X2=0 $Y2=0
cc_591 N_A_1711_85#_c_868_n N_A_1494_539#_c_1047_n 0.00142444f $X=8.94 $Y=1.655
+ $X2=0 $Y2=0
cc_592 N_A_1711_85#_c_869_n N_A_1494_539#_c_1047_n 0.00905623f $X=10.07 $Y=1.74
+ $X2=0 $Y2=0
cc_593 N_A_1711_85#_M1008_g N_A_1494_539#_c_984_n 0.0171633f $X=8.805 $Y=2.905
+ $X2=0 $Y2=0
cc_594 N_A_1711_85#_c_865_n N_A_1494_539#_c_984_n 0.00161135f $X=9.905 $Y=1.59
+ $X2=0 $Y2=0
cc_595 N_A_1711_85#_c_879_n N_A_1494_539#_c_984_n 0.0227469f $X=10.07 $Y=2.84
+ $X2=0 $Y2=0
cc_596 N_A_1711_85#_c_893_p N_A_1494_539#_c_984_n 0.00141778f $X=8.94 $Y=1.655
+ $X2=0 $Y2=0
cc_597 N_A_1711_85#_c_868_n N_A_1494_539#_c_984_n 0.0199051f $X=8.94 $Y=1.655
+ $X2=0 $Y2=0
cc_598 N_A_1711_85#_c_869_n N_A_1494_539#_c_984_n 0.00535511f $X=10.07 $Y=1.74
+ $X2=0 $Y2=0
cc_599 N_A_1711_85#_M1005_g N_A_2365_443#_M1020_g 0.0184541f $X=12.34 $Y=2.59
+ $X2=0 $Y2=0
cc_600 N_A_1711_85#_M1014_g N_A_2365_443#_M1027_g 0.0145305f $X=12.36 $Y=1.235
+ $X2=0 $Y2=0
cc_601 N_A_1711_85#_M1001_g N_A_2365_443#_c_1084_n 0.00121637f $X=11.01 $Y=2.965
+ $X2=13.68 $Y2=0
cc_602 N_A_1711_85#_c_860_n N_A_2365_443#_c_1084_n 9.44109e-19 $X=12.09 $Y=1.83
+ $X2=13.68 $Y2=0
cc_603 N_A_1711_85#_M1005_g N_A_2365_443#_c_1084_n 0.0158627f $X=12.34 $Y=2.59
+ $X2=13.68 $Y2=0
cc_604 N_A_1711_85#_M1010_g N_A_2365_443#_c_1078_n 0.00353218f $X=11.01 $Y=1.07
+ $X2=6.96 $Y2=0
cc_605 N_A_1711_85#_c_860_n N_A_2365_443#_c_1078_n 0.0115591f $X=12.09 $Y=1.83
+ $X2=6.96 $Y2=0
cc_606 N_A_1711_85#_M1014_g N_A_2365_443#_c_1078_n 0.0162876f $X=12.36 $Y=1.235
+ $X2=6.96 $Y2=0
cc_607 N_A_1711_85#_c_864_n N_A_2365_443#_c_1078_n 0.00435507f $X=12.35 $Y=1.83
+ $X2=6.96 $Y2=0
cc_608 N_A_1711_85#_c_864_n N_A_2365_443#_c_1079_n 0.0441217f $X=12.35 $Y=1.83
+ $X2=0 $Y2=0
cc_609 N_A_1711_85#_c_864_n N_A_2365_443#_c_1080_n 0.0212641f $X=12.35 $Y=1.83
+ $X2=0 $Y2=0
cc_610 N_A_1711_85#_M1001_g N_A_2365_443#_c_1087_n 0.00310603f $X=11.01 $Y=2.965
+ $X2=0 $Y2=0
cc_611 N_A_1711_85#_c_860_n N_A_2365_443#_c_1087_n 0.0114226f $X=12.09 $Y=1.83
+ $X2=0 $Y2=0
cc_612 N_A_1711_85#_M1005_g N_A_2365_443#_c_1087_n 0.00662382f $X=12.34 $Y=2.59
+ $X2=0 $Y2=0
cc_613 N_A_1711_85#_c_864_n N_A_2365_443#_c_1087_n 0.00417344f $X=12.35 $Y=1.83
+ $X2=0 $Y2=0
cc_614 N_A_1711_85#_c_860_n N_A_2365_443#_c_1103_n 0.0259571f $X=12.09 $Y=1.83
+ $X2=0 $Y2=0
cc_615 N_A_1711_85#_c_864_n N_A_2365_443#_c_1103_n 0.00238473f $X=12.35 $Y=1.83
+ $X2=0 $Y2=0
cc_616 N_A_1711_85#_M1008_g N_VPWR_c_1134_n 0.0555024f $X=8.805 $Y=2.905 $X2=0
+ $Y2=0
cc_617 N_A_1711_85#_c_879_n N_VPWR_c_1134_n 0.0328768f $X=10.07 $Y=2.84 $X2=0
+ $Y2=0
cc_618 N_A_1711_85#_M1001_g N_VPWR_c_1137_n 0.0605836f $X=11.01 $Y=2.965 $X2=0
+ $Y2=0
cc_619 N_A_1711_85#_c_860_n N_VPWR_c_1137_n 0.0126213f $X=12.09 $Y=1.83 $X2=0
+ $Y2=0
cc_620 N_A_1711_85#_M1005_g N_VPWR_c_1137_n 0.00512254f $X=12.34 $Y=2.59 $X2=0
+ $Y2=0
cc_621 N_A_1711_85#_M1005_g N_VPWR_c_1140_n 0.0682053f $X=12.34 $Y=2.59 $X2=0
+ $Y2=0
cc_622 N_A_1711_85#_c_864_n N_VPWR_c_1140_n 6.03453e-19 $X=12.35 $Y=1.83 $X2=0
+ $Y2=0
cc_623 N_A_1711_85#_M1001_g N_VPWR_c_1143_n 0.0120207f $X=11.01 $Y=2.965 $X2=0
+ $Y2=0
cc_624 N_A_1711_85#_M1005_g N_VPWR_c_1143_n 0.00584154f $X=12.34 $Y=2.59 $X2=0
+ $Y2=0
cc_625 N_A_1711_85#_c_879_n N_VPWR_c_1143_n 0.0400422f $X=10.07 $Y=2.84 $X2=0
+ $Y2=0
cc_626 N_A_1711_85#_M1010_g Q 0.00762126f $X=11.01 $Y=1.07 $X2=0 $Y2=0
cc_627 N_A_1711_85#_M1001_g Q 0.00824262f $X=11.01 $Y=2.965 $X2=0 $Y2=0
cc_628 N_A_1711_85#_c_862_n Q 0.0160592f $X=10.76 $Y=1.83 $X2=0 $Y2=0
cc_629 N_A_1711_85#_c_863_n Q 0.0292466f $X=11.01 $Y=1.83 $X2=0 $Y2=0
cc_630 N_A_1711_85#_c_879_n Q 0.00606278f $X=10.07 $Y=2.84 $X2=0 $Y2=0
cc_631 N_A_1711_85#_c_869_n Q 0.029151f $X=10.07 $Y=1.74 $X2=0 $Y2=0
cc_632 N_A_1711_85#_M1001_g Q 0.035316f $X=11.01 $Y=2.965 $X2=0.24 $Y2=0
cc_633 N_A_1711_85#_M1010_g N_Q_c_1256_n 0.0191296f $X=11.01 $Y=1.07 $X2=0 $Y2=0
cc_634 N_A_1711_85#_c_866_n N_Q_c_1256_n 0.0560601f $X=10.07 $Y=0.7 $X2=0 $Y2=0
cc_635 N_A_1711_85#_M1010_g Q 0.00618786f $X=11.01 $Y=1.07 $X2=0 $Y2=0
cc_636 N_A_1711_85#_c_862_n Q 0.0102906f $X=10.76 $Y=1.83 $X2=0 $Y2=0
cc_637 N_A_1711_85#_c_869_n Q 0.00397605f $X=10.07 $Y=1.74 $X2=0 $Y2=0
cc_638 N_A_1711_85#_M1001_g N_Q_c_1262_n 0.00618786f $X=11.01 $Y=2.965 $X2=0
+ $Y2=0
cc_639 N_A_1711_85#_c_862_n N_Q_c_1262_n 0.0103264f $X=10.76 $Y=1.83 $X2=0 $Y2=0
cc_640 N_A_1711_85#_c_879_n N_Q_c_1262_n 0.103887f $X=10.07 $Y=2.84 $X2=0 $Y2=0
cc_641 N_A_1711_85#_c_869_n N_Q_c_1262_n 0.00341927f $X=10.07 $Y=1.74 $X2=0
+ $Y2=0
cc_642 N_A_1711_85#_M1016_g N_VGND_c_1308_n 0.0580449f $X=8.805 $Y=0.765 $X2=0
+ $Y2=0
cc_643 N_A_1711_85#_c_865_n N_VGND_c_1308_n 0.0476367f $X=9.905 $Y=1.59 $X2=0
+ $Y2=0
cc_644 N_A_1711_85#_c_866_n N_VGND_c_1308_n 0.0586492f $X=10.07 $Y=0.7 $X2=0
+ $Y2=0
cc_645 N_A_1711_85#_c_893_p N_VGND_c_1308_n 0.0266932f $X=8.94 $Y=1.655 $X2=0
+ $Y2=0
cc_646 N_A_1711_85#_c_868_n N_VGND_c_1308_n 0.00197001f $X=8.94 $Y=1.655 $X2=0
+ $Y2=0
cc_647 N_A_1711_85#_M1010_g N_VGND_c_1310_n 0.0510701f $X=11.01 $Y=1.07 $X2=0
+ $Y2=0
cc_648 N_A_1711_85#_c_860_n N_VGND_c_1310_n 0.013916f $X=12.09 $Y=1.83 $X2=0
+ $Y2=0
cc_649 N_A_1711_85#_M1014_g N_VGND_c_1310_n 0.00457714f $X=12.36 $Y=1.235 $X2=0
+ $Y2=0
cc_650 N_A_1711_85#_M1014_g N_VGND_c_1312_n 0.0487781f $X=12.36 $Y=1.235 $X2=0
+ $Y2=0
cc_651 N_A_1711_85#_M1016_g N_VGND_c_1314_n 0.0109908f $X=8.805 $Y=0.765 $X2=0
+ $Y2=0
cc_652 N_A_1711_85#_M1010_g N_VGND_c_1314_n 0.0147965f $X=11.01 $Y=1.07 $X2=0
+ $Y2=0
cc_653 N_A_1711_85#_M1014_g N_VGND_c_1314_n 0.00612244f $X=12.36 $Y=1.235 $X2=0
+ $Y2=0
cc_654 N_A_1711_85#_c_866_n N_VGND_c_1314_n 0.0317391f $X=10.07 $Y=0.7 $X2=0
+ $Y2=0
cc_655 N_A_1494_539#_M1003_g N_VPWR_c_1134_n 0.027156f $X=9.68 $Y=3.195 $X2=0
+ $Y2=0
cc_656 N_A_1494_539#_c_992_n N_VPWR_c_1134_n 0.0658013f $X=9.395 $Y=2.41 $X2=0
+ $Y2=0
cc_657 N_A_1494_539#_c_993_n N_VPWR_c_1134_n 0.00759982f $X=8.595 $Y=2.41 $X2=0
+ $Y2=0
cc_658 N_A_1494_539#_c_984_n N_VPWR_c_1134_n 0.00161905f $X=9.56 $Y=2.005 $X2=0
+ $Y2=0
cc_659 N_A_1494_539#_M1003_g N_VPWR_c_1143_n 0.0289411f $X=9.68 $Y=3.195 $X2=0
+ $Y2=0
cc_660 N_A_1494_539#_c_990_n N_VPWR_c_1143_n 0.024174f $X=7.61 $Y=3.37 $X2=0
+ $Y2=0
cc_661 N_A_1494_539#_M1003_g Q 0.00215212f $X=9.68 $Y=3.195 $X2=0.24 $Y2=0
cc_662 N_A_1494_539#_M1009_g N_Q_c_1256_n 0.00192078f $X=9.68 $Y=0.93 $X2=0
+ $Y2=0
cc_663 N_A_1494_539#_c_984_n N_Q_c_1262_n 0.00182116f $X=9.56 $Y=2.005 $X2=0
+ $Y2=0
cc_664 N_A_1494_539#_M1009_g N_VGND_c_1308_n 0.0504437f $X=9.68 $Y=0.93 $X2=0
+ $Y2=0
cc_665 N_A_1494_539#_c_979_n N_VGND_c_1308_n 0.0116452f $X=8.425 $Y=0.6 $X2=0
+ $Y2=0
cc_666 N_A_1494_539#_c_983_n N_VGND_c_1308_n 0.0463156f $X=8.51 $Y=2.325 $X2=0
+ $Y2=0
cc_667 N_A_1494_539#_M1009_g N_VGND_c_1314_n 0.0122927f $X=9.68 $Y=0.93 $X2=0
+ $Y2=0
cc_668 N_A_1494_539#_c_979_n N_VGND_c_1314_n 0.0536722f $X=8.425 $Y=0.6 $X2=0
+ $Y2=0
cc_669 N_A_1494_539#_c_981_n N_VGND_c_1314_n 0.0225267f $X=7.795 $Y=0.6 $X2=0
+ $Y2=0
cc_670 N_A_1494_539#_c_979_n A_1669_111# 8.39422e-19 $X=8.425 $Y=0.6 $X2=0 $Y2=0
cc_671 N_A_1494_539#_c_983_n A_1669_111# 0.00382391f $X=8.51 $Y=2.325 $X2=0
+ $Y2=0
cc_672 N_A_2365_443#_c_1084_n N_VPWR_c_1137_n 0.0655371f $X=11.95 $Y=2.36 $X2=0
+ $Y2=0
cc_673 N_A_2365_443#_M1020_g N_VPWR_c_1140_n 0.0702557f $X=13.235 $Y=2.965 $X2=0
+ $Y2=0
cc_674 N_A_2365_443#_c_1079_n N_VPWR_c_1140_n 0.0754782f $X=13.135 $Y=1.83 $X2=0
+ $Y2=0
cc_675 N_A_2365_443#_c_1080_n N_VPWR_c_1140_n 9.86162e-19 $X=13.135 $Y=1.83
+ $X2=0 $Y2=0
cc_676 N_A_2365_443#_c_1087_n N_VPWR_c_1140_n 0.0613912f $X=11.95 $Y=2.195 $X2=0
+ $Y2=0
cc_677 N_A_2365_443#_M1020_g N_VPWR_c_1143_n 0.0130327f $X=13.235 $Y=2.965 $X2=0
+ $Y2=0
cc_678 N_A_2365_443#_c_1084_n N_VPWR_c_1143_n 0.0141253f $X=11.95 $Y=2.36 $X2=0
+ $Y2=0
cc_679 N_A_2365_443#_M1020_g Q_N 0.00579133f $X=13.235 $Y=2.965 $X2=0 $Y2=0
cc_680 N_A_2365_443#_M1027_g Q_N 0.0236277f $X=13.255 $Y=1.07 $X2=0 $Y2=0
cc_681 N_A_2365_443#_c_1079_n Q_N 0.0250026f $X=13.135 $Y=1.83 $X2=0 $Y2=0
cc_682 N_A_2365_443#_c_1080_n Q_N 0.0249251f $X=13.135 $Y=1.83 $X2=0 $Y2=0
cc_683 N_A_2365_443#_M1020_g Q_N 0.00496571f $X=13.235 $Y=2.965 $X2=0.24 $Y2=0
cc_684 N_A_2365_443#_M1020_g Q_N 0.0260206f $X=13.235 $Y=2.965 $X2=0 $Y2=0
cc_685 N_A_2365_443#_c_1078_n N_VGND_c_1310_n 0.0399591f $X=11.97 $Y=1.235 $X2=0
+ $Y2=0
cc_686 N_A_2365_443#_M1027_g N_VGND_c_1312_n 0.0532767f $X=13.255 $Y=1.07 $X2=0
+ $Y2=0
cc_687 N_A_2365_443#_c_1078_n N_VGND_c_1312_n 0.0364263f $X=11.97 $Y=1.235 $X2=0
+ $Y2=0
cc_688 N_A_2365_443#_c_1079_n N_VGND_c_1312_n 0.0754782f $X=13.135 $Y=1.83 $X2=0
+ $Y2=0
cc_689 N_A_2365_443#_c_1080_n N_VGND_c_1312_n 0.00158962f $X=13.135 $Y=1.83
+ $X2=0 $Y2=0
cc_690 N_A_2365_443#_M1027_g N_VGND_c_1314_n 0.0141765f $X=13.255 $Y=1.07 $X2=0
+ $Y2=0
cc_691 N_A_2365_443#_c_1078_n N_VGND_c_1314_n 0.0152237f $X=11.97 $Y=1.235 $X2=0
+ $Y2=0
cc_692 N_VPWR_c_1143_n N_A_709_111#_c_1225_n 0.00151101f $X=13.13 $Y=3.59 $X2=0
+ $Y2=0
cc_693 N_VPWR_c_1143_n Q 0.0488721f $X=13.13 $Y=3.59 $X2=0 $Y2=0
cc_694 N_VPWR_c_1137_n N_Q_c_1262_n 0.112748f $X=11.4 $Y=2.36 $X2=0 $Y2=0
cc_695 N_VPWR_c_1140_n Q_N 0.0995832f $X=12.845 $Y=2.34 $X2=0 $Y2=0
cc_696 N_VPWR_c_1143_n Q_N 0.0451876f $X=13.13 $Y=3.59 $X2=0 $Y2=0
cc_697 N_A_709_111#_c_1229_n N_VGND_c_1314_n 0.020053f $X=3.685 $Y=0.775 $X2=0
+ $Y2=0
cc_698 N_Q_c_1256_n N_VGND_c_1310_n 0.0616937f $X=10.62 $Y=0.84 $X2=0 $Y2=0
cc_699 N_Q_c_1256_n N_VGND_c_1314_n 0.0185753f $X=10.62 $Y=0.84 $X2=0 $Y2=0
cc_700 Q_N N_VGND_c_1312_n 0.0533341f $X=13.595 $Y=0.84 $X2=0 $Y2=0
cc_701 Q_N N_VGND_c_1314_n 0.0144846f $X=13.595 $Y=0.84 $X2=0 $Y2=0
cc_702 N_VGND_c_1306_n A_1021_111# 0.00359873f $X=6.05 $Y=0.8 $X2=0 $Y2=0
cc_703 N_VGND_c_1314_n A_1021_111# 0.00333633f $X=13.15 $Y=0.48 $X2=0 $Y2=0
