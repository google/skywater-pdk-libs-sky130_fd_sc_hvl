# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hvl__sdlclkp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN GATE
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 1.535000 1.805000 2.125000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.590000 0.515000 10.955000 1.215000 ;
        RECT 10.590000 1.895000 10.955000 3.735000 ;
        RECT 10.685000 1.215000 10.955000 1.895000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 1.535000 0.925000 2.125000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  1.170000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.320000 1.465000 4.650000 1.975000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 11.040000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 11.040000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 11.040000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 11.040000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 11.040000 0.085000 ;
      RECT 0.000000  3.985000 11.040000 4.155000 ;
      RECT 0.290000  0.840000  0.620000 1.195000 ;
      RECT 0.290000  1.195000  2.145000 1.365000 ;
      RECT 0.290000  2.295000  0.620000 3.445000 ;
      RECT 0.290000  3.445000  1.985000 3.615000 ;
      RECT 0.290000  3.615000  4.290000 3.815000 ;
      RECT 0.730000  0.365000  1.740000 0.625000 ;
      RECT 1.070000  0.625000  1.400000 1.025000 ;
      RECT 1.850000  0.840000  2.145000 1.195000 ;
      RECT 1.850000  2.295000  2.145000 3.055000 ;
      RECT 1.975000  1.365000  2.145000 2.295000 ;
      RECT 2.115000  0.365000  3.770000 0.535000 ;
      RECT 2.115000  0.535000  2.825000 0.670000 ;
      RECT 2.155000  3.225000  3.455000 3.445000 ;
      RECT 2.555000  1.555000  3.065000 1.885000 ;
      RECT 2.630000  0.840000  2.960000 1.555000 ;
      RECT 2.630000  1.885000  2.960000 3.055000 ;
      RECT 3.180000  0.705000  3.430000 1.080000 ;
      RECT 3.235000  1.080000  3.430000 2.145000 ;
      RECT 3.235000  2.145000  4.650000 2.315000 ;
      RECT 3.235000  2.315000  3.455000 3.225000 ;
      RECT 3.600000  0.535000  3.770000 1.125000 ;
      RECT 3.600000  1.125000  5.030000 1.295000 ;
      RECT 3.600000  1.295000  3.930000 1.965000 ;
      RECT 3.625000  3.445000  4.290000 3.615000 ;
      RECT 3.940000  0.255000  4.885000 0.535000 ;
      RECT 3.940000  0.535000  4.610000 0.625000 ;
      RECT 3.940000  0.625000  4.290000 0.955000 ;
      RECT 3.960000  2.485000  4.290000 3.445000 ;
      RECT 4.480000  2.315000  4.650000 3.385000 ;
      RECT 4.480000  3.385000  6.475000 3.555000 ;
      RECT 4.780000  0.705000  5.030000 1.125000 ;
      RECT 4.820000  1.295000  5.030000 3.005000 ;
      RECT 4.820000  3.005000  6.135000 3.215000 ;
      RECT 5.055000  0.255000  5.620000 0.535000 ;
      RECT 5.335000  0.535000  5.620000 1.195000 ;
      RECT 5.335000  1.195000  7.450000 1.365000 ;
      RECT 5.335000  1.365000  5.505000 2.330000 ;
      RECT 5.335000  2.330000  5.620000 2.660000 ;
      RECT 5.675000  1.615000  6.265000 1.945000 ;
      RECT 5.790000  0.255000  7.110000 0.625000 ;
      RECT 6.095000  1.945000  6.265000 2.425000 ;
      RECT 6.095000  2.425000  6.475000 2.595000 ;
      RECT 6.305000  2.595000  6.475000 3.385000 ;
      RECT 6.475000  1.535000  6.805000 1.875000 ;
      RECT 6.475000  1.875000  7.890000 2.085000 ;
      RECT 6.645000  3.445000  9.025000 3.615000 ;
      RECT 6.645000  3.615000 10.420000 3.815000 ;
      RECT 6.780000  0.625000  7.110000 1.025000 ;
      RECT 6.780000  2.330000  7.110000 3.445000 ;
      RECT 7.085000  1.365000  7.450000 1.655000 ;
      RECT 7.280000  0.355000  7.870000 0.670000 ;
      RECT 7.280000  0.670000  7.450000 1.195000 ;
      RECT 7.620000  0.840000  7.890000 1.615000 ;
      RECT 7.620000  1.615000  8.745000 1.825000 ;
      RECT 7.620000  1.825000  7.890000 1.875000 ;
      RECT 7.620000  2.085000  7.890000 2.660000 ;
      RECT 8.040000  0.255000 10.420000 0.625000 ;
      RECT 8.110000  0.885000  9.140000 1.215000 ;
      RECT 8.110000  2.225000  8.440000 3.445000 ;
      RECT 8.415000  1.385000  8.745000 1.615000 ;
      RECT 8.415000  1.825000  8.745000 2.055000 ;
      RECT 8.915000  1.215000  9.140000 1.385000 ;
      RECT 8.915000  1.385000 10.515000 1.555000 ;
      RECT 8.915000  1.555000  9.140000 2.955000 ;
      RECT 9.195000  3.125000  9.560000 3.445000 ;
      RECT 9.310000  1.725000  9.640000 2.025000 ;
      RECT 9.310000  2.025000  9.560000 3.125000 ;
      RECT 9.730000  0.625000 10.060000 1.215000 ;
      RECT 9.730000  2.195000 10.060000 3.445000 ;
      RECT 9.730000  3.445000 10.420000 3.615000 ;
      RECT 9.905000  1.555000 10.515000 1.725000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.380000  3.475000  0.550000 3.645000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.740000  3.475000  0.910000 3.645000 ;
      RECT  0.790000  0.425000  0.960000 0.595000 ;
      RECT  1.100000  3.475000  1.270000 3.645000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.150000  0.425000  1.320000 0.595000 ;
      RECT  1.460000  3.475000  1.630000 3.645000 ;
      RECT  1.510000  0.425000  1.680000 0.595000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  1.820000  3.615000  1.990000 3.785000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.180000  3.615000  2.350000 3.785000 ;
      RECT  2.540000  3.615000  2.710000 3.785000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.955000  3.615000  3.125000 3.785000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.315000  3.615000  3.485000 3.785000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.675000  3.475000  3.845000 3.645000 ;
      RECT  3.955000  0.425000  4.125000 0.595000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.035000  3.475000  4.205000 3.645000 ;
      RECT  4.315000  0.425000  4.485000 0.595000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.675000  0.355000  4.845000 0.525000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.830000  0.355000  6.000000 0.525000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.190000  0.355000  6.360000 0.525000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.550000  0.425000  6.720000 0.595000 ;
      RECT  6.675000  3.475000  6.845000 3.645000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  6.910000  0.425000  7.080000 0.595000 ;
      RECT  7.035000  3.475000  7.205000 3.645000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.395000  3.545000  7.565000 3.715000 ;
      RECT  7.755000  3.545000  7.925000 3.715000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.060000  0.355000  8.230000 0.525000 ;
      RECT  8.115000  3.475000  8.285000 3.645000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.420000  0.355000  8.590000 0.525000 ;
      RECT  8.475000  3.475000  8.645000 3.645000 ;
      RECT  8.780000  0.355000  8.950000 0.525000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.140000  0.355000  9.310000 0.525000 ;
      RECT  9.155000  3.615000  9.325000 3.785000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.500000  0.425000  9.670000 0.595000 ;
      RECT  9.515000  3.615000  9.685000 3.785000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.860000  0.425000 10.030000 0.595000 ;
      RECT  9.875000  3.475000 10.045000 3.645000 ;
      RECT 10.220000  0.425000 10.390000 0.595000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.475000 10.405000 3.645000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
  END
END sky130_fd_sc_hvl__sdlclkp_1
