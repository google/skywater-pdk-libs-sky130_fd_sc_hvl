* File: sky130_fd_sc_hvl__dlrtp_1.pxi.spice
* Created: Wed Sep  2 09:05:56 2020
* 
x_PM_SKY130_FD_SC_HVL__DLRTP_1%VNB N_VNB_M1019_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__DLRTP_1%VNB
x_PM_SKY130_FD_SC_HVL__DLRTP_1%VPB N_VPB_M1014_b VPB N_VPB_c_74_p VPB
+ PM_SKY130_FD_SC_HVL__DLRTP_1%VPB
x_PM_SKY130_FD_SC_HVL__DLRTP_1%D D D N_D_M1019_g N_D_M1014_g
+ PM_SKY130_FD_SC_HVL__DLRTP_1%D
x_PM_SKY130_FD_SC_HVL__DLRTP_1%GATE GATE GATE GATE N_GATE_M1007_g N_GATE_M1005_g
+ PM_SKY130_FD_SC_HVL__DLRTP_1%GATE
x_PM_SKY130_FD_SC_HVL__DLRTP_1%A_345_107# N_A_345_107#_M1007_d
+ N_A_345_107#_M1005_d N_A_345_107#_c_187_n N_A_345_107#_c_188_n
+ N_A_345_107#_M1004_g N_A_345_107#_c_200_n N_A_345_107#_c_191_n
+ N_A_345_107#_c_203_n N_A_345_107#_c_204_n N_A_345_107#_c_192_n
+ N_A_345_107#_c_193_n N_A_345_107#_c_194_n N_A_345_107#_c_196_n
+ N_A_345_107#_c_197_n N_A_345_107#_M1018_g N_A_345_107#_M1001_g
+ N_A_345_107#_M1016_g PM_SKY130_FD_SC_HVL__DLRTP_1%A_345_107#
x_PM_SKY130_FD_SC_HVL__DLRTP_1%A_32_107# N_A_32_107#_M1019_s N_A_32_107#_M1014_s
+ N_A_32_107#_M1008_g N_A_32_107#_M1010_g N_A_32_107#_c_301_n
+ N_A_32_107#_c_303_n N_A_32_107#_c_304_n N_A_32_107#_c_305_n
+ N_A_32_107#_c_306_n N_A_32_107#_c_307_n N_A_32_107#_c_308_n
+ PM_SKY130_FD_SC_HVL__DLRTP_1%A_32_107#
x_PM_SKY130_FD_SC_HVL__DLRTP_1%A_462_107# N_A_462_107#_M1018_s
+ N_A_462_107#_M1001_s N_A_462_107#_M1006_g N_A_462_107#_c_372_n
+ N_A_462_107#_c_364_n N_A_462_107#_c_366_n N_A_462_107#_c_367_n
+ N_A_462_107#_c_373_n N_A_462_107#_c_374_n N_A_462_107#_c_368_n
+ N_A_462_107#_c_369_n N_A_462_107#_c_376_n N_A_462_107#_c_377_n
+ N_A_462_107#_M1012_g N_A_462_107#_c_378_n
+ PM_SKY130_FD_SC_HVL__DLRTP_1%A_462_107#
x_PM_SKY130_FD_SC_HVL__DLRTP_1%A_1138_81# N_A_1138_81#_M1000_s
+ N_A_1138_81#_M1011_d N_A_1138_81#_c_470_n N_A_1138_81#_M1017_g
+ N_A_1138_81#_M1015_g N_A_1138_81#_c_479_n N_A_1138_81#_c_473_n
+ N_A_1138_81#_c_493_p N_A_1138_81#_c_465_n N_A_1138_81#_c_474_n
+ N_A_1138_81#_c_475_n N_A_1138_81#_c_476_n N_A_1138_81#_c_466_n
+ N_A_1138_81#_c_516_p N_A_1138_81#_M1009_g N_A_1138_81#_M1013_g
+ N_A_1138_81#_c_469_n PM_SKY130_FD_SC_HVL__DLRTP_1%A_1138_81#
x_PM_SKY130_FD_SC_HVL__DLRTP_1%A_917_107# N_A_917_107#_M1012_d
+ N_A_917_107#_M1016_d N_A_917_107#_M1011_g N_A_917_107#_c_555_n
+ N_A_917_107#_M1000_g N_A_917_107#_c_566_n N_A_917_107#_c_567_n
+ N_A_917_107#_c_570_n N_A_917_107#_c_557_n N_A_917_107#_c_572_n
+ N_A_917_107#_c_558_n N_A_917_107#_c_559_n N_A_917_107#_c_560_n
+ N_A_917_107#_c_561_n N_A_917_107#_c_563_n N_A_917_107#_c_621_n
+ N_A_917_107#_c_564_n PM_SKY130_FD_SC_HVL__DLRTP_1%A_917_107#
x_PM_SKY130_FD_SC_HVL__DLRTP_1%RESET_B RESET_B RESET_B RESET_B N_RESET_B_c_661_n
+ N_RESET_B_M1002_g N_RESET_B_M1003_g PM_SKY130_FD_SC_HVL__DLRTP_1%RESET_B
x_PM_SKY130_FD_SC_HVL__DLRTP_1%VPWR N_VPWR_M1014_d N_VPWR_M1001_d N_VPWR_M1013_d
+ N_VPWR_M1002_d VPWR N_VPWR_c_694_n N_VPWR_c_697_n N_VPWR_c_700_n
+ N_VPWR_c_703_n N_VPWR_c_706_n PM_SKY130_FD_SC_HVL__DLRTP_1%VPWR
x_PM_SKY130_FD_SC_HVL__DLRTP_1%Q N_Q_M1015_d N_Q_M1017_d Q Q Q Q Q Q Q
+ N_Q_c_755_n N_Q_c_761_n PM_SKY130_FD_SC_HVL__DLRTP_1%Q
x_PM_SKY130_FD_SC_HVL__DLRTP_1%VGND N_VGND_M1019_d N_VGND_M1018_d N_VGND_M1009_d
+ N_VGND_M1003_d VGND N_VGND_c_774_n N_VGND_c_776_n N_VGND_c_778_n
+ N_VGND_c_780_n N_VGND_c_782_n PM_SKY130_FD_SC_HVL__DLRTP_1%VGND
cc_1 N_VNB_M1019_b N_D_M1019_g 0.120745f $X=-0.33 $Y=-0.265 $X2=0.695 $Y2=0.745
cc_2 N_VNB_c_2_p N_D_M1019_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.695 $Y2=0.745
cc_3 N_VNB_M1019_b GATE 0.00851108f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_4 N_VNB_M1019_b N_GATE_M1007_g 0.128119f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=2.095
cc_5 N_VNB_c_2_p N_GATE_M1007_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.695 $Y2=2.095
cc_6 N_VNB_M1019_b N_A_345_107#_c_187_n 0.0438159f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_7 N_VNB_M1019_b N_A_345_107#_c_188_n 0.0155806f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=2.095
cc_8 N_VNB_M1019_b N_A_345_107#_M1004_g 0.0936111f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=3.195
cc_9 N_VNB_c_2_p N_A_345_107#_M1004_g 0.0023273f $X=0.24 $Y=0 $X2=0.695
+ $Y2=3.195
cc_10 N_VNB_M1019_b N_A_345_107#_c_191_n 0.00860932f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1019_b N_A_345_107#_c_192_n 0.020264f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1019_b N_A_345_107#_c_193_n 0.00431015f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1019_b N_A_345_107#_c_194_n 0.0296936f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_c_2_p N_A_345_107#_c_194_n 0.0010966f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_15 N_VNB_M1019_b N_A_345_107#_c_196_n 0.00880816f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_16 N_VNB_M1019_b N_A_345_107#_c_197_n 0.0112468f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_17 N_VNB_M1019_b N_A_345_107#_M1018_g 0.129681f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_c_2_p N_A_345_107#_M1018_g 9.58849e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_19 N_VNB_M1019_b N_A_32_107#_M1008_g 0.0707076f $X=-0.33 $Y=-0.265 $X2=0.735
+ $Y2=2.095
cc_20 N_VNB_c_2_p N_A_32_107#_M1008_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.735
+ $Y2=2.095
cc_21 N_VNB_M1019_b N_A_32_107#_c_301_n 0.0555095f $X=-0.33 $Y=-0.265 $X2=0.735
+ $Y2=2.405
cc_22 N_VNB_c_2_p N_A_32_107#_c_301_n 5.81195e-19 $X=0.24 $Y=0 $X2=0.735
+ $Y2=2.405
cc_23 N_VNB_M1019_b N_A_32_107#_c_303_n 0.0067175f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_24 N_VNB_M1019_b N_A_32_107#_c_304_n 0.0159515f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_25 N_VNB_M1019_b N_A_32_107#_c_305_n 0.0268928f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_26 N_VNB_M1019_b N_A_32_107#_c_306_n 0.0420231f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_27 N_VNB_M1019_b N_A_32_107#_c_307_n 0.00770964f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_28 N_VNB_M1019_b N_A_32_107#_c_308_n 0.0050765f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_29 N_VNB_M1019_b N_A_462_107#_c_364_n 0.00885801f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_30 N_VNB_c_2_p N_A_462_107#_c_364_n 6.32411e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_31 N_VNB_M1019_b N_A_462_107#_c_366_n 0.00988001f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_32 N_VNB_M1019_b N_A_462_107#_c_367_n 0.00387481f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_33 N_VNB_M1019_b N_A_462_107#_c_368_n 0.00810768f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_M1019_b N_A_462_107#_c_369_n 0.00771145f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_35 N_VNB_M1019_b N_A_462_107#_M1012_g 0.0839084f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_36 N_VNB_c_2_p N_A_462_107#_M1012_g 0.0023273f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_37 N_VNB_M1019_b N_A_1138_81#_M1015_g 0.0715731f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=3.195
cc_38 N_VNB_c_2_p N_A_1138_81#_M1015_g 0.00128467f $X=0.24 $Y=0 $X2=0.695
+ $Y2=3.195
cc_39 N_VNB_M1019_b N_A_1138_81#_c_465_n 0.0074163f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_M1019_b N_A_1138_81#_c_466_n 0.0186607f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_41 N_VNB_c_2_p N_A_1138_81#_c_466_n 0.00102439f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_42 N_VNB_M1019_b N_A_1138_81#_M1009_g 0.112286f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_M1019_b N_A_1138_81#_c_469_n 0.0537087f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_44 N_VNB_M1019_b N_A_917_107#_M1011_g 0.00713544f $X=-0.33 $Y=-0.265
+ $X2=0.735 $Y2=2.095
cc_45 N_VNB_M1019_b N_A_917_107#_c_555_n 0.0503298f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=3.195
cc_46 N_VNB_c_2_p N_A_917_107#_c_555_n 0.0023273f $X=0.24 $Y=0 $X2=0.695
+ $Y2=3.195
cc_47 N_VNB_M1019_b N_A_917_107#_c_557_n 0.00177939f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_M1019_b N_A_917_107#_c_558_n 0.00148236f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_49 N_VNB_M1019_b N_A_917_107#_c_559_n 0.00628447f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_M1019_b N_A_917_107#_c_560_n 0.0130208f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_51 N_VNB_M1019_b N_A_917_107#_c_561_n 0.0194072f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_52 N_VNB_c_2_p N_A_917_107#_c_561_n 0.00138851f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_53 N_VNB_M1019_b N_A_917_107#_c_563_n 8.82068e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_54 N_VNB_M1019_b N_A_917_107#_c_564_n 0.129493f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_55 N_VNB_M1019_b RESET_B 0.0020581f $X=-0.33 $Y=-0.265 $X2=0.635 $Y2=1.95
cc_56 N_VNB_M1019_b RESET_B 0.00790662f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_57 N_VNB_M1019_b N_RESET_B_c_661_n 0.0358811f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=2.095
cc_58 N_VNB_M1019_b N_RESET_B_M1003_g 0.0907482f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_59 N_VNB_c_2_p N_RESET_B_M1003_g 0.0023273f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_60 N_VNB_M1019_b N_Q_c_755_n 0.063857f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_61 N_VNB_c_2_p N_Q_c_755_n 8.31735e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_62 N_VNB_M1019_b N_VGND_c_774_n 0.0496364f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_63 N_VNB_c_2_p N_VGND_c_774_n 0.00269373f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_64 N_VNB_M1019_b N_VGND_c_776_n 0.0466961f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_65 N_VNB_c_2_p N_VGND_c_776_n 0.0027102f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_66 N_VNB_M1019_b N_VGND_c_778_n 0.0590394f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_67 N_VNB_c_2_p N_VGND_c_778_n 0.00269545f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_68 N_VNB_M1019_b N_VGND_c_780_n 0.0389793f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_69 N_VNB_c_2_p N_VGND_c_780_n 0.00166879f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_70 N_VNB_M1019_b N_VGND_c_782_n 0.147611f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_71 N_VNB_c_2_p N_VGND_c_782_n 1.02698f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_72 N_VPB_M1014_b N_D_M1019_g 0.118301f $X=-0.33 $Y=1.885 $X2=0.695 $Y2=0.745
cc_73 VPB N_D_M1019_g 6.11586e-19 $X=0 $Y=3.955 $X2=0.695 $Y2=0.745
cc_74 N_VPB_c_74_p N_D_M1019_g 0.00512296f $X=9.36 $Y=4.07 $X2=0.695 $Y2=0.745
cc_75 N_VPB_M1014_b N_GATE_M1007_g 0.126026f $X=-0.33 $Y=1.885 $X2=0.695
+ $Y2=2.095
cc_76 VPB N_GATE_M1007_g 9.99895e-19 $X=0 $Y=3.955 $X2=0.695 $Y2=2.095
cc_77 N_VPB_c_74_p N_GATE_M1007_g 0.00643888f $X=9.36 $Y=4.07 $X2=0.695
+ $Y2=2.095
cc_78 N_VPB_M1014_b N_A_345_107#_c_200_n 0.0232635f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_79 VPB N_A_345_107#_c_200_n 8.58775e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_80 N_VPB_c_74_p N_A_345_107#_c_200_n 0.0101785f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_81 N_VPB_M1014_b N_A_345_107#_c_203_n 0.0244201f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_82 N_VPB_M1014_b N_A_345_107#_c_204_n 0.00369566f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_83 N_VPB_M1014_b N_A_345_107#_c_196_n 0.002009f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_84 N_VPB_M1014_b N_A_345_107#_c_197_n 0.0812515f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_85 N_VPB_c_74_p N_A_345_107#_c_197_n 0.0102891f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_86 N_VPB_M1014_b N_A_345_107#_M1018_g 0.0888906f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_87 N_VPB_c_74_p N_A_345_107#_M1018_g 0.00499334f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_88 N_VPB_M1014_b N_A_32_107#_M1010_g 0.0678723f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_89 N_VPB_c_74_p N_A_32_107#_M1010_g 0.0035523f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_90 N_VPB_M1014_b N_A_32_107#_c_303_n 0.0756926f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_91 VPB N_A_32_107#_c_303_n 6.11207e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_92 N_VPB_c_74_p N_A_32_107#_c_303_n 0.00776898f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_93 N_VPB_M1014_b N_A_32_107#_c_306_n 0.00695392f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_94 N_VPB_M1014_b N_A_462_107#_c_372_n 0.0107675f $X=-0.33 $Y=1.885 $X2=0.695
+ $Y2=3.195
cc_95 N_VPB_M1014_b N_A_462_107#_c_373_n 0.00483489f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_96 N_VPB_M1014_b N_A_462_107#_c_374_n 0.00484175f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_97 N_VPB_M1014_b N_A_462_107#_c_368_n 0.00171633f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_98 N_VPB_M1014_b N_A_462_107#_c_376_n 0.00946936f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_99 N_VPB_M1014_b N_A_462_107#_c_377_n 0.0472953f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_100 N_VPB_M1014_b N_A_462_107#_c_378_n 0.0416988f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_101 N_VPB_M1014_b N_A_1138_81#_c_470_n 0.0401266f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_102 VPB N_A_1138_81#_c_470_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_103 N_VPB_c_74_p N_A_1138_81#_c_470_n 0.0162989f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_104 N_VPB_M1014_b N_A_1138_81#_c_473_n 0.00856641f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_105 N_VPB_M1014_b N_A_1138_81#_c_474_n 0.00557903f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_106 N_VPB_M1014_b N_A_1138_81#_c_475_n 0.00491892f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_107 N_VPB_M1014_b N_A_1138_81#_c_476_n 0.00815367f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_108 N_VPB_M1014_b N_A_1138_81#_M1009_g 0.0774285f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_109 N_VPB_M1014_b N_A_1138_81#_c_469_n 0.0424929f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_110 N_VPB_M1014_b N_A_917_107#_M1011_g 0.0603771f $X=-0.33 $Y=1.885 $X2=0.735
+ $Y2=2.095
cc_111 N_VPB_M1014_b N_A_917_107#_c_566_n 0.0142605f $X=-0.33 $Y=1.885 $X2=0.735
+ $Y2=2.035
cc_112 N_VPB_M1014_b N_A_917_107#_c_567_n 0.00245378f $X=-0.33 $Y=1.885
+ $X2=0.735 $Y2=2.405
cc_113 N_VPB_M1014_b N_A_917_107#_c_559_n 0.00552314f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_114 N_VPB_M1014_b N_RESET_B_c_661_n 0.0576855f $X=-0.33 $Y=1.885 $X2=0.695
+ $Y2=2.095
cc_115 N_VPB_M1014_b N_VPWR_c_694_n 0.0165123f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_694_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_117 N_VPB_c_74_p N_VPWR_c_694_n 0.0409968f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_118 N_VPB_M1014_b N_VPWR_c_697_n 0.0273337f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_697_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_120 N_VPB_c_74_p N_VPWR_c_697_n 0.0409968f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_121 N_VPB_M1014_b N_VPWR_c_700_n 0.0626284f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_700_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_123 N_VPB_c_74_p N_VPWR_c_700_n 0.0409968f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_124 N_VPB_M1014_b N_VPWR_c_703_n 0.0286727f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_703_n 0.00335473f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_126 N_VPB_c_74_p N_VPWR_c_703_n 0.0490696f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_127 N_VPB_M1014_b N_VPWR_c_706_n 0.167104f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_706_n 1.02593f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_129 N_VPB_c_74_p N_VPWR_c_706_n 0.0534074f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_130 N_VPB_M1014_b Q 0.0631548f $X=-0.33 $Y=1.885 $X2=0.695 $Y2=3.195
cc_131 VPB Q 0.00230357f $X=0 $Y=3.955 $X2=0.695 $Y2=3.195
cc_132 N_VPB_c_74_p Q 0.0389027f $X=9.36 $Y=4.07 $X2=0.695 $Y2=3.195
cc_133 N_VPB_M1014_b N_Q_c_755_n 0.0129568f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_134 N_VPB_M1014_b N_Q_c_761_n 0.0238583f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_135 N_D_M1019_g GATE 0.021795f $X=0.695 $Y=0.745 $X2=0 $Y2=0
cc_136 D N_GATE_M1007_g 0.00434665f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_137 N_D_M1019_g N_GATE_M1007_g 0.119531f $X=0.695 $Y=0.745 $X2=0 $Y2=0
cc_138 N_D_M1019_g N_A_32_107#_c_301_n 0.0261201f $X=0.695 $Y=0.745 $X2=9.36
+ $Y2=0
cc_139 D N_A_32_107#_c_303_n 0.0496842f $X=0.635 $Y=1.95 $X2=4.8 $Y2=0
cc_140 N_D_M1019_g N_A_32_107#_c_303_n 0.0407584f $X=0.695 $Y=0.745 $X2=4.8
+ $Y2=0
cc_141 D N_A_32_107#_c_304_n 0.0238298f $X=0.635 $Y=1.95 $X2=4.8 $Y2=0.057
cc_142 N_D_M1019_g N_A_32_107#_c_304_n 0.0368003f $X=0.695 $Y=0.745 $X2=4.8
+ $Y2=0.057
cc_143 N_D_M1019_g N_A_32_107#_c_308_n 3.77577e-19 $X=0.695 $Y=0.745 $X2=0 $Y2=0
cc_144 D N_VPWR_c_694_n 0.0264771f $X=0.635 $Y=1.95 $X2=9.36 $Y2=0
cc_145 N_D_M1019_g N_VPWR_c_694_n 0.0564557f $X=0.695 $Y=0.745 $X2=9.36 $Y2=0
cc_146 N_D_M1019_g N_VPWR_c_706_n 0.00864979f $X=0.695 $Y=0.745 $X2=0 $Y2=0
cc_147 N_D_M1019_g N_VGND_c_774_n 0.0402835f $X=0.695 $Y=0.745 $X2=9.36 $Y2=0
cc_148 N_D_M1019_g N_VGND_c_782_n 0.00892534f $X=0.695 $Y=0.745 $X2=0 $Y2=0
cc_149 N_GATE_M1007_g N_A_345_107#_c_200_n 0.05602f $X=1.475 $Y=0.745 $X2=9.36
+ $Y2=0
cc_150 GATE N_A_345_107#_c_191_n 0.0120469f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_151 N_GATE_M1007_g N_A_345_107#_c_191_n 0.00743135f $X=1.475 $Y=0.745 $X2=0
+ $Y2=0
cc_152 N_GATE_M1007_g N_A_345_107#_c_204_n 0.0132671f $X=1.475 $Y=0.745 $X2=4.8
+ $Y2=0
cc_153 GATE N_A_345_107#_c_193_n 0.0066556f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_GATE_M1007_g N_A_345_107#_c_193_n 0.0045768f $X=1.475 $Y=0.745 $X2=0
+ $Y2=0
cc_155 GATE N_A_345_107#_c_194_n 0.00718216f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_156 N_GATE_M1007_g N_A_345_107#_c_194_n 0.0104826f $X=1.475 $Y=0.745 $X2=0
+ $Y2=0
cc_157 GATE N_A_32_107#_c_301_n 0.0153456f $X=1.595 $Y=1.21 $X2=9.36 $Y2=0
cc_158 GATE N_A_32_107#_c_304_n 0.0696576f $X=1.595 $Y=1.21 $X2=4.8 $Y2=0.057
cc_159 N_GATE_M1007_g N_A_32_107#_c_304_n 0.0321856f $X=1.475 $Y=0.745 $X2=4.8
+ $Y2=0.057
cc_160 N_GATE_M1007_g N_A_32_107#_c_305_n 0.00130965f $X=1.475 $Y=0.745 $X2=0
+ $Y2=0
cc_161 GATE N_A_32_107#_c_308_n 0.0121081f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_162 N_GATE_M1007_g N_A_32_107#_c_308_n 0.0142419f $X=1.475 $Y=0.745 $X2=0
+ $Y2=0
cc_163 N_GATE_M1007_g N_A_462_107#_c_372_n 0.00205999f $X=1.475 $Y=0.745 $X2=0
+ $Y2=0
cc_164 N_GATE_M1007_g N_A_462_107#_c_364_n 7.12395e-19 $X=1.475 $Y=0.745
+ $X2=9.36 $Y2=0
cc_165 N_GATE_M1007_g N_A_462_107#_c_367_n 3.48386e-19 $X=1.475 $Y=0.745 $X2=0
+ $Y2=0
cc_166 N_GATE_M1007_g N_A_462_107#_c_374_n 7.193e-19 $X=1.475 $Y=0.745 $X2=4.8
+ $Y2=0
cc_167 N_GATE_M1007_g N_VPWR_c_694_n 0.0611728f $X=1.475 $Y=0.745 $X2=9.36 $Y2=0
cc_168 N_GATE_M1007_g N_VPWR_c_706_n 0.0117355f $X=1.475 $Y=0.745 $X2=0 $Y2=0
cc_169 GATE N_VGND_c_774_n 0.0675615f $X=1.595 $Y=1.21 $X2=9.36 $Y2=0
cc_170 N_GATE_M1007_g N_VGND_c_774_n 0.0357941f $X=1.475 $Y=0.745 $X2=9.36 $Y2=0
cc_171 GATE N_VGND_c_782_n 0.00861672f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_172 N_GATE_M1007_g N_VGND_c_782_n 0.00646356f $X=1.475 $Y=0.745 $X2=0 $Y2=0
cc_173 N_A_345_107#_c_192_n N_A_32_107#_M1008_g 0.0129737f $X=3.835 $Y=1.41
+ $X2=0 $Y2=0
cc_174 N_A_345_107#_c_196_n N_A_32_107#_M1008_g 0.00223582f $X=4.27 $Y=1.77
+ $X2=0 $Y2=0
cc_175 N_A_345_107#_M1018_g N_A_32_107#_M1008_g 0.0359267f $X=2.845 $Y=0.745
+ $X2=0 $Y2=0
cc_176 N_A_345_107#_c_203_n N_A_32_107#_M1010_g 0.0241186f $X=3.835 $Y=2.11
+ $X2=0 $Y2=0
cc_177 N_A_345_107#_c_196_n N_A_32_107#_M1010_g 0.00524175f $X=4.27 $Y=1.77
+ $X2=0 $Y2=0
cc_178 N_A_345_107#_c_197_n N_A_32_107#_M1010_g 0.0608605f $X=4.27 $Y=1.77 $X2=0
+ $Y2=0
cc_179 N_A_345_107#_M1018_g N_A_32_107#_M1010_g 0.0523716f $X=2.845 $Y=0.745
+ $X2=0 $Y2=0
cc_180 N_A_345_107#_c_203_n N_A_32_107#_c_305_n 0.111314f $X=3.835 $Y=2.11 $X2=0
+ $Y2=0
cc_181 N_A_345_107#_c_204_n N_A_32_107#_c_305_n 0.0190597f $X=2.03 $Y=2.11 $X2=0
+ $Y2=0
cc_182 N_A_345_107#_c_192_n N_A_32_107#_c_305_n 0.102732f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_183 N_A_345_107#_c_193_n N_A_32_107#_c_305_n 0.0134479f $X=2.145 $Y=1.41
+ $X2=0 $Y2=0
cc_184 N_A_345_107#_c_196_n N_A_32_107#_c_305_n 0.0134486f $X=4.27 $Y=1.77 $X2=0
+ $Y2=0
cc_185 N_A_345_107#_M1018_g N_A_32_107#_c_305_n 0.0277217f $X=2.845 $Y=0.745
+ $X2=0 $Y2=0
cc_186 N_A_345_107#_c_188_n N_A_32_107#_c_306_n 0.0608605f $X=4.585 $Y=1.68
+ $X2=0 $Y2=0
cc_187 N_A_345_107#_c_203_n N_A_32_107#_c_306_n 0.0019113f $X=3.835 $Y=2.11
+ $X2=0 $Y2=0
cc_188 N_A_345_107#_c_192_n N_A_32_107#_c_306_n 0.0134327f $X=3.835 $Y=1.41
+ $X2=0 $Y2=0
cc_189 N_A_345_107#_c_196_n N_A_32_107#_c_306_n 0.0210704f $X=4.27 $Y=1.77 $X2=0
+ $Y2=0
cc_190 N_A_345_107#_M1018_g N_A_32_107#_c_306_n 0.0367665f $X=2.845 $Y=0.745
+ $X2=0 $Y2=0
cc_191 N_A_345_107#_c_204_n N_A_32_107#_c_308_n 0.00768214f $X=2.03 $Y=2.11
+ $X2=0 $Y2=0
cc_192 N_A_345_107#_c_200_n N_A_462_107#_c_372_n 0.0433374f $X=1.865 $Y=2.945
+ $X2=0 $Y2=0
cc_193 N_A_345_107#_M1018_g N_A_462_107#_c_372_n 0.0204855f $X=2.845 $Y=0.745
+ $X2=0 $Y2=0
cc_194 N_A_345_107#_c_194_n N_A_462_107#_c_364_n 0.03055f $X=2.06 $Y=0.745
+ $X2=9.36 $Y2=0
cc_195 N_A_345_107#_M1018_g N_A_462_107#_c_364_n 0.0141412f $X=2.845 $Y=0.745
+ $X2=9.36 $Y2=0
cc_196 N_A_345_107#_c_192_n N_A_462_107#_c_366_n 0.0807219f $X=3.835 $Y=1.41
+ $X2=0 $Y2=0
cc_197 N_A_345_107#_c_196_n N_A_462_107#_c_366_n 0.0201316f $X=4.27 $Y=1.77
+ $X2=0 $Y2=0
cc_198 N_A_345_107#_M1018_g N_A_462_107#_c_366_n 0.0235038f $X=2.845 $Y=0.745
+ $X2=0 $Y2=0
cc_199 N_A_345_107#_c_191_n N_A_462_107#_c_367_n 0.0104032f $X=2.06 $Y=1.325
+ $X2=0 $Y2=0
cc_200 N_A_345_107#_c_192_n N_A_462_107#_c_367_n 0.0199928f $X=3.835 $Y=1.41
+ $X2=0 $Y2=0
cc_201 N_A_345_107#_c_194_n N_A_462_107#_c_367_n 0.00141515f $X=2.06 $Y=0.745
+ $X2=0 $Y2=0
cc_202 N_A_345_107#_M1018_g N_A_462_107#_c_367_n 0.00394456f $X=2.845 $Y=0.745
+ $X2=0 $Y2=0
cc_203 N_A_345_107#_c_187_n N_A_462_107#_c_373_n 6.22937e-19 $X=4.98 $Y=1.68
+ $X2=0 $Y2=0
cc_204 N_A_345_107#_c_203_n N_A_462_107#_c_373_n 0.0807223f $X=3.835 $Y=2.11
+ $X2=0 $Y2=0
cc_205 N_A_345_107#_c_196_n N_A_462_107#_c_373_n 0.0450251f $X=4.27 $Y=1.77
+ $X2=0 $Y2=0
cc_206 N_A_345_107#_c_197_n N_A_462_107#_c_373_n 0.0441983f $X=4.27 $Y=1.77
+ $X2=0 $Y2=0
cc_207 N_A_345_107#_M1018_g N_A_462_107#_c_373_n 0.0282719f $X=2.845 $Y=0.745
+ $X2=0 $Y2=0
cc_208 N_A_345_107#_c_200_n N_A_462_107#_c_374_n 0.011172f $X=1.865 $Y=2.945
+ $X2=4.8 $Y2=0
cc_209 N_A_345_107#_c_203_n N_A_462_107#_c_374_n 0.0265557f $X=3.835 $Y=2.11
+ $X2=4.8 $Y2=0
cc_210 N_A_345_107#_M1018_g N_A_462_107#_c_374_n 0.0023611f $X=2.845 $Y=0.745
+ $X2=4.8 $Y2=0
cc_211 N_A_345_107#_c_187_n N_A_462_107#_c_368_n 0.0160832f $X=4.98 $Y=1.68
+ $X2=4.8 $Y2=0.057
cc_212 N_A_345_107#_M1004_g N_A_462_107#_c_368_n 0.00577781f $X=5.23 $Y=0.745
+ $X2=4.8 $Y2=0.057
cc_213 N_A_345_107#_c_196_n N_A_462_107#_c_368_n 0.0336636f $X=4.27 $Y=1.77
+ $X2=4.8 $Y2=0.057
cc_214 N_A_345_107#_c_197_n N_A_462_107#_c_368_n 0.00605806f $X=4.27 $Y=1.77
+ $X2=4.8 $Y2=0.057
cc_215 N_A_345_107#_c_187_n N_A_462_107#_c_369_n 9.7e-19 $X=4.98 $Y=1.68 $X2=4.8
+ $Y2=0.058
cc_216 N_A_345_107#_c_188_n N_A_462_107#_c_369_n 0.00147349f $X=4.585 $Y=1.68
+ $X2=4.8 $Y2=0.058
cc_217 N_A_345_107#_M1004_g N_A_462_107#_c_369_n 0.00143594f $X=5.23 $Y=0.745
+ $X2=4.8 $Y2=0.058
cc_218 N_A_345_107#_c_196_n N_A_462_107#_c_369_n 0.022938f $X=4.27 $Y=1.77
+ $X2=4.8 $Y2=0.058
cc_219 N_A_345_107#_c_187_n N_A_462_107#_c_376_n 0.00339612f $X=4.98 $Y=1.68
+ $X2=0 $Y2=0
cc_220 N_A_345_107#_c_196_n N_A_462_107#_c_376_n 0.019324f $X=4.27 $Y=1.77 $X2=0
+ $Y2=0
cc_221 N_A_345_107#_c_197_n N_A_462_107#_c_376_n 0.0073857f $X=4.27 $Y=1.77
+ $X2=0 $Y2=0
cc_222 N_A_345_107#_c_187_n N_A_462_107#_c_377_n 0.0450016f $X=4.98 $Y=1.68
+ $X2=0 $Y2=0
cc_223 N_A_345_107#_c_197_n N_A_462_107#_c_377_n 0.0203584f $X=4.27 $Y=1.77
+ $X2=0 $Y2=0
cc_224 N_A_345_107#_c_188_n N_A_462_107#_M1012_g 0.0330968f $X=4.585 $Y=1.68
+ $X2=0 $Y2=0
cc_225 N_A_345_107#_M1004_g N_A_462_107#_M1012_g 0.023235f $X=5.23 $Y=0.745
+ $X2=0 $Y2=0
cc_226 N_A_345_107#_c_196_n N_A_462_107#_M1012_g 0.00133047f $X=4.27 $Y=1.77
+ $X2=0 $Y2=0
cc_227 N_A_345_107#_c_197_n N_A_462_107#_c_378_n 0.0176742f $X=4.27 $Y=1.77
+ $X2=0 $Y2=0
cc_228 N_A_345_107#_M1004_g N_A_1138_81#_c_479_n 2.24396e-19 $X=5.23 $Y=0.745
+ $X2=9.36 $Y2=0
cc_229 N_A_345_107#_M1004_g N_A_1138_81#_M1009_g 0.0899136f $X=5.23 $Y=0.745
+ $X2=0 $Y2=0
cc_230 N_A_345_107#_c_197_n N_A_917_107#_c_566_n 0.0109662f $X=4.27 $Y=1.77
+ $X2=0 $Y2=0
cc_231 N_A_345_107#_c_197_n N_A_917_107#_c_570_n 0.00519821f $X=4.27 $Y=1.77
+ $X2=0 $Y2=0
cc_232 N_A_345_107#_M1004_g N_A_917_107#_c_557_n 0.00776886f $X=5.23 $Y=0.745
+ $X2=0 $Y2=0
cc_233 N_A_345_107#_M1004_g N_A_917_107#_c_572_n 0.0128119f $X=5.23 $Y=0.745
+ $X2=4.8 $Y2=0
cc_234 N_A_345_107#_c_187_n N_A_917_107#_c_558_n 3.17269e-19 $X=4.98 $Y=1.68
+ $X2=0 $Y2=0
cc_235 N_A_345_107#_M1004_g N_A_917_107#_c_558_n 0.00688368f $X=5.23 $Y=0.745
+ $X2=0 $Y2=0
cc_236 N_A_345_107#_c_187_n N_A_917_107#_c_559_n 0.00726848f $X=4.98 $Y=1.68
+ $X2=4.8 $Y2=0.058
cc_237 N_A_345_107#_M1004_g N_A_917_107#_c_559_n 0.00953789f $X=5.23 $Y=0.745
+ $X2=4.8 $Y2=0.058
cc_238 N_A_345_107#_c_187_n N_A_917_107#_c_561_n 0.00488184f $X=4.98 $Y=1.68
+ $X2=0 $Y2=0
cc_239 N_A_345_107#_M1004_g N_A_917_107#_c_561_n 0.0186293f $X=5.23 $Y=0.745
+ $X2=0 $Y2=0
cc_240 N_A_345_107#_M1004_g N_A_917_107#_c_563_n 0.00694558f $X=5.23 $Y=0.745
+ $X2=0 $Y2=0
cc_241 N_A_345_107#_c_200_n N_VPWR_c_694_n 0.0605993f $X=1.865 $Y=2.945 $X2=9.36
+ $Y2=0
cc_242 N_A_345_107#_c_197_n N_VPWR_c_697_n 0.00338454f $X=4.27 $Y=1.77 $X2=4.8
+ $Y2=0.058
cc_243 N_A_345_107#_M1018_g N_VPWR_c_697_n 0.0419815f $X=2.845 $Y=0.745 $X2=4.8
+ $Y2=0.058
cc_244 N_A_345_107#_c_200_n N_VPWR_c_706_n 0.0367193f $X=1.865 $Y=2.945 $X2=0
+ $Y2=0
cc_245 N_A_345_107#_c_197_n N_VPWR_c_706_n 0.016332f $X=4.27 $Y=1.77 $X2=0 $Y2=0
cc_246 N_A_345_107#_M1018_g N_VPWR_c_706_n 0.00672879f $X=2.845 $Y=0.745 $X2=0
+ $Y2=0
cc_247 N_A_345_107#_c_194_n N_VGND_c_774_n 0.036741f $X=2.06 $Y=0.745 $X2=9.36
+ $Y2=0
cc_248 N_A_345_107#_M1018_g N_VGND_c_776_n 0.0263602f $X=2.845 $Y=0.745 $X2=4.8
+ $Y2=0.058
cc_249 N_A_345_107#_M1004_g N_VGND_c_778_n 0.00782651f $X=5.23 $Y=0.745 $X2=0
+ $Y2=0
cc_250 N_A_345_107#_M1004_g N_VGND_c_782_n 0.0145098f $X=5.23 $Y=0.745 $X2=0
+ $Y2=0
cc_251 N_A_345_107#_c_191_n N_VGND_c_782_n 4.53342e-19 $X=2.06 $Y=1.325 $X2=0
+ $Y2=0
cc_252 N_A_345_107#_c_194_n N_VGND_c_782_n 0.0300567f $X=2.06 $Y=0.745 $X2=0
+ $Y2=0
cc_253 N_A_345_107#_M1018_g N_VGND_c_782_n 0.00586905f $X=2.845 $Y=0.745 $X2=0
+ $Y2=0
cc_254 N_A_32_107#_M1008_g N_A_462_107#_c_366_n 0.0259423f $X=3.625 $Y=0.745
+ $X2=0 $Y2=0
cc_255 N_A_32_107#_c_306_n N_A_462_107#_c_366_n 3.61041e-19 $X=3.49 $Y=1.76
+ $X2=0 $Y2=0
cc_256 N_A_32_107#_M1010_g N_A_462_107#_c_373_n 0.0293175f $X=3.625 $Y=2.83
+ $X2=0 $Y2=0
cc_257 N_A_32_107#_M1008_g N_A_462_107#_c_369_n 0.00111867f $X=3.625 $Y=0.745
+ $X2=4.8 $Y2=0.058
cc_258 N_A_32_107#_M1008_g N_A_462_107#_M1012_g 0.0712966f $X=3.625 $Y=0.745
+ $X2=0 $Y2=0
cc_259 N_A_32_107#_M1010_g N_A_917_107#_c_566_n 0.00106623f $X=3.625 $Y=2.83
+ $X2=0 $Y2=0
cc_260 N_A_32_107#_M1010_g N_A_917_107#_c_570_n 5.139e-19 $X=3.625 $Y=2.83 $X2=0
+ $Y2=0
cc_261 N_A_32_107#_c_303_n N_VPWR_c_694_n 0.0366474f $X=0.305 $Y=2.945 $X2=9.36
+ $Y2=0
cc_262 N_A_32_107#_M1010_g N_VPWR_c_697_n 0.0475895f $X=3.625 $Y=2.83 $X2=4.8
+ $Y2=0.058
cc_263 N_A_32_107#_M1014_s N_VPWR_c_706_n 0.00221032f $X=0.16 $Y=2.82 $X2=0
+ $Y2=0
cc_264 N_A_32_107#_M1010_g N_VPWR_c_706_n 0.00411567f $X=3.625 $Y=2.83 $X2=0
+ $Y2=0
cc_265 N_A_32_107#_c_303_n N_VPWR_c_706_n 0.028278f $X=0.305 $Y=2.945 $X2=0
+ $Y2=0
cc_266 N_A_32_107#_c_301_n N_VGND_c_774_n 0.0231654f $X=0.305 $Y=0.745 $X2=9.36
+ $Y2=0
cc_267 N_A_32_107#_c_304_n N_VGND_c_774_n 9.25196e-19 $X=1.625 $Y=1.665 $X2=9.36
+ $Y2=0
cc_268 N_A_32_107#_M1008_g N_VGND_c_776_n 0.0332758f $X=3.625 $Y=0.745 $X2=4.8
+ $Y2=0.058
cc_269 N_A_32_107#_M1019_s N_VGND_c_782_n 0.00221032f $X=0.16 $Y=0.535 $X2=0
+ $Y2=0
cc_270 N_A_32_107#_M1008_g N_VGND_c_782_n 0.0042168f $X=3.625 $Y=0.745 $X2=0
+ $Y2=0
cc_271 N_A_32_107#_c_301_n N_VGND_c_782_n 0.0264336f $X=0.305 $Y=0.745 $X2=0
+ $Y2=0
cc_272 N_A_462_107#_c_377_n N_A_1138_81#_M1009_g 0.0679742f $X=5.01 $Y=2.13
+ $X2=0 $Y2=0
cc_273 N_A_462_107#_c_376_n N_A_917_107#_M1016_d 0.00302109f $X=5.01 $Y=2.13
+ $X2=0 $Y2=0
cc_274 N_A_462_107#_c_378_n N_A_917_107#_c_566_n 0.00316525f $X=5.152 $Y=2.345
+ $X2=0 $Y2=0
cc_275 N_A_462_107#_c_376_n N_A_917_107#_c_567_n 0.00878025f $X=5.01 $Y=2.13
+ $X2=9.36 $Y2=0
cc_276 N_A_462_107#_c_377_n N_A_917_107#_c_567_n 0.00161343f $X=5.01 $Y=2.13
+ $X2=9.36 $Y2=0
cc_277 N_A_462_107#_c_378_n N_A_917_107#_c_567_n 0.0336359f $X=5.152 $Y=2.345
+ $X2=9.36 $Y2=0
cc_278 N_A_462_107#_c_373_n N_A_917_107#_c_570_n 0.00177995f $X=4.615 $Y=2.46
+ $X2=0 $Y2=0
cc_279 N_A_462_107#_c_376_n N_A_917_107#_c_570_n 0.0164313f $X=5.01 $Y=2.13
+ $X2=0 $Y2=0
cc_280 N_A_462_107#_c_377_n N_A_917_107#_c_570_n 0.00137418f $X=5.01 $Y=2.13
+ $X2=0 $Y2=0
cc_281 N_A_462_107#_c_369_n N_A_917_107#_c_557_n 0.00658319f $X=4.34 $Y=1.23
+ $X2=0 $Y2=0
cc_282 N_A_462_107#_M1012_g N_A_917_107#_c_557_n 0.00138521f $X=4.335 $Y=0.745
+ $X2=0 $Y2=0
cc_283 N_A_462_107#_c_376_n N_A_917_107#_c_572_n 9.64928e-19 $X=5.01 $Y=2.13
+ $X2=4.8 $Y2=0
cc_284 N_A_462_107#_c_377_n N_A_917_107#_c_572_n 6.65012e-19 $X=5.01 $Y=2.13
+ $X2=4.8 $Y2=0
cc_285 N_A_462_107#_c_369_n N_A_917_107#_c_558_n 0.0126598f $X=4.34 $Y=1.23
+ $X2=0 $Y2=0
cc_286 N_A_462_107#_c_376_n N_A_917_107#_c_558_n 0.00445268f $X=5.01 $Y=2.13
+ $X2=0 $Y2=0
cc_287 N_A_462_107#_M1012_g N_A_917_107#_c_558_n 7.93318e-19 $X=4.335 $Y=0.745
+ $X2=0 $Y2=0
cc_288 N_A_462_107#_c_368_n N_A_917_107#_c_559_n 0.0165479f $X=4.7 $Y=1.965
+ $X2=4.8 $Y2=0.058
cc_289 N_A_462_107#_c_369_n N_A_917_107#_c_559_n 0.00159024f $X=4.34 $Y=1.23
+ $X2=4.8 $Y2=0.058
cc_290 N_A_462_107#_c_376_n N_A_917_107#_c_559_n 0.031246f $X=5.01 $Y=2.13
+ $X2=4.8 $Y2=0.058
cc_291 N_A_462_107#_c_377_n N_A_917_107#_c_559_n 0.0124257f $X=5.01 $Y=2.13
+ $X2=4.8 $Y2=0.058
cc_292 N_A_462_107#_c_378_n N_A_917_107#_c_559_n 0.0172078f $X=5.152 $Y=2.345
+ $X2=4.8 $Y2=0.058
cc_293 N_A_462_107#_c_369_n N_A_917_107#_c_561_n 0.0092442f $X=4.34 $Y=1.23
+ $X2=0 $Y2=0
cc_294 N_A_462_107#_M1012_g N_A_917_107#_c_561_n 0.013933f $X=4.335 $Y=0.745
+ $X2=0 $Y2=0
cc_295 N_A_462_107#_c_373_n N_VPWR_M1001_d 0.00180746f $X=4.615 $Y=2.46 $X2=0
+ $Y2=0
cc_296 N_A_462_107#_c_372_n N_VPWR_c_697_n 0.0394618f $X=2.455 $Y=2.58 $X2=4.8
+ $Y2=0.058
cc_297 N_A_462_107#_c_373_n N_VPWR_c_697_n 0.0615323f $X=4.615 $Y=2.46 $X2=4.8
+ $Y2=0.058
cc_298 N_A_462_107#_c_377_n N_VPWR_c_700_n 7.05769e-19 $X=5.01 $Y=2.13 $X2=0
+ $Y2=0
cc_299 N_A_462_107#_c_378_n N_VPWR_c_700_n 7.77477e-19 $X=5.152 $Y=2.345 $X2=0
+ $Y2=0
cc_300 N_A_462_107#_c_372_n N_VPWR_c_706_n 0.0181496f $X=2.455 $Y=2.58 $X2=0
+ $Y2=0
cc_301 N_A_462_107#_c_378_n N_VPWR_c_706_n 0.0134517f $X=5.152 $Y=2.345 $X2=0
+ $Y2=0
cc_302 N_A_462_107#_c_373_n A_775_491# 0.00366293f $X=4.615 $Y=2.46 $X2=0 $Y2=0
cc_303 N_A_462_107#_c_364_n N_VGND_c_776_n 0.0206222f $X=2.455 $Y=0.745 $X2=4.8
+ $Y2=0.058
cc_304 N_A_462_107#_c_366_n N_VGND_c_776_n 0.0593584f $X=4.185 $Y=1.06 $X2=4.8
+ $Y2=0.058
cc_305 N_A_462_107#_M1012_g N_VGND_c_776_n 0.00296386f $X=4.335 $Y=0.745 $X2=4.8
+ $Y2=0.058
cc_306 N_A_462_107#_M1018_s N_VGND_c_782_n 0.00254395f $X=2.31 $Y=0.535 $X2=0
+ $Y2=0
cc_307 N_A_462_107#_c_364_n N_VGND_c_782_n 0.0234066f $X=2.455 $Y=0.745 $X2=0
+ $Y2=0
cc_308 N_A_462_107#_c_366_n N_VGND_c_782_n 0.0272816f $X=4.185 $Y=1.06 $X2=0
+ $Y2=0
cc_309 N_A_462_107#_c_369_n N_VGND_c_782_n 0.017927f $X=4.34 $Y=1.23 $X2=0 $Y2=0
cc_310 N_A_462_107#_M1012_g N_VGND_c_782_n 0.0194876f $X=4.335 $Y=0.745 $X2=0
+ $Y2=0
cc_311 N_A_1138_81#_c_479_n N_A_917_107#_M1011_g 6.06951e-19 $X=5.975 $Y=1.63
+ $X2=0 $Y2=0
cc_312 N_A_1138_81#_c_473_n N_A_917_107#_M1011_g 0.033663f $X=6.96 $Y=1.99 $X2=0
+ $Y2=0
cc_313 N_A_1138_81#_c_465_n N_A_917_107#_M1011_g 0.00556646f $X=7.045 $Y=1.905
+ $X2=0 $Y2=0
cc_314 N_A_1138_81#_c_474_n N_A_917_107#_M1011_g 0.0123286f $X=7.175 $Y=2.205
+ $X2=0 $Y2=0
cc_315 N_A_1138_81#_c_475_n N_A_917_107#_M1011_g 0.0306275f $X=7.225 $Y=2.34
+ $X2=0 $Y2=0
cc_316 N_A_1138_81#_M1009_g N_A_917_107#_M1011_g 0.0286275f $X=5.94 $Y=0.745
+ $X2=0 $Y2=0
cc_317 N_A_1138_81#_c_465_n N_A_917_107#_c_555_n 0.00293358f $X=7.045 $Y=1.905
+ $X2=0.24 $Y2=0
cc_318 N_A_1138_81#_c_466_n N_A_917_107#_c_555_n 0.0167752f $X=6.92 $Y=0.745
+ $X2=0.24 $Y2=0
cc_319 N_A_1138_81#_M1009_g N_A_917_107#_c_567_n 6.44081e-19 $X=5.94 $Y=0.745
+ $X2=9.36 $Y2=0
cc_320 N_A_1138_81#_M1009_g N_A_917_107#_c_557_n 6.80723e-19 $X=5.94 $Y=0.745
+ $X2=0 $Y2=0
cc_321 N_A_1138_81#_c_479_n N_A_917_107#_c_559_n 0.0193884f $X=5.975 $Y=1.63
+ $X2=4.8 $Y2=0.058
cc_322 N_A_1138_81#_c_493_p N_A_917_107#_c_559_n 0.00920426f $X=6.14 $Y=1.99
+ $X2=4.8 $Y2=0.058
cc_323 N_A_1138_81#_M1009_g N_A_917_107#_c_559_n 0.0173632f $X=5.94 $Y=0.745
+ $X2=4.8 $Y2=0.058
cc_324 N_A_1138_81#_c_479_n N_A_917_107#_c_560_n 0.0234404f $X=5.975 $Y=1.63
+ $X2=4.8 $Y2=0.058
cc_325 N_A_1138_81#_c_473_n N_A_917_107#_c_560_n 0.0097304f $X=6.96 $Y=1.99
+ $X2=4.8 $Y2=0.058
cc_326 N_A_1138_81#_M1009_g N_A_917_107#_c_560_n 0.0294832f $X=5.94 $Y=0.745
+ $X2=4.8 $Y2=0.058
cc_327 N_A_1138_81#_M1009_g N_A_917_107#_c_561_n 4.085e-19 $X=5.94 $Y=0.745
+ $X2=0 $Y2=0
cc_328 N_A_1138_81#_c_479_n N_A_917_107#_c_621_n 0.00928073f $X=5.975 $Y=1.63
+ $X2=0 $Y2=0
cc_329 N_A_1138_81#_c_473_n N_A_917_107#_c_621_n 0.0239448f $X=6.96 $Y=1.99
+ $X2=0 $Y2=0
cc_330 N_A_1138_81#_c_465_n N_A_917_107#_c_621_n 0.0382514f $X=7.045 $Y=1.905
+ $X2=0 $Y2=0
cc_331 N_A_1138_81#_c_466_n N_A_917_107#_c_621_n 0.00190709f $X=6.92 $Y=0.745
+ $X2=0 $Y2=0
cc_332 N_A_1138_81#_M1009_g N_A_917_107#_c_621_n 0.00204273f $X=5.94 $Y=0.745
+ $X2=0 $Y2=0
cc_333 N_A_1138_81#_c_479_n N_A_917_107#_c_564_n 0.00132035f $X=5.975 $Y=1.63
+ $X2=0 $Y2=0
cc_334 N_A_1138_81#_c_473_n N_A_917_107#_c_564_n 0.00455724f $X=6.96 $Y=1.99
+ $X2=0 $Y2=0
cc_335 N_A_1138_81#_c_465_n N_A_917_107#_c_564_n 0.0398329f $X=7.045 $Y=1.905
+ $X2=0 $Y2=0
cc_336 N_A_1138_81#_c_474_n N_A_917_107#_c_564_n 0.00707848f $X=7.175 $Y=2.205
+ $X2=0 $Y2=0
cc_337 N_A_1138_81#_c_476_n N_A_917_107#_c_564_n 4.44732e-19 $X=8.3 $Y=2.12
+ $X2=0 $Y2=0
cc_338 N_A_1138_81#_c_466_n N_A_917_107#_c_564_n 0.0100584f $X=6.92 $Y=0.745
+ $X2=0 $Y2=0
cc_339 N_A_1138_81#_M1009_g N_A_917_107#_c_564_n 0.0455403f $X=5.94 $Y=0.745
+ $X2=0 $Y2=0
cc_340 N_A_1138_81#_M1015_g RESET_B 0.00306412f $X=8.915 $Y=0.91 $X2=0 $Y2=0
cc_341 N_A_1138_81#_c_466_n RESET_B 0.027012f $X=6.92 $Y=0.745 $X2=0 $Y2=0
cc_342 N_A_1138_81#_M1015_g RESET_B 0.00389247f $X=8.915 $Y=0.91 $X2=0 $Y2=0
cc_343 N_A_1138_81#_c_465_n RESET_B 0.0165737f $X=7.045 $Y=1.905 $X2=0 $Y2=0
cc_344 N_A_1138_81#_c_476_n RESET_B 0.0413217f $X=8.3 $Y=2.12 $X2=0 $Y2=0
cc_345 N_A_1138_81#_c_516_p RESET_B 0.0117873f $X=8.465 $Y=1.83 $X2=0 $Y2=0
cc_346 N_A_1138_81#_c_469_n RESET_B 0.00337612f $X=8.915 $Y=1.855 $X2=0 $Y2=0
cc_347 N_A_1138_81#_c_465_n N_RESET_B_c_661_n 0.00295972f $X=7.045 $Y=1.905
+ $X2=0 $Y2=0
cc_348 N_A_1138_81#_c_474_n N_RESET_B_c_661_n 0.00643371f $X=7.175 $Y=2.205
+ $X2=0 $Y2=0
cc_349 N_A_1138_81#_c_475_n N_RESET_B_c_661_n 0.0214736f $X=7.225 $Y=2.34 $X2=0
+ $Y2=0
cc_350 N_A_1138_81#_c_476_n N_RESET_B_c_661_n 0.0295313f $X=8.3 $Y=2.12 $X2=0
+ $Y2=0
cc_351 N_A_1138_81#_c_516_p N_RESET_B_c_661_n 0.00154627f $X=8.465 $Y=1.83 $X2=0
+ $Y2=0
cc_352 N_A_1138_81#_c_469_n N_RESET_B_c_661_n 0.0348242f $X=8.915 $Y=1.855 $X2=0
+ $Y2=0
cc_353 N_A_1138_81#_M1015_g N_RESET_B_M1003_g 0.0193317f $X=8.915 $Y=0.91 $X2=0
+ $Y2=0
cc_354 N_A_1138_81#_c_476_n N_RESET_B_M1003_g 0.00446081f $X=8.3 $Y=2.12 $X2=0
+ $Y2=0
cc_355 N_A_1138_81#_c_466_n N_RESET_B_M1003_g 0.00155691f $X=6.92 $Y=0.745 $X2=0
+ $Y2=0
cc_356 N_A_1138_81#_c_469_n N_RESET_B_M1003_g 8.09768e-19 $X=8.915 $Y=1.855
+ $X2=0 $Y2=0
cc_357 N_A_1138_81#_c_473_n N_VPWR_c_700_n 0.0376571f $X=6.96 $Y=1.99 $X2=0
+ $Y2=0
cc_358 N_A_1138_81#_c_493_p N_VPWR_c_700_n 0.0262475f $X=6.14 $Y=1.99 $X2=0
+ $Y2=0
cc_359 N_A_1138_81#_c_475_n N_VPWR_c_700_n 0.038062f $X=7.225 $Y=2.34 $X2=0
+ $Y2=0
cc_360 N_A_1138_81#_M1009_g N_VPWR_c_700_n 0.0731046f $X=5.94 $Y=0.745 $X2=0
+ $Y2=0
cc_361 N_A_1138_81#_c_470_n N_VPWR_c_703_n 0.060007f $X=8.51 $Y=2.105 $X2=0
+ $Y2=0
cc_362 N_A_1138_81#_c_475_n N_VPWR_c_703_n 0.047969f $X=7.225 $Y=2.34 $X2=0
+ $Y2=0
cc_363 N_A_1138_81#_c_476_n N_VPWR_c_703_n 0.0506481f $X=8.3 $Y=2.12 $X2=0 $Y2=0
cc_364 N_A_1138_81#_c_516_p N_VPWR_c_703_n 0.0155063f $X=8.465 $Y=1.83 $X2=0
+ $Y2=0
cc_365 N_A_1138_81#_c_470_n N_VPWR_c_706_n 0.013214f $X=8.51 $Y=2.105 $X2=0
+ $Y2=0
cc_366 N_A_1138_81#_c_475_n N_VPWR_c_706_n 0.0183081f $X=7.225 $Y=2.34 $X2=0
+ $Y2=0
cc_367 N_A_1138_81#_M1009_g N_VPWR_c_706_n 4.30453e-19 $X=5.94 $Y=0.745 $X2=0
+ $Y2=0
cc_368 N_A_1138_81#_c_470_n Q 0.0230529f $X=8.51 $Y=2.105 $X2=0 $Y2=0
cc_369 N_A_1138_81#_c_470_n N_Q_c_755_n 0.0016249f $X=8.51 $Y=2.105 $X2=4.8
+ $Y2=0.057
cc_370 N_A_1138_81#_M1015_g N_Q_c_755_n 0.0381621f $X=8.915 $Y=0.91 $X2=4.8
+ $Y2=0.057
cc_371 N_A_1138_81#_c_516_p N_Q_c_755_n 0.014835f $X=8.465 $Y=1.83 $X2=4.8
+ $Y2=0.057
cc_372 N_A_1138_81#_c_469_n N_Q_c_755_n 0.0265245f $X=8.915 $Y=1.855 $X2=4.8
+ $Y2=0.057
cc_373 N_A_1138_81#_c_470_n N_Q_c_761_n 0.0151395f $X=8.51 $Y=2.105 $X2=0 $Y2=0
cc_374 N_A_1138_81#_c_516_p N_Q_c_761_n 0.00176972f $X=8.465 $Y=1.83 $X2=0 $Y2=0
cc_375 N_A_1138_81#_c_469_n N_Q_c_761_n 0.020503f $X=8.915 $Y=1.855 $X2=0 $Y2=0
cc_376 N_A_1138_81#_c_466_n N_VGND_c_778_n 0.0307575f $X=6.92 $Y=0.745 $X2=0
+ $Y2=0
cc_377 N_A_1138_81#_M1009_g N_VGND_c_778_n 0.0498108f $X=5.94 $Y=0.745 $X2=0
+ $Y2=0
cc_378 N_A_1138_81#_M1015_g N_VGND_c_780_n 0.0538744f $X=8.915 $Y=0.91 $X2=0
+ $Y2=0
cc_379 N_A_1138_81#_c_516_p N_VGND_c_780_n 0.0168968f $X=8.465 $Y=1.83 $X2=0
+ $Y2=0
cc_380 N_A_1138_81#_c_469_n N_VGND_c_780_n 0.0100995f $X=8.915 $Y=1.855 $X2=0
+ $Y2=0
cc_381 N_A_1138_81#_M1015_g N_VGND_c_782_n 0.0159812f $X=8.915 $Y=0.91 $X2=0
+ $Y2=0
cc_382 N_A_1138_81#_c_466_n N_VGND_c_782_n 0.0287222f $X=6.92 $Y=0.745 $X2=0
+ $Y2=0
cc_383 N_A_917_107#_c_555_n RESET_B 0.00988692f $X=7.31 $Y=1.065 $X2=0 $Y2=0
cc_384 N_A_917_107#_c_564_n RESET_B 0.0128071f $X=6.835 $Y=1.435 $X2=0 $Y2=0
cc_385 N_A_917_107#_c_564_n RESET_B 0.00104689f $X=6.835 $Y=1.435 $X2=0 $Y2=0
cc_386 N_A_917_107#_c_564_n N_RESET_B_c_661_n 0.0545483f $X=6.835 $Y=1.435 $X2=0
+ $Y2=0
cc_387 N_A_917_107#_c_555_n N_RESET_B_M1003_g 0.0681078f $X=7.31 $Y=1.065 $X2=0
+ $Y2=0
cc_388 N_A_917_107#_M1011_g N_VPWR_c_700_n 0.0319005f $X=6.835 $Y=2.59 $X2=0
+ $Y2=0
cc_389 N_A_917_107#_c_567_n N_VPWR_c_700_n 0.00768914f $X=5.355 $Y=2.81 $X2=0
+ $Y2=0
cc_390 N_A_917_107#_c_559_n N_VPWR_c_700_n 0.0260149f $X=5.44 $Y=2.725 $X2=0
+ $Y2=0
cc_391 N_A_917_107#_M1011_g N_VPWR_c_703_n 6.30651e-19 $X=6.835 $Y=2.59 $X2=0
+ $Y2=0
cc_392 N_A_917_107#_M1011_g N_VPWR_c_706_n 0.0122219f $X=6.835 $Y=2.59 $X2=0
+ $Y2=0
cc_393 N_A_917_107#_c_566_n N_VPWR_c_706_n 0.0176598f $X=4.725 $Y=2.895 $X2=0
+ $Y2=0
cc_394 N_A_917_107#_c_567_n N_VPWR_c_706_n 0.0211801f $X=5.355 $Y=2.81 $X2=0
+ $Y2=0
cc_395 N_A_917_107#_c_555_n N_VGND_c_778_n 0.00261609f $X=7.31 $Y=1.065 $X2=0
+ $Y2=0
cc_396 N_A_917_107#_c_560_n N_VGND_c_778_n 0.0662492f $X=6.45 $Y=1.26 $X2=0
+ $Y2=0
cc_397 N_A_917_107#_c_561_n N_VGND_c_778_n 0.0191233f $X=5.05 $Y=0.745 $X2=0
+ $Y2=0
cc_398 N_A_917_107#_c_621_n N_VGND_c_778_n 0.00362506f $X=6.615 $Y=1.28 $X2=0
+ $Y2=0
cc_399 N_A_917_107#_c_564_n N_VGND_c_778_n 0.00199981f $X=6.835 $Y=1.435 $X2=0
+ $Y2=0
cc_400 N_A_917_107#_M1012_d N_VGND_c_782_n 0.00129126f $X=4.585 $Y=0.535 $X2=0
+ $Y2=0
cc_401 N_A_917_107#_c_555_n N_VGND_c_782_n 0.0289761f $X=7.31 $Y=1.065 $X2=0
+ $Y2=0
cc_402 N_A_917_107#_c_557_n N_VGND_c_782_n 4.52779e-19 $X=5.05 $Y=1.175 $X2=0
+ $Y2=0
cc_403 N_A_917_107#_c_572_n N_VGND_c_782_n 0.00608199f $X=5.355 $Y=1.26 $X2=0
+ $Y2=0
cc_404 N_A_917_107#_c_560_n N_VGND_c_782_n 0.00372618f $X=6.45 $Y=1.26 $X2=0
+ $Y2=0
cc_405 N_A_917_107#_c_561_n N_VGND_c_782_n 0.0344812f $X=5.05 $Y=0.745 $X2=0
+ $Y2=0
cc_406 N_A_917_107#_c_563_n N_VGND_c_782_n 0.00583674f $X=5.44 $Y=1.26 $X2=0
+ $Y2=0
cc_407 N_A_917_107#_c_621_n N_VGND_c_782_n 0.00944702f $X=6.615 $Y=1.28 $X2=0
+ $Y2=0
cc_408 N_A_917_107#_c_564_n N_VGND_c_782_n 0.0070366f $X=6.835 $Y=1.435 $X2=0
+ $Y2=0
cc_409 N_RESET_B_c_661_n N_VPWR_c_703_n 0.0525158f $X=7.68 $Y=1.77 $X2=0 $Y2=0
cc_410 N_RESET_B_c_661_n N_VPWR_c_706_n 0.00584154f $X=7.68 $Y=1.77 $X2=0 $Y2=0
cc_411 RESET_B N_VGND_c_780_n 0.0363473f $X=7.835 $Y=0.84 $X2=0 $Y2=0
cc_412 N_RESET_B_M1003_g N_VGND_c_780_n 0.011881f $X=8.02 $Y=0.745 $X2=0 $Y2=0
cc_413 RESET_B N_VGND_c_782_n 0.0309023f $X=7.835 $Y=0.84 $X2=0 $Y2=0
cc_414 N_RESET_B_M1003_g N_VGND_c_782_n 0.0227308f $X=8.02 $Y=0.745 $X2=0 $Y2=0
cc_415 RESET_B A_1512_107# 0.00149154f $X=7.835 $Y=0.84 $X2=0 $Y2=0
cc_416 N_VPWR_c_706_n Q 0.0837f $X=8.405 $Y=3.59 $X2=0.24 $Y2=4.07
cc_417 N_VPWR_c_703_n N_Q_c_761_n 0.0893061f $X=8.12 $Y=2.47 $X2=0 $Y2=0
cc_418 N_Q_c_755_n N_VGND_c_780_n 0.0459558f $X=9.305 $Y=0.66 $X2=0 $Y2=0
cc_419 N_Q_c_755_n N_VGND_c_782_n 0.0340863f $X=9.305 $Y=0.66 $X2=0 $Y2=0
cc_420 N_VGND_c_782_n A_775_107# 0.00226189f $X=8.775 $Y=0.48 $X2=0 $Y2=0
cc_421 N_VGND_c_778_n A_1096_107# 0.00493749f $X=6.38 $Y=0.48 $X2=0 $Y2=0
cc_422 N_VGND_c_782_n A_1096_107# 8.85468e-19 $X=8.775 $Y=0.48 $X2=0 $Y2=0
cc_423 N_VGND_c_782_n A_1512_107# 0.00184558f $X=8.775 $Y=0.48 $X2=0 $Y2=0
