* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__einvp_1 A TE VGND VNB VPB VPWR Z
M1000 Z A a_413_443# VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=5.4e+11p ps=3.72e+06u
M1001 a_413_123# TE VGND VNB nhv w=750000u l=500000u
+  ad=2.7e+11p pd=2.22e+06u as=3.5865e+11p ps=2.76e+06u
M1002 VPWR TE a_30_189# VPB phv w=750000u l=500000u
+  ad=4.9875e+11p pd=3.76e+06u as=2.1375e+11p ps=2.07e+06u
M1003 Z A a_413_123# VNB nhv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
M1004 a_413_443# a_30_189# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND TE a_30_189# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
.ends
