* File: sky130_fd_sc_hvl__lsbufhv2hv_lh_1.pxi.spice
* Created: Fri Aug 28 09:36:43 2020
* 
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%VNB N_VNB_M1011_b VNB VNB N_VNB_c_6_p
+ N_VNB_c_38_p VNB VNB PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%VNB
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%VPB N_VPB_X16_noxref_D1 N_VPB_M1003_b VPB
+ N_VPB_c_78_n N_VPB_c_87_p N_VPB_c_79_n VPB
+ PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%VPB
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%LOWHVPWR N_LOWHVPWR_M1014_d
+ N_LOWHVPWR_M1014_b N_LOWHVPWR_c_138_n LOWHVPWR N_LOWHVPWR_c_145_p LOWHVPWR
+ PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%LOWHVPWR
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A N_A_c_184_n N_A_M1011_g N_A_M1014_g
+ N_A_c_187_n A A N_A_c_189_n PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A_626_141# N_A_626_141#_M1011_s
+ N_A_626_141#_M1014_s N_A_626_141#_c_217_n N_A_626_141#_M1000_g
+ N_A_626_141#_M1006_g N_A_626_141#_M1009_g N_A_626_141#_c_219_n
+ N_A_626_141#_M1002_g N_A_626_141#_c_220_n N_A_626_141#_M1007_g
+ N_A_626_141#_c_221_n N_A_626_141#_M1013_g N_A_626_141#_c_222_n
+ N_A_626_141#_c_223_n N_A_626_141#_c_224_n N_A_626_141#_c_225_n
+ N_A_626_141#_c_226_n N_A_626_141#_c_227_n N_A_626_141#_c_254_n
+ N_A_626_141#_c_228_n PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A_626_141#
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A_847_1221# N_A_847_1221#_M1000_d
+ N_A_847_1221#_M1007_d N_A_847_1221#_M1005_s N_A_847_1221#_c_315_n
+ N_A_847_1221#_M1003_g N_A_847_1221#_c_318_n N_A_847_1221#_c_328_n
+ N_A_847_1221#_c_330_n N_A_847_1221#_c_312_n N_A_847_1221#_c_334_n
+ N_A_847_1221#_c_313_n N_A_847_1221#_c_321_n N_A_847_1221#_c_314_n
+ N_A_847_1221#_c_323_n PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A_847_1221#
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A_935_141# N_A_935_141#_M1006_d
+ N_A_935_141#_M1009_d N_A_935_141#_c_373_n N_A_935_141#_M1008_g
+ N_A_935_141#_c_374_n N_A_935_141#_M1010_g N_A_935_141#_c_375_n
+ N_A_935_141#_M1012_g N_A_935_141#_c_376_n N_A_935_141#_M1015_g
+ N_A_935_141#_c_377_n N_A_935_141#_c_386_n N_A_935_141#_c_378_n
+ N_A_935_141#_c_379_n N_A_935_141#_c_380_n N_A_935_141#_c_392_n
+ N_A_935_141#_c_381_n N_A_935_141#_c_394_n N_A_935_141#_c_382_n
+ N_A_935_141#_c_383_n PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A_935_141#
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A_1353_107# N_A_1353_107#_M1008_s
+ N_A_1353_107#_M1012_s N_A_1353_107#_M1003_s N_A_1353_107#_c_450_n
+ N_A_1353_107#_M1001_g N_A_1353_107#_M1004_g N_A_1353_107#_M1005_g
+ N_A_1353_107#_c_461_n N_A_1353_107#_c_453_n N_A_1353_107#_c_494_n
+ N_A_1353_107#_c_474_n N_A_1353_107#_c_454_n N_A_1353_107#_c_465_n
+ N_A_1353_107#_c_466_n N_A_1353_107#_c_467_n N_A_1353_107#_c_500_n
+ N_A_1353_107#_c_455_n N_A_1353_107#_c_470_n N_A_1353_107#_c_471_n
+ N_A_1353_107#_c_472_n N_A_1353_107#_c_456_n
+ PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A_1353_107#
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%VPWR N_VPWR_M1003_d N_VPWR_M1005_d
+ N_VPWR_c_540_n N_VPWR_c_543_n VPWR VPWR N_VPWR_c_544_n N_VPWR_c_547_n
+ N_VPWR_c_538_n N_VPWR_c_539_n VPWR VPWR
+ PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%VPWR
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%X N_X_M1004_d N_X_M1001_d X X X X X
+ N_X_c_605_n PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%X
x_PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%VGND N_VGND_M1000_s N_VGND_M1011_d
+ N_VGND_M1002_s N_VGND_M1008_d N_VGND_M1013_s N_VGND_M1010_d N_VGND_M1015_d
+ N_VGND_M1004_s N_VGND_c_618_n N_VGND_c_620_n N_VGND_c_622_n N_VGND_c_624_n
+ N_VGND_c_626_n N_VGND_c_628_n N_VGND_c_630_n N_VGND_c_632_n N_VGND_c_634_n
+ N_VGND_c_636_n VGND VGND N_VGND_c_638_n N_VGND_c_639_n N_VGND_c_666_n
+ N_VGND_c_640_n N_VGND_c_641_n N_VGND_c_705_n N_VGND_c_642_n N_VGND_c_643_n
+ N_VGND_c_645_n N_VGND_c_647_n VGND VGND
+ PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%VGND
cc_1 N_VNB_M1011_b N_VPB_c_78_n 0.0021751f $X=-0.33 $Y=-0.265 $X2=0.24 $Y2=4.07
cc_2 N_VNB_M1011_b N_VPB_c_79_n 0.0836863f $X=-0.33 $Y=-0.265 $X2=10.32 $Y2=4.07
cc_3 N_VNB_M1011_b LOWHVPWR 0.159673f $X=-0.33 $Y=-0.265 $X2=0.24 $Y2=4.07
cc_4 N_VNB_M1011_b N_A_c_184_n 0.0408743f $X=-0.33 $Y=-0.265 $X2=0 $Y2=3.985
cc_5 N_VNB_M1011_b N_A_M1011_g 0.0603069f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_c_6_p N_A_M1011_g 0.00133274f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_7 N_VNB_M1011_b N_A_c_187_n 0.020992f $X=-0.33 $Y=-0.265 $X2=0 $Y2=3.955
cc_8 N_VNB_M1011_b A 0.0248803f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_M1011_b N_A_c_189_n 0.0818371f $X=-0.33 $Y=-0.265 $X2=0.24 $Y2=4.07
cc_10 N_VNB_M1011_b N_A_626_141#_c_217_n 0.0411781f $X=-0.33 $Y=-0.265 $X2=-0.33
+ $Y2=1.885
cc_11 N_VNB_M1011_b N_A_626_141#_M1006_g 0.0575209f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1011_b N_A_626_141#_c_219_n 0.0358616f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1011_b N_A_626_141#_c_220_n 0.0358616f $X=-0.33 $Y=-0.265 $X2=8.88
+ $Y2=4.07
cc_14 N_VNB_M1011_b N_A_626_141#_c_221_n 0.041717f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_15 N_VNB_M1011_b N_A_626_141#_c_222_n 0.042392f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_16 N_VNB_M1011_b N_A_626_141#_c_223_n 0.0555285f $X=-0.33 $Y=-0.265 $X2=8.88
+ $Y2=4.07
cc_17 N_VNB_M1011_b N_A_626_141#_c_224_n 0.010074f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1011_b N_A_626_141#_c_225_n 0.0399436f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_19 N_VNB_M1011_b N_A_626_141#_c_226_n 0.027992f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_20 N_VNB_M1011_b N_A_626_141#_c_227_n 0.0588454f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_21 N_VNB_M1011_b N_A_626_141#_c_228_n 0.334761f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_22 N_VNB_M1011_b N_A_847_1221#_c_312_n 0.00309886f $X=-0.33 $Y=-0.265
+ $X2=10.32 $Y2=4.07
cc_23 N_VNB_M1011_b N_A_847_1221#_c_313_n 0.0459015f $X=-0.33 $Y=-0.265 $X2=4.8
+ $Y2=4.068
cc_24 N_VNB_M1011_b N_A_847_1221#_c_314_n 0.0134401f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_25 N_VNB_M1011_b N_A_935_141#_c_373_n 0.0396454f $X=-0.33 $Y=-0.265 $X2=-0.33
+ $Y2=1.885
cc_26 N_VNB_M1011_b N_A_935_141#_c_374_n 0.0358616f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_27 N_VNB_M1011_b N_A_935_141#_c_375_n 0.0358616f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_28 N_VNB_M1011_b N_A_935_141#_c_376_n 0.202798f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_29 N_VNB_M1011_b N_A_935_141#_c_377_n 0.0203873f $X=-0.33 $Y=-0.265 $X2=8.88
+ $Y2=4.07
cc_30 N_VNB_M1011_b N_A_935_141#_c_378_n 0.0361133f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_31 N_VNB_M1011_b N_A_935_141#_c_379_n 0.00730387f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_32 N_VNB_M1011_b N_A_935_141#_c_380_n 0.00390048f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_33 N_VNB_M1011_b N_A_935_141#_c_381_n 0.0217586f $X=-0.33 $Y=-0.265 $X2=4.8
+ $Y2=4.068
cc_34 N_VNB_M1011_b N_A_935_141#_c_382_n 0.00739552f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_35 N_VNB_M1011_b N_A_935_141#_c_383_n 0.0823775f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_36 N_VNB_M1011_b N_A_1353_107#_c_450_n 0.0459087f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_37 N_VNB_M1011_b N_A_1353_107#_M1004_g 0.0793374f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_38 N_VNB_c_38_p N_A_1353_107#_M1004_g 0.00161049f $X=10.32 $Y=8.14 $X2=0
+ $Y2=0
cc_39 N_VNB_M1011_b N_A_1353_107#_c_453_n 0.024481f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_40 N_VNB_M1011_b N_A_1353_107#_c_454_n 0.00643837f $X=-0.33 $Y=-0.265
+ $X2=8.88 $Y2=4.07
cc_41 N_VNB_M1011_b N_A_1353_107#_c_455_n 0.0133586f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_42 N_VNB_M1011_b N_A_1353_107#_c_456_n 0.036449f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_M1011_b N_VPWR_c_538_n 0.098711f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_44 N_VNB_M1011_b N_VPWR_c_539_n 0.275264f $X=-0.33 $Y=-0.265 $X2=4.8 $Y2=4.07
cc_45 N_VNB_M1011_b N_X_c_605_n 0.0630727f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_46 N_VNB_c_38_p N_X_c_605_n 7.98897e-19 $X=10.32 $Y=8.14 $X2=0 $Y2=0
cc_47 N_VNB_M1011_b N_VGND_c_618_n 0.0718145f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_48 N_VNB_c_38_p N_VGND_c_618_n 0.00332742f $X=10.32 $Y=8.14 $X2=10.32
+ $Y2=4.07
cc_49 N_VNB_M1011_b N_VGND_c_620_n 0.0481389f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_50 N_VNB_c_38_p N_VGND_c_620_n 0.00198821f $X=10.32 $Y=8.14 $X2=10.32
+ $Y2=4.07
cc_51 N_VNB_M1011_b N_VGND_c_622_n 0.135335f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_52 N_VNB_c_6_p N_VGND_c_622_n 0.00514627f $X=10.32 $Y=0 $X2=10.32 $Y2=4.07
cc_53 N_VNB_M1011_b N_VGND_c_624_n 0.0495906f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_54 N_VNB_c_6_p N_VGND_c_624_n 0.00198821f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_55 N_VNB_M1011_b N_VGND_c_626_n 0.119953f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_56 N_VNB_c_38_p N_VGND_c_626_n 0.00531562f $X=10.32 $Y=8.14 $X2=0.24 $Y2=4.07
cc_57 N_VNB_M1011_b N_VGND_c_628_n 0.0718145f $X=-0.33 $Y=-0.265 $X2=4.8
+ $Y2=4.07
cc_58 N_VNB_c_6_p N_VGND_c_628_n 0.00332742f $X=10.32 $Y=0 $X2=4.8 $Y2=4.07
cc_59 N_VNB_M1011_b N_VGND_c_630_n 0.119953f $X=-0.33 $Y=-0.265 $X2=5.28
+ $Y2=4.07
cc_60 N_VNB_c_6_p N_VGND_c_630_n 0.00531562f $X=10.32 $Y=0 $X2=5.28 $Y2=4.07
cc_61 N_VNB_M1011_b N_VGND_c_632_n 0.0443345f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_62 N_VNB_c_38_p N_VGND_c_632_n 0.00198821f $X=10.32 $Y=8.14 $X2=0 $Y2=0
cc_63 N_VNB_M1011_b N_VGND_c_634_n 0.0459379f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_64 N_VNB_c_6_p N_VGND_c_634_n 0.00198821f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_65 N_VNB_M1011_b N_VGND_c_636_n 0.0443345f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_66 N_VNB_c_6_p N_VGND_c_636_n 0.00198821f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_67 N_VNB_M1011_b N_VGND_c_638_n 0.0774259f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_68 N_VNB_M1011_b N_VGND_c_639_n 0.00698685f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_69 N_VNB_M1011_b N_VGND_c_640_n 0.0421704f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_70 N_VNB_M1011_b N_VGND_c_641_n 0.0682032f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_71 N_VNB_M1011_b N_VGND_c_642_n 0.0734992f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_72 N_VNB_M1011_b N_VGND_c_643_n 0.338665f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_73 N_VNB_c_6_p N_VGND_c_643_n 1.11411f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_74 N_VNB_M1011_b N_VGND_c_645_n 0.0680644f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_75 N_VNB_c_38_p N_VGND_c_645_n 0.00159492f $X=10.32 $Y=8.14 $X2=0 $Y2=0
cc_76 N_VNB_M1011_b N_VGND_c_647_n 0.394369f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_77 N_VNB_c_38_p N_VGND_c_647_n 1.11838f $X=10.32 $Y=8.14 $X2=0 $Y2=0
cc_78 N_VPB_c_79_n N_LOWHVPWR_M1014_b 0.0291872f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_79 N_VPB_c_79_n N_LOWHVPWR_c_138_n 0.0595146f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_80 N_VPB_X16_noxref_D1 LOWHVPWR 0.050189f $X=-0.33 $Y=1.885 $X2=0.24 $Y2=0
cc_81 N_VPB_M1003_b LOWHVPWR 0.0690009f $X=7.27 $Y=2.465 $X2=0.24 $Y2=0
cc_82 N_VPB_c_79_n N_A_626_141#_c_223_n 0.0312993f $X=10.32 $Y=4.07 $X2=10.32
+ $Y2=8.14
cc_83 N_VPB_M1003_b N_A_847_1221#_c_315_n 0.0226258f $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_84 N_VPB_M1003_b N_A_847_1221#_M1003_g 0.0854755f $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_85 N_VPB_c_87_p N_A_847_1221#_M1003_g 0.00484292f $X=10.32 $Y=4.07 $X2=0
+ $Y2=0
cc_86 N_VPB_M1003_b N_A_847_1221#_c_318_n 0.0967283f $X=7.27 $Y=2.465 $X2=0.24
+ $Y2=0
cc_87 N_VPB_c_79_n N_A_847_1221#_c_318_n 0.00607296f $X=10.32 $Y=4.07 $X2=0.24
+ $Y2=0
cc_88 N_VPB_M1003_b N_A_847_1221#_c_313_n 0.059422f $X=7.27 $Y=2.465 $X2=0 $Y2=0
cc_89 N_VPB_M1003_b N_A_847_1221#_c_321_n 0.0598451f $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_90 N_VPB_c_79_n N_A_847_1221#_c_321_n 0.0256052f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_91 N_VPB_M1003_b N_A_847_1221#_c_323_n 0.00754345f $X=7.27 $Y=2.465 $X2=4.8
+ $Y2=0.058
cc_92 N_VPB_c_79_n N_A_847_1221#_c_323_n 0.0110089f $X=10.32 $Y=4.07 $X2=4.8
+ $Y2=0.058
cc_93 N_VPB_M1003_b N_A_935_141#_c_376_n 0.0449607f $X=7.27 $Y=2.465 $X2=0.24
+ $Y2=0
cc_94 N_VPB_M1003_b N_A_1353_107#_c_450_n 0.0190575f $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_95 N_VPB_M1003_b N_A_1353_107#_M1001_g 0.0611611f $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_96 N_VPB_c_87_p N_A_1353_107#_M1001_g 0.0175739f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_97 N_VPB_c_79_n N_A_1353_107#_M1001_g 0.00970178f $X=10.32 $Y=4.07 $X2=0
+ $Y2=0
cc_98 N_VPB_M1003_b N_A_1353_107#_c_461_n 0.0948383f $X=7.27 $Y=2.465 $X2=10.32
+ $Y2=0
cc_99 N_VPB_c_87_p N_A_1353_107#_c_461_n 0.00778503f $X=10.32 $Y=4.07 $X2=10.32
+ $Y2=0
cc_100 N_VPB_c_79_n N_A_1353_107#_c_461_n 0.00964562f $X=10.32 $Y=4.07 $X2=10.32
+ $Y2=0
cc_101 N_VPB_M1003_b N_A_1353_107#_c_453_n 0.0024481f $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_102 N_VPB_M1003_b N_A_1353_107#_c_465_n 0.0155783f $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_103 N_VPB_M1003_b N_A_1353_107#_c_466_n 0.0216195f $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_104 N_VPB_M1003_b N_A_1353_107#_c_467_n 0.0252804f $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_105 N_VPB_c_87_p N_A_1353_107#_c_467_n 0.0120574f $X=10.32 $Y=4.07 $X2=0
+ $Y2=0
cc_106 N_VPB_c_79_n N_A_1353_107#_c_467_n 0.0244469f $X=10.32 $Y=4.07 $X2=0
+ $Y2=0
cc_107 N_VPB_M1003_b N_A_1353_107#_c_470_n 4.76607e-19 $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_108 N_VPB_M1003_b N_A_1353_107#_c_471_n 0.0263402f $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_109 N_VPB_M1003_b N_A_1353_107#_c_472_n 0.128346f $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_VPB_M1003_b N_A_1353_107#_c_456_n 0.00270883f $X=7.27 $Y=2.465 $X2=0
+ $Y2=0
cc_111 N_VPB_M1003_b N_VPWR_c_540_n 0.00227194f $X=7.27 $Y=2.465 $X2=0 $Y2=0
cc_112 N_VPB_c_87_p N_VPWR_c_540_n 0.028048f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_113 N_VPB_c_79_n N_VPWR_c_540_n 0.0020337f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_114 N_VPB_M1003_b N_VPWR_c_543_n 0.0239839f $X=7.27 $Y=2.465 $X2=-0.33
+ $Y2=-0.265
cc_115 N_VPB_M1003_b N_VPWR_c_544_n 0.00121452f $X=7.27 $Y=2.465 $X2=0.24 $Y2=0
cc_116 N_VPB_c_87_p N_VPWR_c_544_n 0.019481f $X=10.32 $Y=4.07 $X2=0.24 $Y2=0
cc_117 N_VPB_c_79_n N_VPWR_c_544_n 0.00152922f $X=10.32 $Y=4.07 $X2=0.24 $Y2=0
cc_118 N_VPB_M1003_b N_VPWR_c_547_n 0.0562562f $X=7.27 $Y=2.465 $X2=10.32 $Y2=0
cc_119 N_VPB_c_87_p N_VPWR_c_547_n 0.0254284f $X=10.32 $Y=4.07 $X2=10.32 $Y2=0
cc_120 N_VPB_c_79_n N_VPWR_c_547_n 0.00166879f $X=10.32 $Y=4.07 $X2=10.32 $Y2=0
cc_121 N_VPB_X16_noxref_D1 N_VPWR_c_538_n 0.0336658f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_122 N_VPB_M1003_b N_VPWR_c_538_n 0.0499984f $X=7.27 $Y=2.465 $X2=0 $Y2=0
cc_123 N_VPB_c_78_n N_VPWR_c_538_n 0.00613319f $X=0.24 $Y=4.07 $X2=0 $Y2=0
cc_124 N_VPB_c_87_p N_VPWR_c_538_n 0.0118549f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_125 N_VPB_c_79_n N_VPWR_c_538_n 1.10385f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_126 N_VPB_X16_noxref_D1 N_VPWR_c_539_n 0.0565882f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_127 N_VPB_M1003_b N_VPWR_c_539_n 0.0402136f $X=7.27 $Y=2.465 $X2=0 $Y2=0
cc_128 N_VPB_c_78_n N_VPWR_c_539_n 0.00613319f $X=0.24 $Y=4.07 $X2=0 $Y2=0
cc_129 N_VPB_c_87_p N_VPWR_c_539_n 0.00850276f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_130 N_VPB_c_79_n N_VPWR_c_539_n 1.11909f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_131 N_VPB_M1003_b N_X_c_605_n 0.0670968f $X=7.27 $Y=2.465 $X2=0 $Y2=0
cc_132 N_VPB_c_87_p N_X_c_605_n 0.0158392f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_133 N_VPB_c_79_n N_X_c_605_n 0.00101808f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_134 N_LOWHVPWR_M1014_b N_A_c_184_n 0.0233928f $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_135 N_LOWHVPWR_M1014_b N_A_M1014_g 0.0583521f $X=2.8 $Y=2.015 $X2=-0.33
+ $Y2=-0.265
cc_136 N_LOWHVPWR_c_138_n N_A_M1014_g 0.00724845f $X=4.695 $Y=3.52 $X2=-0.33
+ $Y2=-0.265
cc_137 LOWHVPWR N_A_M1014_g 0.0182732f $X=0.07 $Y=3.02 $X2=-0.33 $Y2=-0.265
cc_138 N_LOWHVPWR_c_145_p N_A_M1014_g 0.0382962f $X=4.035 $Y=2.49 $X2=-0.33
+ $Y2=-0.265
cc_139 N_LOWHVPWR_M1014_b N_A_c_187_n 0.00146233f $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_140 N_LOWHVPWR_M1014_b N_A_c_189_n 0.00602715f $X=2.8 $Y=2.015 $X2=0.24 $Y2=0
cc_141 N_LOWHVPWR_M1014_b N_A_626_141#_M1009_g 0.0610725f $X=2.8 $Y=2.015
+ $X2=0.24 $Y2=0
cc_142 N_LOWHVPWR_c_138_n N_A_626_141#_M1009_g 0.0150117f $X=4.695 $Y=3.52
+ $X2=0.24 $Y2=0
cc_143 LOWHVPWR N_A_626_141#_M1009_g 0.0203751f $X=0.07 $Y=3.02 $X2=0.24 $Y2=0
cc_144 N_LOWHVPWR_c_145_p N_A_626_141#_M1009_g 0.0392499f $X=4.035 $Y=2.49
+ $X2=0.24 $Y2=0
cc_145 N_LOWHVPWR_M1014_b N_A_626_141#_c_223_n 0.0881397f $X=2.8 $Y=2.015
+ $X2=10.32 $Y2=8.14
cc_146 N_LOWHVPWR_c_138_n N_A_626_141#_c_223_n 0.0507377f $X=4.695 $Y=3.52
+ $X2=10.32 $Y2=8.14
cc_147 LOWHVPWR N_A_626_141#_c_223_n 0.0478141f $X=0.07 $Y=3.02 $X2=10.32
+ $Y2=8.14
cc_148 N_LOWHVPWR_c_145_p N_A_626_141#_c_223_n 0.0452275f $X=4.035 $Y=2.49
+ $X2=10.32 $Y2=8.14
cc_149 N_LOWHVPWR_c_145_p N_A_626_141#_c_224_n 0.0294514f $X=4.035 $Y=2.49 $X2=0
+ $Y2=0
cc_150 N_LOWHVPWR_M1014_b N_A_626_141#_c_225_n 0.00649522f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_151 LOWHVPWR N_A_847_1221#_M1003_g 0.0159233f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_152 LOWHVPWR N_A_847_1221#_c_318_n 0.00117082f $X=0.07 $Y=3.02 $X2=0.24 $Y2=0
cc_153 LOWHVPWR N_A_847_1221#_c_323_n 0.00448365f $X=0.07 $Y=3.02 $X2=4.8
+ $Y2=0.058
cc_154 LOWHVPWR N_A_935_141#_c_376_n 0.00131056f $X=0.07 $Y=3.02 $X2=0.24 $Y2=0
cc_155 N_LOWHVPWR_M1014_b N_A_935_141#_c_386_n 0.0255441f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_156 N_LOWHVPWR_c_138_n N_A_935_141#_c_386_n 0.00641004f $X=4.695 $Y=3.52
+ $X2=0 $Y2=0
cc_157 LOWHVPWR N_A_935_141#_c_386_n 0.0336116f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_158 N_LOWHVPWR_c_145_p N_A_935_141#_c_386_n 0.028744f $X=4.035 $Y=2.49 $X2=0
+ $Y2=0
cc_159 N_LOWHVPWR_M1014_b N_A_935_141#_c_380_n 0.0190927f $X=2.8 $Y=2.015
+ $X2=0.24 $Y2=8.14
cc_160 LOWHVPWR N_A_935_141#_c_380_n 0.012615f $X=0.07 $Y=3.02 $X2=0.24 $Y2=8.14
cc_161 N_LOWHVPWR_M1014_b N_A_935_141#_c_392_n 0.00750794f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_162 N_LOWHVPWR_c_145_p N_A_935_141#_c_392_n 0.00751668f $X=4.035 $Y=2.49
+ $X2=0 $Y2=0
cc_163 LOWHVPWR N_A_935_141#_c_394_n 0.0297219f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_164 LOWHVPWR N_A_935_141#_c_382_n 0.0125456f $X=0.07 $Y=3.02 $X2=4.8 $Y2=0
cc_165 LOWHVPWR N_A_935_141#_c_383_n 0.037513f $X=0.07 $Y=3.02 $X2=4.8 $Y2=0.058
cc_166 LOWHVPWR N_A_1353_107#_c_474_n 0.0200805f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_167 LOWHVPWR N_A_1353_107#_c_454_n 0.0116369f $X=0.07 $Y=3.02 $X2=10.32
+ $Y2=8.14
cc_168 LOWHVPWR N_A_1353_107#_c_466_n 0.05867f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_169 LOWHVPWR N_A_1353_107#_c_467_n 0.0168006f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_170 LOWHVPWR N_A_1353_107#_c_470_n 0.00268926f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_171 LOWHVPWR N_VPWR_c_547_n 0.0666751f $X=0.07 $Y=3.02 $X2=10.32 $Y2=0
cc_172 N_LOWHVPWR_M1014_b N_VPWR_c_538_n 0.0196315f $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_173 N_LOWHVPWR_c_138_n N_VPWR_c_538_n 0.0891245f $X=4.695 $Y=3.52 $X2=0 $Y2=0
cc_174 LOWHVPWR N_VPWR_c_538_n 1.10321f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_175 N_LOWHVPWR_c_145_p N_VPWR_c_538_n 4.74994e-19 $X=4.035 $Y=2.49 $X2=0
+ $Y2=0
cc_176 N_LOWHVPWR_c_138_n N_VPWR_c_539_n 0.00618556f $X=4.695 $Y=3.52 $X2=0
+ $Y2=0
cc_177 N_A_M1011_g N_A_626_141#_M1006_g 0.0227397f $X=3.645 $Y=1.08 $X2=0
+ $Y2=8.025
cc_178 N_A_M1014_g N_A_626_141#_M1009_g 0.0227397f $X=3.645 $Y=2.72 $X2=0.24
+ $Y2=0
cc_179 N_A_c_184_n N_A_626_141#_c_222_n 0.00929641f $X=3.395 $Y=1.87 $X2=0.24
+ $Y2=8.14
cc_180 N_A_M1011_g N_A_626_141#_c_222_n 0.0345799f $X=3.645 $Y=1.08 $X2=0.24
+ $Y2=8.14
cc_181 N_A_c_187_n N_A_626_141#_c_222_n 0.00183495f $X=3.645 $Y=1.87 $X2=0.24
+ $Y2=8.14
cc_182 A N_A_626_141#_c_222_n 0.0113411f $X=2.555 $Y=1.58 $X2=0.24 $Y2=8.14
cc_183 N_A_c_189_n N_A_626_141#_c_222_n 0.00167153f $X=2.66 $Y=1.695 $X2=0.24
+ $Y2=8.14
cc_184 N_A_c_184_n N_A_626_141#_c_223_n 0.00929641f $X=3.395 $Y=1.87 $X2=10.32
+ $Y2=8.14
cc_185 N_A_M1014_g N_A_626_141#_c_223_n 0.0421868f $X=3.645 $Y=2.72 $X2=10.32
+ $Y2=8.14
cc_186 N_A_c_187_n N_A_626_141#_c_223_n 0.00183495f $X=3.645 $Y=1.87 $X2=10.32
+ $Y2=8.14
cc_187 A N_A_626_141#_c_223_n 0.0108046f $X=2.555 $Y=1.58 $X2=10.32 $Y2=8.14
cc_188 N_A_c_189_n N_A_626_141#_c_223_n 0.00157601f $X=2.66 $Y=1.695 $X2=10.32
+ $Y2=8.14
cc_189 N_A_c_187_n N_A_626_141#_c_224_n 0.0494497f $X=3.645 $Y=1.87 $X2=0 $Y2=0
cc_190 N_A_c_187_n N_A_626_141#_c_225_n 0.0227397f $X=3.645 $Y=1.87 $X2=0 $Y2=0
cc_191 N_A_c_184_n N_A_626_141#_c_254_n 0.0119558f $X=3.395 $Y=1.87 $X2=4.8
+ $Y2=8.14
cc_192 N_A_c_187_n N_A_626_141#_c_254_n 5.88527e-19 $X=3.645 $Y=1.87 $X2=4.8
+ $Y2=8.14
cc_193 A N_A_626_141#_c_254_n 0.0131201f $X=2.555 $Y=1.58 $X2=4.8 $Y2=8.14
cc_194 N_A_M1014_g N_VPWR_c_538_n 8.98934e-19 $X=3.645 $Y=2.72 $X2=0 $Y2=0
cc_195 N_A_M1011_g N_VGND_c_639_n 0.0416092f $X=3.645 $Y=1.08 $X2=0 $Y2=0
cc_196 N_A_M1011_g N_VGND_c_643_n 0.0204436f $X=3.645 $Y=1.08 $X2=0 $Y2=0
cc_197 N_A_626_141#_c_217_n N_A_847_1221#_c_328_n 0.0381272f $X=3.985 $Y=5.995
+ $X2=0 $Y2=0
cc_198 N_A_626_141#_c_219_n N_A_847_1221#_c_328_n 0.0401197f $X=4.765 $Y=5.995
+ $X2=0 $Y2=0
cc_199 N_A_626_141#_c_227_n N_A_847_1221#_c_330_n 0.084463f $X=5.495 $Y=5.33
+ $X2=0 $Y2=0
cc_200 N_A_626_141#_c_228_n N_A_847_1221#_c_330_n 0.0948653f $X=5.545 $Y=5.58
+ $X2=0 $Y2=0
cc_201 N_A_626_141#_c_227_n N_A_847_1221#_c_312_n 0.0276921f $X=5.495 $Y=5.33
+ $X2=0 $Y2=0
cc_202 N_A_626_141#_c_228_n N_A_847_1221#_c_312_n 0.0287562f $X=5.545 $Y=5.58
+ $X2=0 $Y2=0
cc_203 N_A_626_141#_c_220_n N_A_847_1221#_c_334_n 0.0401197f $X=5.545 $Y=5.995
+ $X2=0.24 $Y2=8.14
cc_204 N_A_626_141#_c_221_n N_A_847_1221#_c_334_n 0.0401197f $X=6.325 $Y=5.995
+ $X2=0.24 $Y2=8.14
cc_205 N_A_626_141#_c_228_n N_A_847_1221#_c_313_n 0.059011f $X=5.545 $Y=5.58
+ $X2=0 $Y2=0
cc_206 N_A_626_141#_c_228_n N_A_847_1221#_c_314_n 0.0175374f $X=5.545 $Y=5.58
+ $X2=0 $Y2=0
cc_207 N_A_626_141#_M1006_g N_A_935_141#_c_377_n 0.0121585f $X=4.425 $Y=1.08
+ $X2=0 $Y2=0
cc_208 N_A_626_141#_M1009_g N_A_935_141#_c_386_n 0.0153965f $X=4.425 $Y=2.72
+ $X2=0 $Y2=0
cc_209 N_A_626_141#_M1006_g N_A_935_141#_c_379_n 0.00845053f $X=4.425 $Y=1.08
+ $X2=0.24 $Y2=8.14
cc_210 N_A_626_141#_c_224_n N_A_935_141#_c_379_n 0.0113212f $X=4.68 $Y=1.87
+ $X2=0.24 $Y2=8.14
cc_211 N_A_626_141#_c_225_n N_A_935_141#_c_379_n 0.00393092f $X=4.68 $Y=1.87
+ $X2=0.24 $Y2=8.14
cc_212 N_A_626_141#_M1009_g N_A_935_141#_c_392_n 0.0163873f $X=4.425 $Y=2.72
+ $X2=0 $Y2=0
cc_213 N_A_626_141#_c_224_n N_A_935_141#_c_392_n 0.0160252f $X=4.68 $Y=1.87
+ $X2=0 $Y2=0
cc_214 N_A_626_141#_c_225_n N_A_935_141#_c_392_n 0.00415632f $X=4.68 $Y=1.87
+ $X2=0 $Y2=0
cc_215 N_A_626_141#_M1006_g N_A_935_141#_c_381_n 0.0058909f $X=4.425 $Y=1.08
+ $X2=0 $Y2=0
cc_216 N_A_626_141#_M1009_g N_A_935_141#_c_381_n 0.00280396f $X=4.425 $Y=2.72
+ $X2=0 $Y2=0
cc_217 N_A_626_141#_c_224_n N_A_935_141#_c_381_n 0.00944185f $X=4.68 $Y=1.87
+ $X2=0 $Y2=0
cc_218 N_A_626_141#_c_225_n N_A_935_141#_c_381_n 0.00407226f $X=4.68 $Y=1.87
+ $X2=0 $Y2=0
cc_219 N_A_626_141#_M1009_g N_A_935_141#_c_382_n 5.63146e-19 $X=4.425 $Y=2.72
+ $X2=4.8 $Y2=0
cc_220 N_A_626_141#_c_223_n N_VPWR_c_538_n 0.0387554f $X=3.255 $Y=2.49 $X2=0
+ $Y2=0
cc_221 N_A_626_141#_c_223_n N_VPWR_c_539_n 0.0625354f $X=3.255 $Y=2.49 $X2=0
+ $Y2=0
cc_222 N_A_626_141#_c_227_n N_VPWR_c_539_n 0.0856203f $X=5.495 $Y=5.33 $X2=0
+ $Y2=0
cc_223 N_A_626_141#_c_228_n N_VPWR_c_539_n 0.0267012f $X=5.545 $Y=5.58 $X2=0
+ $Y2=0
cc_224 N_A_626_141#_c_217_n N_VGND_c_618_n 0.0146836f $X=3.985 $Y=5.995 $X2=0
+ $Y2=0
cc_225 N_A_626_141#_c_219_n N_VGND_c_618_n 0.0146836f $X=4.765 $Y=5.995 $X2=0
+ $Y2=0
cc_226 N_A_626_141#_c_217_n N_VGND_c_620_n 0.0034209f $X=3.985 $Y=5.995 $X2=0
+ $Y2=0
cc_227 N_A_626_141#_M1006_g N_VGND_c_622_n 0.0104183f $X=4.425 $Y=1.08 $X2=0
+ $Y2=0
cc_228 N_A_626_141#_c_220_n N_VGND_c_626_n 0.0146836f $X=5.545 $Y=5.995 $X2=0.24
+ $Y2=8.14
cc_229 N_A_626_141#_c_221_n N_VGND_c_626_n 0.0181045f $X=6.325 $Y=5.995 $X2=0.24
+ $Y2=8.14
cc_230 N_A_626_141#_c_219_n N_VGND_c_632_n 0.00322203f $X=4.765 $Y=5.995 $X2=0
+ $Y2=0
cc_231 N_A_626_141#_c_220_n N_VGND_c_632_n 0.00322203f $X=5.545 $Y=5.995 $X2=0
+ $Y2=0
cc_232 N_A_626_141#_c_217_n N_VGND_c_638_n 0.0628109f $X=3.985 $Y=5.995 $X2=5.28
+ $Y2=8.14
cc_233 N_A_626_141#_c_219_n N_VGND_c_638_n 0.00132352f $X=4.765 $Y=5.995
+ $X2=5.28 $Y2=8.14
cc_234 N_A_626_141#_c_226_n N_VGND_c_638_n 0.00466914f $X=3.42 $Y=5.33 $X2=5.28
+ $Y2=8.14
cc_235 N_A_626_141#_c_227_n N_VGND_c_638_n 0.0166722f $X=5.495 $Y=5.33 $X2=5.28
+ $Y2=8.14
cc_236 N_A_626_141#_M1006_g N_VGND_c_639_n 0.0415973f $X=4.425 $Y=1.08 $X2=0
+ $Y2=0
cc_237 N_A_626_141#_c_222_n N_VGND_c_639_n 0.0373914f $X=3.255 $Y=0.85 $X2=0
+ $Y2=0
cc_238 N_A_626_141#_c_224_n N_VGND_c_639_n 0.0342051f $X=4.68 $Y=1.87 $X2=0
+ $Y2=0
cc_239 N_A_626_141#_c_217_n N_VGND_c_666_n 0.00129485f $X=3.985 $Y=5.995 $X2=0
+ $Y2=0
cc_240 N_A_626_141#_c_219_n N_VGND_c_666_n 0.0567946f $X=4.765 $Y=5.995 $X2=0
+ $Y2=0
cc_241 N_A_626_141#_c_220_n N_VGND_c_666_n 0.0567946f $X=5.545 $Y=5.995 $X2=0
+ $Y2=0
cc_242 N_A_626_141#_c_221_n N_VGND_c_666_n 0.00129485f $X=6.325 $Y=5.995 $X2=0
+ $Y2=0
cc_243 N_A_626_141#_c_228_n N_VGND_c_666_n 0.00272398f $X=5.545 $Y=5.58 $X2=0
+ $Y2=0
cc_244 N_A_626_141#_c_220_n N_VGND_c_641_n 0.00129485f $X=5.545 $Y=5.995 $X2=0
+ $Y2=0
cc_245 N_A_626_141#_c_221_n N_VGND_c_641_n 0.0582646f $X=6.325 $Y=5.995 $X2=0
+ $Y2=0
cc_246 N_A_626_141#_M1006_g N_VGND_c_643_n 0.0204309f $X=4.425 $Y=1.08 $X2=0
+ $Y2=0
cc_247 N_A_626_141#_c_222_n N_VGND_c_643_n 0.0143529f $X=3.255 $Y=0.85 $X2=0
+ $Y2=0
cc_248 N_A_626_141#_c_217_n N_VGND_c_647_n 0.0157032f $X=3.985 $Y=5.995 $X2=0
+ $Y2=0
cc_249 N_A_626_141#_c_219_n N_VGND_c_647_n 0.0157032f $X=4.765 $Y=5.995 $X2=0
+ $Y2=0
cc_250 N_A_626_141#_c_220_n N_VGND_c_647_n 0.0157032f $X=5.545 $Y=5.995 $X2=0
+ $Y2=0
cc_251 N_A_626_141#_c_221_n N_VGND_c_647_n 0.0157032f $X=6.325 $Y=5.995 $X2=0
+ $Y2=0
cc_252 N_A_847_1221#_M1003_g N_A_935_141#_c_376_n 0.072143f $X=8.465 $Y=3.025
+ $X2=0.24 $Y2=0
cc_253 N_A_847_1221#_c_318_n N_A_1353_107#_c_461_n 0.0130406f $X=7.965 $Y=3.77
+ $X2=10.32 $Y2=0
cc_254 N_A_847_1221#_c_321_n N_A_1353_107#_c_461_n 0.0106527f $X=7.825 $Y=4.57
+ $X2=10.32 $Y2=0
cc_255 N_A_847_1221#_c_323_n N_A_1353_107#_c_461_n 5.69156e-19 $X=7.88 $Y=3.77
+ $X2=10.32 $Y2=0
cc_256 N_A_847_1221#_M1003_g N_A_1353_107#_c_474_n 0.00108076f $X=8.465 $Y=3.025
+ $X2=0 $Y2=0
cc_257 N_A_847_1221#_M1003_g N_A_1353_107#_c_465_n 0.0158589f $X=8.465 $Y=3.025
+ $X2=0 $Y2=0
cc_258 N_A_847_1221#_M1003_g N_A_1353_107#_c_466_n 0.0395212f $X=8.465 $Y=3.025
+ $X2=0 $Y2=0
cc_259 N_A_847_1221#_c_318_n N_A_1353_107#_c_466_n 0.00587983f $X=7.965 $Y=3.77
+ $X2=0 $Y2=0
cc_260 N_A_847_1221#_c_323_n N_A_1353_107#_c_466_n 0.0233751f $X=7.88 $Y=3.77
+ $X2=0 $Y2=0
cc_261 N_A_847_1221#_c_315_n N_A_1353_107#_c_467_n 0.0111141f $X=8.13 $Y=3.605
+ $X2=0 $Y2=0
cc_262 N_A_847_1221#_M1003_g N_A_1353_107#_c_467_n 0.0204045f $X=8.465 $Y=3.025
+ $X2=0 $Y2=0
cc_263 N_A_847_1221#_c_318_n N_A_1353_107#_c_467_n 0.0132073f $X=7.965 $Y=3.77
+ $X2=0 $Y2=0
cc_264 N_A_847_1221#_c_321_n N_A_1353_107#_c_467_n 0.0550062f $X=7.825 $Y=4.57
+ $X2=0 $Y2=0
cc_265 N_A_847_1221#_c_323_n N_A_1353_107#_c_467_n 0.0232561f $X=7.88 $Y=3.77
+ $X2=0 $Y2=0
cc_266 N_A_847_1221#_M1003_g N_A_1353_107#_c_470_n 6.44419e-19 $X=8.465 $Y=3.025
+ $X2=0 $Y2=0
cc_267 N_A_847_1221#_c_321_n N_A_1353_107#_c_471_n 0.020235f $X=7.825 $Y=4.57
+ $X2=0 $Y2=0
cc_268 N_A_847_1221#_c_315_n N_VPWR_c_547_n 0.00116463f $X=8.13 $Y=3.605
+ $X2=10.32 $Y2=0
cc_269 N_A_847_1221#_M1003_g N_VPWR_c_547_n 0.0183254f $X=8.465 $Y=3.025
+ $X2=10.32 $Y2=0
cc_270 N_A_847_1221#_c_315_n N_VPWR_c_538_n 0.00472921f $X=8.13 $Y=3.605 $X2=0
+ $Y2=0
cc_271 N_A_847_1221#_M1003_g N_VPWR_c_538_n 0.00782326f $X=8.465 $Y=3.025 $X2=0
+ $Y2=0
cc_272 N_A_847_1221#_c_318_n N_VPWR_c_538_n 0.0105529f $X=7.965 $Y=3.77 $X2=0
+ $Y2=0
cc_273 N_A_847_1221#_c_321_n N_VPWR_c_538_n 2.14811e-19 $X=7.825 $Y=4.57 $X2=0
+ $Y2=0
cc_274 N_A_847_1221#_c_323_n N_VPWR_c_538_n 0.0363684f $X=7.88 $Y=3.77 $X2=0
+ $Y2=0
cc_275 N_A_847_1221#_M1005_s N_VPWR_c_539_n 0.00137624f $X=7.6 $Y=4.425 $X2=0
+ $Y2=0
cc_276 N_A_847_1221#_c_321_n N_VPWR_c_539_n 0.0543355f $X=7.825 $Y=4.57 $X2=0
+ $Y2=0
cc_277 N_A_847_1221#_c_328_n N_VGND_c_618_n 0.0211458f $X=4.375 $Y=6.25 $X2=0
+ $Y2=0
cc_278 N_A_847_1221#_c_334_n N_VGND_c_626_n 0.0211458f $X=5.935 $Y=6.25 $X2=0.24
+ $Y2=8.14
cc_279 N_A_847_1221#_c_328_n N_VGND_c_638_n 0.0686214f $X=4.375 $Y=6.25 $X2=5.28
+ $Y2=8.14
cc_280 N_A_847_1221#_c_328_n N_VGND_c_666_n 0.0648349f $X=4.375 $Y=6.25 $X2=0
+ $Y2=0
cc_281 N_A_847_1221#_c_330_n N_VGND_c_666_n 0.0425081f $X=5.77 $Y=5.83 $X2=0
+ $Y2=0
cc_282 N_A_847_1221#_c_334_n N_VGND_c_666_n 0.0648349f $X=5.935 $Y=6.25 $X2=0
+ $Y2=0
cc_283 N_A_847_1221#_c_334_n N_VGND_c_641_n 0.0648349f $X=5.935 $Y=6.25 $X2=0
+ $Y2=0
cc_284 N_A_847_1221#_c_313_n N_VGND_c_641_n 0.0476157f $X=7.6 $Y=5.83 $X2=0
+ $Y2=0
cc_285 N_A_847_1221#_c_328_n N_VGND_c_647_n 0.0240827f $X=4.375 $Y=6.25 $X2=0
+ $Y2=0
cc_286 N_A_847_1221#_c_334_n N_VGND_c_647_n 0.0240827f $X=5.935 $Y=6.25 $X2=0
+ $Y2=0
cc_287 N_A_935_141#_c_373_n N_A_1353_107#_c_494_n 0.0401197f $X=6.515 $Y=2.145
+ $X2=0.24 $Y2=8.14
cc_288 N_A_935_141#_c_374_n N_A_1353_107#_c_494_n 0.0401197f $X=7.295 $Y=2.145
+ $X2=0.24 $Y2=8.14
cc_289 N_A_935_141#_c_376_n N_A_1353_107#_c_474_n 0.084984f $X=8.855 $Y=2.145
+ $X2=0 $Y2=0
cc_290 N_A_935_141#_c_376_n N_A_1353_107#_c_454_n 0.0199658f $X=8.855 $Y=2.145
+ $X2=10.32 $Y2=8.14
cc_291 N_A_935_141#_c_394_n N_A_1353_107#_c_454_n 0.0277655f $X=6.405 $Y=2.31
+ $X2=10.32 $Y2=8.14
cc_292 N_A_935_141#_c_376_n N_A_1353_107#_c_466_n 0.00949295f $X=8.855 $Y=2.145
+ $X2=0 $Y2=0
cc_293 N_A_935_141#_c_375_n N_A_1353_107#_c_500_n 0.0401197f $X=8.075 $Y=2.145
+ $X2=4.8 $Y2=0
cc_294 N_A_935_141#_c_376_n N_A_1353_107#_c_500_n 0.0401197f $X=8.855 $Y=2.145
+ $X2=4.8 $Y2=0
cc_295 N_A_935_141#_c_376_n N_A_1353_107#_c_470_n 0.039042f $X=8.855 $Y=2.145
+ $X2=0 $Y2=0
cc_296 N_A_935_141#_c_376_n N_VPWR_c_547_n 0.00591526f $X=8.855 $Y=2.145
+ $X2=10.32 $Y2=0
cc_297 N_A_935_141#_c_386_n N_VPWR_c_538_n 0.0010968f $X=4.815 $Y=2.49 $X2=0
+ $Y2=0
cc_298 N_A_935_141#_c_377_n N_VGND_c_622_n 0.0147545f $X=4.815 $Y=0.85 $X2=0
+ $Y2=0
cc_299 N_A_935_141#_c_373_n N_VGND_c_628_n 0.0146836f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_300 N_A_935_141#_c_374_n N_VGND_c_628_n 0.0146836f $X=7.295 $Y=2.145 $X2=0
+ $Y2=0
cc_301 N_A_935_141#_c_375_n N_VGND_c_630_n 0.0146836f $X=8.075 $Y=2.145 $X2=0
+ $Y2=0
cc_302 N_A_935_141#_c_376_n N_VGND_c_630_n 0.0181045f $X=8.855 $Y=2.145 $X2=0
+ $Y2=0
cc_303 N_A_935_141#_c_373_n N_VGND_c_634_n 0.00348095f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_304 N_A_935_141#_c_374_n N_VGND_c_636_n 0.00322203f $X=7.295 $Y=2.145
+ $X2=5.28 $Y2=0
cc_305 N_A_935_141#_c_375_n N_VGND_c_636_n 0.00322203f $X=8.075 $Y=2.145
+ $X2=5.28 $Y2=0
cc_306 N_A_935_141#_c_377_n N_VGND_c_639_n 0.0217496f $X=4.815 $Y=0.85 $X2=0
+ $Y2=0
cc_307 N_A_935_141#_c_379_n N_VGND_c_639_n 0.0165367f $X=4.98 $Y=1.31 $X2=0
+ $Y2=0
cc_308 N_A_935_141#_c_373_n N_VGND_c_640_n 0.0582646f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_309 N_A_935_141#_c_374_n N_VGND_c_640_n 0.00129485f $X=7.295 $Y=2.145 $X2=0
+ $Y2=0
cc_310 N_A_935_141#_c_378_n N_VGND_c_640_n 0.0304579f $X=5.33 $Y=1.31 $X2=0
+ $Y2=0
cc_311 N_A_935_141#_c_381_n N_VGND_c_640_n 0.0435029f $X=5.495 $Y=2.145 $X2=0
+ $Y2=0
cc_312 N_A_935_141#_c_394_n N_VGND_c_640_n 0.0457912f $X=6.405 $Y=2.31 $X2=0
+ $Y2=0
cc_313 N_A_935_141#_c_383_n N_VGND_c_640_n 0.00991638f $X=6.265 $Y=2.31 $X2=0
+ $Y2=0
cc_314 N_A_935_141#_c_373_n N_VGND_c_705_n 0.00129485f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_315 N_A_935_141#_c_374_n N_VGND_c_705_n 0.0567946f $X=7.295 $Y=2.145 $X2=0
+ $Y2=0
cc_316 N_A_935_141#_c_375_n N_VGND_c_705_n 0.0567946f $X=8.075 $Y=2.145 $X2=0
+ $Y2=0
cc_317 N_A_935_141#_c_376_n N_VGND_c_705_n 0.00362441f $X=8.855 $Y=2.145 $X2=0
+ $Y2=0
cc_318 N_A_935_141#_c_375_n N_VGND_c_642_n 0.00129485f $X=8.075 $Y=2.145 $X2=0
+ $Y2=0
cc_319 N_A_935_141#_c_376_n N_VGND_c_642_n 0.0635146f $X=8.855 $Y=2.145 $X2=0
+ $Y2=0
cc_320 N_A_935_141#_c_373_n N_VGND_c_643_n 0.0157032f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_321 N_A_935_141#_c_374_n N_VGND_c_643_n 0.0157032f $X=7.295 $Y=2.145 $X2=0
+ $Y2=0
cc_322 N_A_935_141#_c_375_n N_VGND_c_643_n 0.0157032f $X=8.075 $Y=2.145 $X2=0
+ $Y2=0
cc_323 N_A_935_141#_c_376_n N_VGND_c_643_n 0.0157032f $X=8.855 $Y=2.145 $X2=0
+ $Y2=0
cc_324 N_A_935_141#_c_377_n N_VGND_c_643_n 0.0120786f $X=4.815 $Y=0.85 $X2=0
+ $Y2=0
cc_325 N_A_935_141#_c_378_n N_VGND_c_643_n 0.0268634f $X=5.33 $Y=1.31 $X2=0
+ $Y2=0
cc_326 N_A_1353_107#_M1001_g N_VPWR_c_540_n 0.0131793f $X=9.895 $Y=5.175 $X2=0
+ $Y2=0
cc_327 N_A_1353_107#_c_450_n N_VPWR_c_543_n 0.0135895f $X=9.645 $Y=6.39
+ $X2=-0.33 $Y2=-0.265
cc_328 N_A_1353_107#_M1001_g N_VPWR_c_543_n 0.048726f $X=9.895 $Y=5.175
+ $X2=-0.33 $Y2=-0.265
cc_329 N_A_1353_107#_c_461_n N_VPWR_c_543_n 0.00629978f $X=8.8 $Y=4.635
+ $X2=-0.33 $Y2=-0.265
cc_330 N_A_1353_107#_c_467_n N_VPWR_c_543_n 0.0126425f $X=8.38 $Y=5.205
+ $X2=-0.33 $Y2=-0.265
cc_331 N_A_1353_107#_c_455_n N_VPWR_c_543_n 0.0259241f $X=8.8 $Y=6.39 $X2=-0.33
+ $Y2=-0.265
cc_332 N_A_1353_107#_c_471_n N_VPWR_c_543_n 0.021884f $X=8.8 $Y=5.37 $X2=-0.33
+ $Y2=-0.265
cc_333 N_A_1353_107#_c_472_n N_VPWR_c_543_n 0.00612879f $X=8.8 $Y=5.37 $X2=-0.33
+ $Y2=-0.265
cc_334 N_A_1353_107#_c_461_n N_VPWR_c_544_n 0.0170233f $X=8.8 $Y=4.635 $X2=0.24
+ $Y2=0
cc_335 N_A_1353_107#_c_467_n N_VPWR_c_544_n 0.0188122f $X=8.38 $Y=5.205 $X2=0.24
+ $Y2=0
cc_336 N_A_1353_107#_c_471_n N_VPWR_c_544_n 0.00554595f $X=8.8 $Y=5.37 $X2=0.24
+ $Y2=0
cc_337 N_A_1353_107#_c_466_n N_VPWR_c_547_n 0.0119353f $X=8.38 $Y=3.125
+ $X2=10.32 $Y2=0
cc_338 N_A_1353_107#_c_467_n N_VPWR_c_547_n 0.0184731f $X=8.38 $Y=5.205
+ $X2=10.32 $Y2=0
cc_339 N_A_1353_107#_M1003_s N_VPWR_c_538_n 0.00118086f $X=7.6 $Y=2.815 $X2=0
+ $Y2=0
cc_340 N_A_1353_107#_c_466_n N_VPWR_c_538_n 0.00486511f $X=8.38 $Y=3.125 $X2=0
+ $Y2=0
cc_341 N_A_1353_107#_c_467_n N_VPWR_c_538_n 0.0374126f $X=8.38 $Y=5.205 $X2=0
+ $Y2=0
cc_342 N_A_1353_107#_M1001_g N_VPWR_c_539_n 0.0196379f $X=9.895 $Y=5.175 $X2=0
+ $Y2=0
cc_343 N_A_1353_107#_c_461_n N_VPWR_c_539_n 0.0202019f $X=8.8 $Y=4.635 $X2=0
+ $Y2=0
cc_344 N_A_1353_107#_c_467_n N_VPWR_c_539_n 0.0357766f $X=8.38 $Y=5.205 $X2=0
+ $Y2=0
cc_345 N_A_1353_107#_c_471_n N_VPWR_c_539_n 0.00959858f $X=8.8 $Y=5.37 $X2=0
+ $Y2=0
cc_346 N_A_1353_107#_M1001_g N_X_c_605_n 0.0525051f $X=9.895 $Y=5.175 $X2=0
+ $Y2=0
cc_347 N_A_1353_107#_M1004_g N_X_c_605_n 0.0378537f $X=9.895 $Y=7.23 $X2=0 $Y2=0
cc_348 N_A_1353_107#_c_453_n N_X_c_605_n 0.0231667f $X=9.895 $Y=6.39 $X2=0 $Y2=0
cc_349 N_A_1353_107#_c_494_n N_VGND_c_628_n 0.0211458f $X=6.905 $Y=0.68 $X2=0
+ $Y2=0
cc_350 N_A_1353_107#_c_500_n N_VGND_c_630_n 0.0211458f $X=8.465 $Y=0.68 $X2=0
+ $Y2=0
cc_351 N_A_1353_107#_c_494_n N_VGND_c_640_n 0.0648349f $X=6.905 $Y=0.68 $X2=0
+ $Y2=0
cc_352 N_A_1353_107#_c_494_n N_VGND_c_705_n 0.0648349f $X=6.905 $Y=0.68 $X2=0
+ $Y2=0
cc_353 N_A_1353_107#_c_474_n N_VGND_c_705_n 0.0425081f $X=8.215 $Y=2.31 $X2=0
+ $Y2=0
cc_354 N_A_1353_107#_c_500_n N_VGND_c_705_n 0.0648349f $X=8.465 $Y=0.68 $X2=0
+ $Y2=0
cc_355 N_A_1353_107#_c_500_n N_VGND_c_642_n 0.0648349f $X=8.465 $Y=0.68 $X2=0
+ $Y2=0
cc_356 N_A_1353_107#_c_494_n N_VGND_c_643_n 0.0240827f $X=6.905 $Y=0.68 $X2=0
+ $Y2=0
cc_357 N_A_1353_107#_c_500_n N_VGND_c_643_n 0.0240827f $X=8.465 $Y=0.68 $X2=0
+ $Y2=0
cc_358 N_A_1353_107#_c_450_n N_VGND_c_645_n 0.017439f $X=9.645 $Y=6.39 $X2=0
+ $Y2=0
cc_359 N_A_1353_107#_M1004_g N_VGND_c_645_n 0.0456555f $X=9.895 $Y=7.23 $X2=0
+ $Y2=0
cc_360 N_A_1353_107#_M1004_g N_VGND_c_647_n 0.0208706f $X=9.895 $Y=7.23 $X2=0
+ $Y2=0
cc_361 N_VPWR_c_540_n N_X_c_605_n 0.0141539f $X=9.505 $Y=4.8 $X2=0 $Y2=0
cc_362 N_VPWR_c_543_n N_X_c_605_n 0.0541691f $X=9.505 $Y=4.97 $X2=0 $Y2=0
cc_363 N_VPWR_c_539_n N_X_c_605_n 0.0434173f $X=9.685 $Y=4.58 $X2=0 $Y2=0
cc_364 N_X_c_605_n N_VGND_c_645_n 0.0356255f $X=10.285 $Y=4.57 $X2=0 $Y2=0
cc_365 N_X_c_605_n N_VGND_c_647_n 0.0326456f $X=10.285 $Y=4.57 $X2=0 $Y2=0
