* NGSPICE file created from sky130_fd_sc_hvl__dfstp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
M1000 VPWR a_1000_81# a_982_529# VPB phv w=420000u l=500000u
+  ad=1.5397e+12p pd=1.406e+07u as=8.82e+10p ps=1.26e+06u
M1001 Q a_2553_203# VPWR VPB phv w=1e+06u l=500000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1002 a_642_107# D VPWR VPB phv w=420000u l=500000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1003 VGND a_1000_81# a_958_107# VNB nhv w=420000u l=500000u
+  ad=9.711e+11p pd=1.012e+07u as=8.82e+10p ps=1.26e+06u
M1004 VGND a_1787_137# a_2553_203# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1005 VPWR a_1787_137# a_2553_203# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u
M1006 a_798_107# a_30_131# a_642_107# VNB nhv w=420000u l=500000u
+  ad=1.26e+11p pd=1.44e+06u as=1.176e+11p ps=1.4e+06u
M1007 a_2031_177# a_1787_137# VGND VNB nhv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1008 Q a_2553_203# VGND VNB nhv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
M1009 a_1000_81# a_798_107# VPWR VPB phv w=420000u l=500000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1010 a_1787_137# SET_B VPWR VPB phv w=420000u l=500000u
+  ad=5.2205e+11p pd=4.35e+06u as=0p ps=0u
M1011 a_1653_515# a_798_107# VPWR VPB phv w=1e+06u l=500000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1012 VPWR a_1787_137# a_2031_177# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=1.848e+11p ps=1.72e+06u
M1013 a_1645_137# a_798_107# VGND VNB nhv w=750000u l=500000u
+  ad=1.575e+11p pd=1.92e+06u as=0p ps=0u
M1014 a_1787_137# a_30_131# a_1653_515# VPB phv w=1e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1787_137# a_340_593# a_1645_137# VNB nhv w=750000u l=500000u
+  ad=2.967e+11p pd=2.52e+06u as=0p ps=0u
M1016 VPWR CLK a_30_131# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u
M1017 VGND CLK a_30_131# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1018 a_1989_203# a_30_131# a_1787_137# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1019 a_2131_203# a_2031_177# a_1989_203# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1020 VGND SET_B a_2131_203# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_982_529# a_30_131# a_798_107# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1022 VGND SET_B a_1268_251# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=2.838e+11p ps=2.34e+06u
M1023 a_958_107# a_340_593# a_798_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_798_107# a_340_593# a_642_107# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1268_251# a_798_107# a_1000_81# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1026 VPWR SET_B a_1000_81# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_642_107# D VGND VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_340_593# a_30_131# VPWR VPB phv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
M1029 a_340_593# a_30_131# VGND VNB nhv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1030 a_1989_515# a_340_593# a_1787_137# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1031 VPWR a_2031_177# a_1989_515# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends

