* File: sky130_fd_sc_hvl__sdfxbp_1.pxi.spice
* Created: Wed Sep  2 09:10:25 2020
* 
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%VNB N_VNB_M1028_b VNB N_VNB_c_2_p
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%VNB
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%VPB N_VPB_M1022_b VPB N_VPB_c_124_p
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%VPB
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%SCE N_SCE_M1022_g N_SCE_M1028_g N_SCE_M1020_g
+ N_SCE_M1018_g SCE SCE SCE SCE SCE N_SCE_c_301_n N_SCE_c_309_n N_SCE_c_314_p
+ N_SCE_c_302_n N_SCE_c_321_p N_SCE_c_334_p PM_SKY130_FD_SC_HVL__SDFXBP_1%SCE
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%SCD SCD N_SCD_M1019_g N_SCD_c_374_n
+ N_SCD_M1000_g PM_SKY130_FD_SC_HVL__SDFXBP_1%SCD
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_30_515# N_A_30_515#_M1028_s
+ N_A_30_515#_M1022_s N_A_30_515#_M1013_g N_A_30_515#_c_399_n
+ N_A_30_515#_M1016_g N_A_30_515#_c_411_n N_A_30_515#_c_400_n
+ N_A_30_515#_c_401_n N_A_30_515#_c_402_n N_A_30_515#_c_404_n
+ N_A_30_515#_c_412_n N_A_30_515#_c_405_n N_A_30_515#_c_431_n
+ N_A_30_515#_c_433_n N_A_30_515#_c_406_n
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%A_30_515#
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%D N_D_M1014_g N_D_M1007_g D D D N_D_c_486_n
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%D
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1124_81# N_A_1124_81#_M1017_d
+ N_A_1124_81#_M1002_d N_A_1124_81#_c_526_n N_A_1124_81#_M1003_g
+ N_A_1124_81#_c_528_n N_A_1124_81#_M1035_g N_A_1124_81#_c_534_n
+ N_A_1124_81#_c_535_n N_A_1124_81#_c_536_n N_A_1124_81#_c_537_n
+ N_A_1124_81#_c_538_n N_A_1124_81#_c_529_n N_A_1124_81#_c_540_n
+ N_A_1124_81#_c_530_n PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1124_81#
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1067_107# N_A_1067_107#_M1003_s
+ N_A_1067_107#_M1005_s N_A_1067_107#_M1035_s N_A_1067_107#_M1025_d
+ N_A_1067_107#_c_618_n N_A_1067_107#_M1012_g N_A_1067_107#_M1001_g
+ N_A_1067_107#_c_619_n N_A_1067_107#_c_620_n N_A_1067_107#_c_621_n
+ N_A_1067_107#_c_630_n N_A_1067_107#_c_631_n N_A_1067_107#_c_622_n
+ N_A_1067_107#_c_623_n N_A_1067_107#_c_632_n N_A_1067_107#_c_633_n
+ N_A_1067_107#_c_634_n N_A_1067_107#_c_624_n N_A_1067_107#_c_625_n
+ N_A_1067_107#_c_637_n PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1067_107#
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1570_457# N_A_1570_457#_M1026_d
+ N_A_1570_457#_M1008_d N_A_1570_457#_M1002_g N_A_1570_457#_M1017_g
+ N_A_1570_457#_c_781_n N_A_1570_457#_M1004_g N_A_1570_457#_c_796_n
+ N_A_1570_457#_M1025_g N_A_1570_457#_c_783_n N_A_1570_457#_M1029_g
+ N_A_1570_457#_c_784_n N_A_1570_457#_c_785_n N_A_1570_457#_c_798_n
+ N_A_1570_457#_c_799_n N_A_1570_457#_c_800_n N_A_1570_457#_c_882_p
+ N_A_1570_457#_c_878_p N_A_1570_457#_c_801_n N_A_1570_457#_c_786_n
+ N_A_1570_457#_c_802_n N_A_1570_457#_c_787_n N_A_1570_457#_c_788_n
+ N_A_1570_457#_c_790_n N_A_1570_457#_c_792_n N_A_1570_457#_c_820_n
+ N_A_1570_457#_c_793_n N_A_1570_457#_c_875_p N_A_1570_457#_c_881_p
+ N_A_1570_457#_c_794_n N_A_1570_457#_c_868_p N_A_1570_457#_c_795_n
+ N_A_1570_457#_c_913_p N_A_1570_457#_M1024_g N_A_1570_457#_c_805_n
+ N_A_1570_457#_c_806_n PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1570_457#
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1726_453# N_A_1726_453#_M1004_s
+ N_A_1726_453#_M1024_s N_A_1726_453#_M1027_g N_A_1726_453#_M1034_g
+ N_A_1726_453#_c_968_n N_A_1726_453#_M1005_g N_A_1726_453#_c_980_n
+ N_A_1726_453#_c_969_n N_A_1726_453#_c_970_n N_A_1726_453#_c_972_n
+ N_A_1726_453#_c_973_n N_A_1726_453#_c_987_n N_A_1726_453#_c_981_n
+ N_A_1726_453#_c_974_n N_A_1726_453#_c_999_n N_A_1726_453#_M1030_g
+ N_A_1726_453#_c_976_n PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1726_453#
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%CLK N_CLK_c_1076_n N_CLK_M1008_g N_CLK_c_1073_n
+ N_CLK_M1026_g CLK CLK PM_SKY130_FD_SC_HVL__SDFXBP_1%CLK
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_2789_147# N_A_2789_147#_M1006_d
+ N_A_2789_147#_M1015_d N_A_2789_147#_M1031_g N_A_2789_147#_c_1122_n
+ N_A_2789_147#_M1023_g N_A_2789_147#_M1010_g N_A_2789_147#_M1009_g
+ N_A_2789_147#_M1032_g N_A_2789_147#_M1033_g N_A_2789_147#_c_1127_n
+ N_A_2789_147#_c_1128_n N_A_2789_147#_c_1118_n N_A_2789_147#_c_1130_n
+ N_A_2789_147#_c_1131_n N_A_2789_147#_c_1134_n N_A_2789_147#_c_1185_p
+ N_A_2789_147#_c_1137_n N_A_2789_147#_c_1138_n N_A_2789_147#_c_1139_n
+ N_A_2789_147#_c_1174_p N_A_2789_147#_c_1120_n
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%A_2789_147#
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_2518_445# N_A_2518_445#_M1005_d
+ N_A_2518_445#_M1034_d N_A_2518_445#_c_1223_n N_A_2518_445#_M1006_g
+ N_A_2518_445#_M1015_g N_A_2518_445#_c_1231_n N_A_2518_445#_c_1232_n
+ N_A_2518_445#_c_1225_n N_A_2518_445#_c_1234_n N_A_2518_445#_c_1235_n
+ N_A_2518_445#_c_1226_n N_A_2518_445#_c_1227_n
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%A_2518_445#
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_3531_107# N_A_3531_107#_M1032_d
+ N_A_3531_107#_M1033_d N_A_3531_107#_M1011_g N_A_3531_107#_M1021_g
+ N_A_3531_107#_c_1305_n N_A_3531_107#_c_1313_n N_A_3531_107#_c_1307_n
+ N_A_3531_107#_c_1308_n N_A_3531_107#_c_1309_n N_A_3531_107#_c_1317_n
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%A_3531_107#
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%VPWR N_VPWR_M1022_d N_VPWR_M1000_d
+ N_VPWR_M1035_d N_VPWR_M1024_d N_VPWR_M1023_d N_VPWR_M1009_d N_VPWR_M1021_s
+ VPWR N_VPWR_c_1343_n N_VPWR_c_1346_n N_VPWR_c_1349_n N_VPWR_c_1352_n
+ N_VPWR_c_1355_n N_VPWR_c_1358_n N_VPWR_c_1361_n N_VPWR_c_1364_n
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%VPWR
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_268_659# N_A_268_659#_M1000_s
+ N_A_268_659#_M1016_s N_A_268_659#_c_1472_n N_A_268_659#_c_1475_n
+ N_A_268_659#_c_1476_n N_A_268_659#_c_1477_n
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%A_268_659#
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_581_659# N_A_581_659#_M1018_d
+ N_A_581_659#_M1007_d N_A_581_659#_c_1504_n N_A_581_659#_c_1505_n
+ N_A_581_659#_c_1508_n N_A_581_659#_c_1511_n N_A_581_659#_c_1512_n
+ N_A_581_659#_c_1521_n N_A_581_659#_c_1513_n
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%A_581_659#
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_567_107# N_A_567_107#_M1020_d
+ N_A_567_107#_M1017_s N_A_567_107#_M1016_d N_A_567_107#_M1027_d
+ N_A_567_107#_c_1550_n N_A_567_107#_c_1551_n N_A_567_107#_c_1563_n
+ N_A_567_107#_c_1584_n N_A_567_107#_c_1564_n N_A_567_107#_c_1565_n
+ N_A_567_107#_c_1568_n N_A_567_107#_c_1552_n N_A_567_107#_c_1553_n
+ N_A_567_107#_c_1555_n N_A_567_107#_c_1618_n N_A_567_107#_c_1619_n
+ N_A_567_107#_c_1621_n N_A_567_107#_c_1557_n N_A_567_107#_c_1624_n
+ N_A_567_107#_c_1572_n N_A_567_107#_c_1628_n N_A_567_107#_c_1629_n
+ N_A_567_107#_c_1664_n N_A_567_107#_c_1558_n N_A_567_107#_c_1573_n
+ N_A_567_107#_c_1559_n N_A_567_107#_c_1634_n N_A_567_107#_c_1673_n
+ N_A_567_107#_c_1576_n N_A_567_107#_c_1561_n N_A_567_107#_c_1579_n
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%A_567_107#
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_2365_445# N_A_2365_445#_M1034_s
+ N_A_2365_445#_M1023_s N_A_2365_445#_c_1742_n N_A_2365_445#_c_1743_n
+ N_A_2365_445#_c_1746_n N_A_2365_445#_c_1749_n
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%A_2365_445#
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%Q N_Q_M1010_s N_Q_M1009_s N_Q_c_1783_n Q Q Q Q
+ N_Q_c_1781_n N_Q_c_1785_n PM_SKY130_FD_SC_HVL__SDFXBP_1%Q
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%Q_N N_Q_N_M1011_d N_Q_N_M1021_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_1809_n PM_SKY130_FD_SC_HVL__SDFXBP_1%Q_N
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%VGND N_VGND_M1028_d N_VGND_M1014_d
+ N_VGND_M1003_d N_VGND_M1004_d N_VGND_M1031_d N_VGND_M1010_d N_VGND_M1011_s
+ VGND N_VGND_c_1822_n N_VGND_c_1824_n N_VGND_c_1826_n N_VGND_c_1828_n
+ N_VGND_c_1830_n N_VGND_c_1832_n N_VGND_c_1834_n N_VGND_c_1836_n
+ PM_SKY130_FD_SC_HVL__SDFXBP_1%VGND
x_PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1454_173# N_A_1454_173#_M1012_d
+ N_A_1454_173#_M1030_d N_A_1454_173#_c_1935_n N_A_1454_173#_c_1937_n
+ N_A_1454_173#_c_1938_n PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1454_173#
cc_1 N_VNB_M1028_b N_SCE_M1028_g 0.0469269f $X=-0.33 $Y=-0.265 $X2=1.095
+ $Y2=0.745
cc_2 N_VNB_c_2_p N_SCE_M1028_g 9.58849e-19 $X=0.24 $Y=0 $X2=1.095 $Y2=0.745
cc_3 N_VNB_M1028_b N_SCE_M1020_g 0.115674f $X=-0.33 $Y=-0.265 $X2=2.585
+ $Y2=0.745
cc_4 N_VNB_c_2_p N_SCE_M1020_g 0.0023273f $X=0.24 $Y=0 $X2=2.585 $Y2=0.745
cc_5 N_VNB_M1028_b N_SCE_c_301_n 0.13009f $X=-0.33 $Y=-0.265 $X2=0.73 $Y2=1.715
cc_6 N_VNB_M1028_b N_SCE_c_302_n 0.0204781f $X=-0.33 $Y=-0.265 $X2=2.425
+ $Y2=1.65
cc_7 N_VNB_M1028_b N_SCD_M1019_g 0.108056f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_8 N_VNB_c_2_p N_SCD_M1019_g 5.86481e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_9 N_VNB_M1028_b N_A_30_515#_M1013_g 0.0487528f $X=-0.33 $Y=-0.265 $X2=2.585
+ $Y2=2.075
cc_10 N_VNB_c_2_p N_A_30_515#_M1013_g 0.0023273f $X=0.24 $Y=0 $X2=2.585
+ $Y2=2.075
cc_11 N_VNB_M1028_b N_A_30_515#_c_399_n 0.00192584f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1028_b N_A_30_515#_c_400_n 0.00682097f $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=1.75
cc_13 N_VNB_M1028_b N_A_30_515#_c_401_n 0.0110419f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_M1028_b N_A_30_515#_c_402_n 0.030504f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_15 N_VNB_c_2_p N_A_30_515#_c_402_n 8.20017e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_16 N_VNB_M1028_b N_A_30_515#_c_404_n 0.0198038f $X=-0.33 $Y=-0.265 $X2=0.88
+ $Y2=1.715
cc_17 N_VNB_M1028_b N_A_30_515#_c_405_n 0.0258345f $X=-0.33 $Y=-0.265 $X2=2.59
+ $Y2=2.26
cc_18 N_VNB_M1028_b N_A_30_515#_c_406_n 0.0728198f $X=-0.33 $Y=-0.265 $X2=0.895
+ $Y2=1.65
cc_19 N_VNB_M1028_b N_D_M1014_g 0.0427468f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=2.785
cc_20 N_VNB_M1028_b N_D_M1007_g 0.00197426f $X=-0.33 $Y=-0.265 $X2=1.095
+ $Y2=0.745
cc_21 N_VNB_M1028_b D 2.22386e-19 $X=-0.33 $Y=-0.265 $X2=2.585 $Y2=2.075
cc_22 N_VNB_M1028_b N_D_c_486_n 0.168248f $X=-0.33 $Y=-0.265 $X2=2.075 $Y2=1.58
cc_23 N_VNB_M1028_b N_A_1124_81#_c_526_n 0.0456338f $X=-0.33 $Y=-0.265 $X2=1.095
+ $Y2=0.745
cc_24 N_VNB_c_2_p N_A_1124_81#_c_526_n 5.98017e-19 $X=0.24 $Y=0 $X2=1.095
+ $Y2=0.745
cc_25 N_VNB_M1028_b N_A_1124_81#_c_528_n 0.0660218f $X=-0.33 $Y=-0.265 $X2=2.585
+ $Y2=0.745
cc_26 N_VNB_M1028_b N_A_1124_81#_c_529_n 0.00411421f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_27 N_VNB_M1028_b N_A_1124_81#_c_530_n 0.00518499f $X=-0.33 $Y=-0.265 $X2=0.88
+ $Y2=1.085
cc_28 N_VNB_M1028_b N_A_1067_107#_c_618_n 0.0451202f $X=-0.33 $Y=-0.265
+ $X2=2.655 $Y2=2.785
cc_29 N_VNB_M1028_b N_A_1067_107#_c_619_n 0.00983132f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_30 N_VNB_M1028_b N_A_1067_107#_c_620_n 0.00748349f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_31 N_VNB_M1028_b N_A_1067_107#_c_621_n 0.00377889f $X=-0.33 $Y=-0.265
+ $X2=0.73 $Y2=1.715
cc_32 N_VNB_M1028_b N_A_1067_107#_c_622_n 0.00619908f $X=-0.33 $Y=-0.265
+ $X2=2.62 $Y2=2.26
cc_33 N_VNB_M1028_b N_A_1067_107#_c_623_n 0.00672881f $X=-0.33 $Y=-0.265
+ $X2=2.59 $Y2=2.26
cc_34 N_VNB_M1028_b N_A_1067_107#_c_624_n 0.0766236f $X=-0.33 $Y=-0.265 $X2=2.59
+ $Y2=2.26
cc_35 N_VNB_M1028_b N_A_1067_107#_c_625_n 9.7518e-19 $X=-0.33 $Y=-0.265 $X2=0.73
+ $Y2=1.65
cc_36 N_VNB_M1028_b N_A_1570_457#_c_781_n 0.0452033f $X=-0.33 $Y=-0.265
+ $X2=2.655 $Y2=3.505
cc_37 N_VNB_c_2_p N_A_1570_457#_c_781_n 9.58849e-19 $X=0.24 $Y=0 $X2=2.655
+ $Y2=3.505
cc_38 N_VNB_M1028_b N_A_1570_457#_c_783_n 0.0387121f $X=-0.33 $Y=-0.265
+ $X2=2.555 $Y2=1.58
cc_39 N_VNB_M1028_b N_A_1570_457#_c_784_n 0.0361314f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_M1028_b N_A_1570_457#_c_785_n 0.0553757f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_41 N_VNB_M1028_b N_A_1570_457#_c_786_n 0.00997126f $X=-0.33 $Y=-0.265
+ $X2=2.425 $Y2=1.65
cc_42 N_VNB_M1028_b N_A_1570_457#_c_787_n 0.00904945f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_M1028_b N_A_1570_457#_c_788_n 0.0937348f $X=-0.33 $Y=-0.265 $X2=0.73
+ $Y2=1.985
cc_44 N_VNB_c_2_p N_A_1570_457#_c_788_n 0.00427487f $X=0.24 $Y=0 $X2=0.73
+ $Y2=1.985
cc_45 N_VNB_M1028_b N_A_1570_457#_c_790_n 0.0100057f $X=-0.33 $Y=-0.265 $X2=0.73
+ $Y2=1.75
cc_46 N_VNB_c_2_p N_A_1570_457#_c_790_n 6.02919e-19 $X=0.24 $Y=0 $X2=0.73
+ $Y2=1.75
cc_47 N_VNB_M1028_b N_A_1570_457#_c_792_n 0.00408115f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_M1028_b N_A_1570_457#_c_793_n 0.0338484f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_49 N_VNB_M1028_b N_A_1570_457#_c_794_n 0.0840011f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_M1028_b N_A_1570_457#_c_795_n 0.0568554f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_51 N_VNB_M1028_b N_A_1726_453#_c_968_n 0.0362216f $X=-0.33 $Y=-0.265
+ $X2=2.655 $Y2=3.505
cc_52 N_VNB_M1028_b N_A_1726_453#_c_969_n 0.0115825f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_53 N_VNB_M1028_b N_A_1726_453#_c_970_n 0.0171918f $X=-0.33 $Y=-0.265 $X2=0.73
+ $Y2=1.715
cc_54 N_VNB_c_2_p N_A_1726_453#_c_970_n 8.20017e-19 $X=0.24 $Y=0 $X2=0.73
+ $Y2=1.715
cc_55 N_VNB_M1028_b N_A_1726_453#_c_972_n 0.0214005f $X=-0.33 $Y=-0.265 $X2=0.88
+ $Y2=2.24
cc_56 N_VNB_M1028_b N_A_1726_453#_c_973_n 0.0124342f $X=-0.33 $Y=-0.265 $X2=2.62
+ $Y2=2.26
cc_57 N_VNB_M1028_b N_A_1726_453#_c_974_n 0.00383736f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_58 N_VNB_M1028_b N_A_1726_453#_M1030_g 0.0816993f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_59 N_VNB_M1028_b N_A_1726_453#_c_976_n 0.108013f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_60 N_VNB_M1028_b N_CLK_c_1073_n 0.023028f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_61 N_VNB_M1028_b N_CLK_M1026_g 0.109555f $X=-0.33 $Y=-0.265 $X2=1.095
+ $Y2=0.745
cc_62 N_VNB_c_2_p N_CLK_M1026_g 5.86481e-19 $X=0.24 $Y=0 $X2=1.095 $Y2=0.745
cc_63 N_VNB_M1028_b N_A_2789_147#_M1031_g 0.080714f $X=-0.33 $Y=-0.265 $X2=2.585
+ $Y2=2.075
cc_64 N_VNB_M1028_b N_A_2789_147#_M1010_g 0.0476678f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_65 N_VNB_c_2_p N_A_2789_147#_M1010_g 9.58849e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_66 N_VNB_M1028_b N_A_2789_147#_M1032_g 0.0813165f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_67 N_VNB_c_2_p N_A_2789_147#_M1032_g 0.00112176f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_68 N_VNB_M1028_b N_A_2789_147#_c_1118_n 0.0296777f $X=-0.33 $Y=-0.265
+ $X2=2.62 $Y2=2.075
cc_69 N_VNB_c_2_p N_A_2789_147#_c_1118_n 0.00112468f $X=0.24 $Y=0 $X2=2.62
+ $Y2=2.075
cc_70 N_VNB_M1028_b N_A_2789_147#_c_1120_n 0.0792325f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_71 N_VNB_M1028_b N_A_2518_445#_c_1223_n 0.0537103f $X=-0.33 $Y=-0.265
+ $X2=1.095 $Y2=0.745
cc_72 N_VNB_c_2_p N_A_2518_445#_c_1223_n 0.00221559f $X=0.24 $Y=0 $X2=1.095
+ $Y2=0.745
cc_73 N_VNB_M1028_b N_A_2518_445#_c_1225_n 0.00641156f $X=-0.33 $Y=-0.265
+ $X2=2.555 $Y2=1.58
cc_74 N_VNB_M1028_b N_A_2518_445#_c_1226_n 0.00473637f $X=-0.33 $Y=-0.265
+ $X2=0.88 $Y2=2.24
cc_75 N_VNB_M1028_b N_A_2518_445#_c_1227_n 0.0799411f $X=-0.33 $Y=-0.265
+ $X2=2.62 $Y2=2.785
cc_76 N_VNB_M1028_b N_A_3531_107#_M1011_g 0.0524616f $X=-0.33 $Y=-0.265
+ $X2=2.585 $Y2=2.075
cc_77 N_VNB_c_2_p N_A_3531_107#_M1011_g 9.58849e-19 $X=0.24 $Y=0 $X2=2.585
+ $Y2=2.075
cc_78 N_VNB_M1028_b N_A_3531_107#_c_1305_n 0.0267782f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=1.58
cc_79 N_VNB_c_2_p N_A_3531_107#_c_1305_n 8.20017e-19 $X=0.24 $Y=0 $X2=0.635
+ $Y2=1.58
cc_80 N_VNB_M1028_b N_A_3531_107#_c_1307_n 0.010258f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_81 N_VNB_M1028_b N_A_3531_107#_c_1308_n 0.00954255f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_82 N_VNB_M1028_b N_A_3531_107#_c_1309_n 0.0583476f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_83 N_VNB_M1028_b N_A_567_107#_c_1550_n 2.40113e-19 $X=-0.33 $Y=-0.265
+ $X2=2.655 $Y2=2.785
cc_84 N_VNB_M1028_b N_A_567_107#_c_1551_n 0.00793695f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_85 N_VNB_M1028_b N_A_567_107#_c_1552_n 0.0193513f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_86 N_VNB_M1028_b N_A_567_107#_c_1553_n 0.0666198f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_87 N_VNB_c_2_p N_A_567_107#_c_1553_n 0.00289338f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_88 N_VNB_M1028_b N_A_567_107#_c_1555_n 0.014726f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_89 N_VNB_c_2_p N_A_567_107#_c_1555_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_90 N_VNB_M1028_b N_A_567_107#_c_1557_n 0.00383119f $X=-0.33 $Y=-0.265
+ $X2=2.59 $Y2=2.26
cc_91 N_VNB_M1028_b N_A_567_107#_c_1558_n 0.0110676f $X=-0.33 $Y=-0.265 $X2=1.68
+ $Y2=1.65
cc_92 N_VNB_M1028_b N_A_567_107#_c_1559_n 0.0133576f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_93 N_VNB_c_2_p N_A_567_107#_c_1559_n 8.67754e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_94 N_VNB_M1028_b N_A_567_107#_c_1561_n 0.0106637f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_95 N_VNB_M1028_b N_Q_c_1781_n 0.022456f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_96 N_VNB_c_2_p N_Q_c_1781_n 8.20017e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_97 N_VNB_M1028_b N_Q_N_c_1809_n 0.063857f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_98 N_VNB_c_2_p N_Q_N_c_1809_n 8.31735e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_99 N_VNB_M1028_b N_VGND_c_1822_n 0.0496364f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_100 N_VNB_c_2_p N_VGND_c_1822_n 0.00269373f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_101 N_VNB_M1028_b N_VGND_c_1824_n 0.0578866f $X=-0.33 $Y=-0.265 $X2=2.62
+ $Y2=2.26
cc_102 N_VNB_c_2_p N_VGND_c_1824_n 0.00262269f $X=0.24 $Y=0 $X2=2.62 $Y2=2.26
cc_103 N_VNB_M1028_b N_VGND_c_1826_n 0.0550114f $X=-0.33 $Y=-0.265 $X2=1.68
+ $Y2=1.65
cc_104 N_VNB_c_2_p N_VGND_c_1826_n 0.0025185f $X=0.24 $Y=0 $X2=1.68 $Y2=1.65
cc_105 N_VNB_M1028_b N_VGND_c_1828_n 0.0468651f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_106 N_VNB_c_2_p N_VGND_c_1828_n 0.00269953f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_107 N_VNB_M1028_b N_VGND_c_1830_n 0.062919f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_108 N_VNB_c_2_p N_VGND_c_1830_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_109 N_VNB_M1028_b N_VGND_c_1832_n 0.0531645f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_110 N_VNB_c_2_p N_VGND_c_1832_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_111 N_VNB_M1028_b N_VGND_c_1834_n 0.0691454f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_112 N_VNB_c_2_p N_VGND_c_1834_n 0.00254859f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_113 N_VNB_M1028_b N_VGND_c_1836_n 0.297766f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_114 N_VNB_c_2_p N_VGND_c_1836_n 2.10493f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_115 N_VNB_M1028_b N_A_1454_173#_c_1935_n 0.0916786f $X=-0.33 $Y=-0.265
+ $X2=1.095 $Y2=0.745
cc_116 N_VNB_c_2_p N_A_1454_173#_c_1935_n 0.00451427f $X=0.24 $Y=0 $X2=1.095
+ $Y2=0.745
cc_117 N_VNB_M1028_b N_A_1454_173#_c_1937_n 0.00916775f $X=-0.33 $Y=-0.265
+ $X2=2.585 $Y2=0.745
cc_118 N_VNB_M1028_b N_A_1454_173#_c_1938_n 0.0167139f $X=-0.33 $Y=-0.265
+ $X2=2.655 $Y2=2.785
cc_119 N_VNB_c_2_p N_A_1454_173#_c_1938_n 6.77859e-19 $X=0.24 $Y=0 $X2=2.655
+ $Y2=2.785
cc_120 N_VPB_M1022_b N_SCE_M1022_g 0.0700931f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=2.785
cc_121 N_VPB_M1022_b N_SCE_M1020_g 0.0169686f $X=-0.33 $Y=1.885 $X2=2.585
+ $Y2=0.745
cc_122 N_VPB_M1022_b N_SCE_M1018_g 0.0782668f $X=-0.33 $Y=1.885 $X2=2.655
+ $Y2=3.505
cc_123 VPB N_SCE_M1018_g 0.00970178f $X=0 $Y=3.955 $X2=2.655 $Y2=3.505
cc_124 N_VPB_c_124_p N_SCE_M1018_g 0.0158633f $X=19.44 $Y=4.07 $X2=2.655
+ $Y2=3.505
cc_125 N_VPB_M1022_b N_SCE_c_301_n 0.0673909f $X=-0.33 $Y=1.885 $X2=0.73
+ $Y2=1.715
cc_126 N_VPB_M1022_b N_SCE_c_309_n 0.0727262f $X=-0.33 $Y=1.885 $X2=2.59
+ $Y2=2.26
cc_127 N_VPB_M1022_b N_SCD_M1019_g 0.160271f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_128 VPB N_SCD_M1019_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_129 N_VPB_c_124_p N_SCD_M1019_g 0.0152133f $X=19.44 $Y=4.07 $X2=0 $Y2=0
cc_130 N_VPB_M1022_b N_SCD_c_374_n 0.00784726f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_131 N_VPB_M1022_b N_A_30_515#_c_399_n 0.0472033f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_132 N_VPB_M1022_b N_A_30_515#_M1016_g 0.0430718f $X=-0.33 $Y=1.885 $X2=2.655
+ $Y2=3.505
cc_133 VPB N_A_30_515#_M1016_g 7.37386e-19 $X=0 $Y=3.955 $X2=2.655 $Y2=3.505
cc_134 N_VPB_c_124_p N_A_30_515#_M1016_g 0.0041461f $X=19.44 $Y=4.07 $X2=2.655
+ $Y2=3.505
cc_135 N_VPB_M1022_b N_A_30_515#_c_411_n 0.106425f $X=-0.33 $Y=1.885 $X2=1.595
+ $Y2=1.58
cc_136 N_VPB_M1022_b N_A_30_515#_c_412_n 0.0283331f $X=-0.33 $Y=1.885 $X2=2.62
+ $Y2=2.26
cc_137 N_VPB_M1022_b N_A_30_515#_c_405_n 0.0323368f $X=-0.33 $Y=1.885 $X2=2.59
+ $Y2=2.26
cc_138 N_VPB_M1022_b N_D_M1007_g 0.144655f $X=-0.33 $Y=1.885 $X2=1.095 $Y2=0.745
cc_139 N_VPB_c_124_p N_D_M1007_g 5.17505e-19 $X=19.44 $Y=4.07 $X2=1.095
+ $Y2=0.745
cc_140 N_VPB_M1022_b D 0.00672348f $X=-0.33 $Y=1.885 $X2=2.585 $Y2=2.075
cc_141 N_VPB_M1022_b N_A_1124_81#_c_528_n 0.17804f $X=-0.33 $Y=1.885 $X2=2.585
+ $Y2=0.745
cc_142 VPB N_A_1124_81#_c_528_n 0.00970178f $X=0 $Y=3.955 $X2=2.585 $Y2=0.745
cc_143 N_VPB_c_124_p N_A_1124_81#_c_528_n 0.0157135f $X=19.44 $Y=4.07 $X2=2.585
+ $Y2=0.745
cc_144 N_VPB_M1022_b N_A_1124_81#_c_534_n 0.016794f $X=-0.33 $Y=1.885 $X2=2.655
+ $Y2=2.785
cc_145 N_VPB_M1022_b N_A_1124_81#_c_535_n 0.00274931f $X=-0.33 $Y=1.885
+ $X2=1.595 $Y2=1.58
cc_146 N_VPB_M1022_b N_A_1124_81#_c_536_n 0.00564869f $X=-0.33 $Y=1.885
+ $X2=2.075 $Y2=1.58
cc_147 N_VPB_M1022_b N_A_1124_81#_c_537_n 4.37313e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_148 N_VPB_M1022_b N_A_1124_81#_c_538_n 0.00239613f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_149 N_VPB_M1022_b N_A_1124_81#_c_529_n 0.00374165f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_150 N_VPB_M1022_b N_A_1124_81#_c_540_n 0.00916587f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_151 N_VPB_M1022_b N_A_1067_107#_M1001_g 0.134202f $X=-0.33 $Y=1.885 $X2=1.115
+ $Y2=1.58
cc_152 VPB N_A_1067_107#_M1001_g 6.77132e-19 $X=0 $Y=3.955 $X2=1.115 $Y2=1.58
cc_153 N_VPB_c_124_p N_A_1067_107#_M1001_g 0.00387149f $X=19.44 $Y=4.07
+ $X2=1.115 $Y2=1.58
cc_154 N_VPB_M1022_b N_A_1067_107#_c_621_n 0.0107004f $X=-0.33 $Y=1.885 $X2=0.73
+ $Y2=1.715
cc_155 N_VPB_M1022_b N_A_1067_107#_c_630_n 0.0125933f $X=-0.33 $Y=1.885 $X2=0.73
+ $Y2=1.715
cc_156 N_VPB_M1022_b N_A_1067_107#_c_631_n 0.00329574f $X=-0.33 $Y=1.885
+ $X2=0.88 $Y2=1.085
cc_157 N_VPB_M1022_b N_A_1067_107#_c_632_n 0.0295859f $X=-0.33 $Y=1.885
+ $X2=0.895 $Y2=1.65
cc_158 N_VPB_M1022_b N_A_1067_107#_c_633_n 0.00362066f $X=-0.33 $Y=1.885 $X2=1.2
+ $Y2=1.65
cc_159 N_VPB_M1022_b N_A_1067_107#_c_634_n 0.00308339f $X=-0.33 $Y=1.885
+ $X2=0.72 $Y2=1.985
cc_160 N_VPB_M1022_b N_A_1067_107#_c_624_n 0.0106281f $X=-0.33 $Y=1.885 $X2=2.59
+ $Y2=2.26
cc_161 N_VPB_M1022_b N_A_1067_107#_c_625_n 0.018f $X=-0.33 $Y=1.885 $X2=0.73
+ $Y2=1.65
cc_162 N_VPB_M1022_b N_A_1067_107#_c_637_n 0.0108646f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_163 N_VPB_M1022_b N_A_1570_457#_c_796_n 0.0391793f $X=-0.33 $Y=1.885
+ $X2=1.115 $Y2=1.58
cc_164 N_VPB_M1022_b N_A_1570_457#_c_785_n 0.0107032f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_165 N_VPB_M1022_b N_A_1570_457#_c_798_n 0.00333892f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_166 N_VPB_M1022_b N_A_1570_457#_c_799_n 0.0461064f $X=-0.33 $Y=1.885 $X2=0.88
+ $Y2=1.715
cc_167 N_VPB_M1022_b N_A_1570_457#_c_800_n 0.0130667f $X=-0.33 $Y=1.885 $X2=0.73
+ $Y2=1.715
cc_168 N_VPB_M1022_b N_A_1570_457#_c_801_n 0.00805484f $X=-0.33 $Y=1.885
+ $X2=2.62 $Y2=2.075
cc_169 N_VPB_M1022_b N_A_1570_457#_c_802_n 0.0099651f $X=-0.33 $Y=1.885 $X2=1.68
+ $Y2=1.65
cc_170 N_VPB_M1022_b N_A_1570_457#_c_793_n 0.0781888f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_171 N_VPB_M1022_b N_A_1570_457#_c_795_n 0.0318112f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_172 N_VPB_M1022_b N_A_1570_457#_c_805_n 0.0329816f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_173 N_VPB_M1022_b N_A_1570_457#_c_806_n 0.0328533f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_174 N_VPB_c_124_p N_A_1570_457#_c_806_n 0.00198372f $X=19.44 $Y=4.07 $X2=0
+ $Y2=0
cc_175 N_VPB_M1022_b N_A_1726_453#_M1027_g 0.039192f $X=-0.33 $Y=1.885 $X2=2.585
+ $Y2=2.075
cc_176 N_VPB_c_124_p N_A_1726_453#_M1027_g 0.00197968f $X=19.44 $Y=4.07
+ $X2=2.585 $Y2=2.075
cc_177 N_VPB_M1022_b N_A_1726_453#_M1034_g 0.043758f $X=-0.33 $Y=1.885 $X2=2.655
+ $Y2=2.785
cc_178 N_VPB_M1022_b N_A_1726_453#_c_980_n 0.0832937f $X=-0.33 $Y=1.885
+ $X2=2.075 $Y2=1.58
cc_179 N_VPB_M1022_b N_A_1726_453#_c_981_n 0.00542303f $X=-0.33 $Y=1.885 $X2=1.2
+ $Y2=1.65
cc_180 N_VPB_M1022_b N_A_1726_453#_c_974_n 0.00826858f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_181 N_VPB_M1022_b N_A_1726_453#_M1030_g 0.0405532f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_182 N_VPB_M1022_b N_A_1726_453#_c_976_n 0.0345455f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_183 N_VPB_M1022_b N_CLK_c_1076_n 0.039688f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=2.24
cc_184 N_VPB_M1022_b N_CLK_c_1073_n 0.0503445f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_185 N_VPB_M1022_b CLK 0.0029637f $X=-0.33 $Y=1.885 $X2=2.585 $Y2=2.075
cc_186 N_VPB_M1022_b N_A_2789_147#_M1031_g 0.0212351f $X=-0.33 $Y=1.885
+ $X2=2.585 $Y2=2.075
cc_187 N_VPB_M1022_b N_A_2789_147#_c_1122_n 0.0404867f $X=-0.33 $Y=1.885
+ $X2=2.585 $Y2=0.745
cc_188 N_VPB_M1022_b N_A_2789_147#_M1009_g 0.0433126f $X=-0.33 $Y=1.885
+ $X2=2.075 $Y2=1.58
cc_189 VPB N_A_2789_147#_M1009_g 6.05038e-19 $X=0 $Y=3.955 $X2=2.075 $Y2=1.58
cc_190 N_VPB_c_124_p N_A_2789_147#_M1009_g 0.0046353f $X=19.44 $Y=4.07 $X2=2.075
+ $Y2=1.58
cc_191 N_VPB_M1022_b N_A_2789_147#_M1033_g 0.0430356f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_192 N_VPB_M1022_b N_A_2789_147#_c_1127_n 0.00650478f $X=-0.33 $Y=1.885
+ $X2=0.73 $Y2=1.715
cc_193 N_VPB_M1022_b N_A_2789_147#_c_1128_n 0.0896971f $X=-0.33 $Y=1.885
+ $X2=0.88 $Y2=2.24
cc_194 N_VPB_M1022_b N_A_2789_147#_c_1118_n 0.00353265f $X=-0.33 $Y=1.885
+ $X2=2.62 $Y2=2.075
cc_195 N_VPB_M1022_b N_A_2789_147#_c_1130_n 0.00785648f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_196 N_VPB_M1022_b N_A_2789_147#_c_1131_n 0.010668f $X=-0.33 $Y=1.885 $X2=2.16
+ $Y2=1.65
cc_197 VPB N_A_2789_147#_c_1131_n 0.00303559f $X=0 $Y=3.955 $X2=2.16 $Y2=1.65
cc_198 N_VPB_c_124_p N_A_2789_147#_c_1131_n 0.0594445f $X=19.44 $Y=4.07 $X2=2.16
+ $Y2=1.65
cc_199 N_VPB_M1022_b N_A_2789_147#_c_1134_n 0.00162883f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_200 VPB N_A_2789_147#_c_1134_n 0.00142553f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_201 N_VPB_c_124_p N_A_2789_147#_c_1134_n 0.0260391f $X=19.44 $Y=4.07 $X2=0
+ $Y2=0
cc_202 N_VPB_M1022_b N_A_2789_147#_c_1137_n 0.00237972f $X=-0.33 $Y=1.885
+ $X2=0.73 $Y2=1.985
cc_203 N_VPB_M1022_b N_A_2789_147#_c_1138_n 0.00959984f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_204 N_VPB_M1022_b N_A_2789_147#_c_1139_n 0.00242348f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_205 N_VPB_M1022_b N_A_2789_147#_c_1120_n 0.0558009f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_206 N_VPB_M1022_b N_A_2518_445#_M1015_g 0.113686f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_207 VPB N_A_2518_445#_M1015_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_208 N_VPB_c_124_p N_A_2518_445#_M1015_g 0.0158724f $X=19.44 $Y=4.07 $X2=0
+ $Y2=0
cc_209 N_VPB_M1022_b N_A_2518_445#_c_1231_n 0.00507357f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_210 N_VPB_M1022_b N_A_2518_445#_c_1232_n 0.00453094f $X=-0.33 $Y=1.885
+ $X2=1.115 $Y2=1.58
cc_211 N_VPB_M1022_b N_A_2518_445#_c_1225_n 2.27616e-19 $X=-0.33 $Y=1.885
+ $X2=2.555 $Y2=1.58
cc_212 N_VPB_M1022_b N_A_2518_445#_c_1234_n 0.0251435f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_213 N_VPB_M1022_b N_A_2518_445#_c_1235_n 3.45447e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_214 N_VPB_M1022_b N_A_2518_445#_c_1227_n 0.0126175f $X=-0.33 $Y=1.885
+ $X2=2.62 $Y2=2.785
cc_215 N_VPB_M1022_b N_A_3531_107#_M1021_g 0.0437682f $X=-0.33 $Y=1.885
+ $X2=2.655 $Y2=2.785
cc_216 VPB N_A_3531_107#_M1021_g 0.00970178f $X=0 $Y=3.955 $X2=2.655 $Y2=2.785
cc_217 N_VPB_c_124_p N_A_3531_107#_M1021_g 0.0167165f $X=19.44 $Y=4.07 $X2=2.655
+ $Y2=2.785
cc_218 N_VPB_M1022_b N_A_3531_107#_c_1313_n 0.0219424f $X=-0.33 $Y=1.885
+ $X2=2.555 $Y2=1.58
cc_219 N_VPB_M1022_b N_A_3531_107#_c_1307_n 0.00189001f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_220 N_VPB_M1022_b N_A_3531_107#_c_1308_n 0.00931119f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_221 N_VPB_M1022_b N_A_3531_107#_c_1309_n 0.0252772f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_222 N_VPB_M1022_b N_A_3531_107#_c_1317_n 0.00501784f $X=-0.33 $Y=1.885
+ $X2=0.88 $Y2=1.085
cc_223 N_VPB_M1022_b N_VPWR_c_1343_n 0.0386849f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1343_n 0.00166879f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_225 N_VPB_c_124_p N_VPWR_c_1343_n 0.0254284f $X=19.44 $Y=4.07 $X2=0 $Y2=0
cc_226 N_VPB_M1022_b N_VPWR_c_1346_n 0.00124766f $X=-0.33 $Y=1.885 $X2=0.88
+ $Y2=1.085
cc_227 VPB N_VPWR_c_1346_n 0.00394105f $X=0 $Y=3.955 $X2=0.88 $Y2=1.085
cc_228 N_VPB_c_124_p N_VPWR_c_1346_n 0.0472737f $X=19.44 $Y=4.07 $X2=0.88
+ $Y2=1.085
cc_229 N_VPB_M1022_b N_VPWR_c_1349_n 0.0160113f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1349_n 0.00279351f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_231 N_VPB_c_124_p N_VPWR_c_1349_n 0.0460952f $X=19.44 $Y=4.07 $X2=0 $Y2=0
cc_232 N_VPB_M1022_b N_VPWR_c_1352_n 0.030529f $X=-0.33 $Y=1.885 $X2=0.73
+ $Y2=1.75
cc_233 VPB N_VPWR_c_1352_n 0.00166879f $X=0 $Y=3.955 $X2=0.73 $Y2=1.75
cc_234 N_VPB_c_124_p N_VPWR_c_1352_n 0.0254284f $X=19.44 $Y=4.07 $X2=0.73
+ $Y2=1.75
cc_235 N_VPB_M1022_b N_VPWR_c_1355_n 0.0139765f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1355_n 0.00310675f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_237 N_VPB_c_124_p N_VPWR_c_1355_n 0.0429406f $X=19.44 $Y=4.07 $X2=0 $Y2=0
cc_238 N_VPB_M1022_b N_VPWR_c_1358_n 0.0448816f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1358_n 0.00166879f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_240 N_VPB_c_124_p N_VPWR_c_1358_n 0.0254284f $X=19.44 $Y=4.07 $X2=0 $Y2=0
cc_241 N_VPB_M1022_b N_VPWR_c_1361_n 0.0419673f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1361_n 0.00219064f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_243 N_VPB_c_124_p N_VPWR_c_1361_n 0.0301848f $X=19.44 $Y=4.07 $X2=0 $Y2=0
cc_244 N_VPB_M1022_b N_VPWR_c_1364_n 0.217853f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1364_n 2.09908f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_246 N_VPB_c_124_p N_VPWR_c_1364_n 0.0919375f $X=19.44 $Y=4.07 $X2=0 $Y2=0
cc_247 N_VPB_M1022_b N_A_268_659#_c_1472_n 0.00567152f $X=-0.33 $Y=1.885
+ $X2=2.585 $Y2=2.075
cc_248 VPB N_A_268_659#_c_1472_n 5.14916e-19 $X=0 $Y=3.955 $X2=2.585 $Y2=2.075
cc_249 N_VPB_c_124_p N_A_268_659#_c_1472_n 0.00887752f $X=19.44 $Y=4.07
+ $X2=2.585 $Y2=2.075
cc_250 N_VPB_M1022_b N_A_268_659#_c_1475_n 0.0326525f $X=-0.33 $Y=1.885
+ $X2=2.585 $Y2=0.745
cc_251 N_VPB_M1022_b N_A_268_659#_c_1476_n 0.00846447f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_252 N_VPB_M1022_b N_A_268_659#_c_1477_n 0.00626963f $X=-0.33 $Y=1.885
+ $X2=2.655 $Y2=3.505
cc_253 N_VPB_M1022_b N_A_581_659#_c_1504_n 0.00611326f $X=-0.33 $Y=1.885
+ $X2=2.585 $Y2=2.075
cc_254 N_VPB_M1022_b N_A_581_659#_c_1505_n 0.0125431f $X=-0.33 $Y=1.885
+ $X2=2.585 $Y2=0.745
cc_255 VPB N_A_581_659#_c_1505_n 0.00266024f $X=0 $Y=3.955 $X2=2.585 $Y2=0.745
cc_256 N_VPB_c_124_p N_A_581_659#_c_1505_n 0.047534f $X=19.44 $Y=4.07 $X2=2.585
+ $Y2=0.745
cc_257 N_VPB_M1022_b N_A_581_659#_c_1508_n 0.00168334f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_258 VPB N_A_581_659#_c_1508_n 0.00109933f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_259 N_VPB_c_124_p N_A_581_659#_c_1508_n 0.0193841f $X=19.44 $Y=4.07 $X2=0
+ $Y2=0
cc_260 N_VPB_M1022_b N_A_581_659#_c_1511_n 8.79395e-19 $X=-0.33 $Y=1.885
+ $X2=2.655 $Y2=3.505
cc_261 N_VPB_M1022_b N_A_581_659#_c_1512_n 0.0121346f $X=-0.33 $Y=1.885
+ $X2=2.655 $Y2=3.505
cc_262 N_VPB_M1022_b N_A_581_659#_c_1513_n 0.00321111f $X=-0.33 $Y=1.885
+ $X2=1.595 $Y2=1.58
cc_263 N_VPB_M1022_b N_A_567_107#_c_1551_n 0.00993279f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_264 N_VPB_M1022_b N_A_567_107#_c_1563_n 0.0169185f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=1.58
cc_265 N_VPB_M1022_b N_A_567_107#_c_1564_n 0.0015486f $X=-0.33 $Y=1.885
+ $X2=2.555 $Y2=1.58
cc_266 N_VPB_M1022_b N_A_567_107#_c_1565_n 0.0205304f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=1.75
cc_267 VPB N_A_567_107#_c_1565_n 0.00576593f $X=0 $Y=3.955 $X2=0.72 $Y2=1.75
cc_268 N_VPB_c_124_p N_A_567_107#_c_1565_n 0.104385f $X=19.44 $Y=4.07 $X2=0.72
+ $Y2=1.75
cc_269 N_VPB_M1022_b N_A_567_107#_c_1568_n 0.00306127f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_270 VPB N_A_567_107#_c_1568_n 0.00110147f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_271 N_VPB_c_124_p N_A_567_107#_c_1568_n 0.0223208f $X=19.44 $Y=4.07 $X2=0
+ $Y2=0
cc_272 N_VPB_M1022_b N_A_567_107#_c_1552_n 0.00376788f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_273 N_VPB_M1022_b N_A_567_107#_c_1572_n 0.0112807f $X=-0.33 $Y=1.885 $X2=2.62
+ $Y2=2.075
cc_274 N_VPB_M1022_b N_A_567_107#_c_1573_n 0.0126397f $X=-0.33 $Y=1.885 $X2=2.16
+ $Y2=1.65
cc_275 VPB N_A_567_107#_c_1573_n 0.00315096f $X=0 $Y=3.955 $X2=2.16 $Y2=1.65
cc_276 N_VPB_c_124_p N_A_567_107#_c_1573_n 0.0297641f $X=19.44 $Y=4.07 $X2=2.16
+ $Y2=1.65
cc_277 N_VPB_M1022_b N_A_567_107#_c_1576_n 0.00150615f $X=-0.33 $Y=1.885
+ $X2=2.59 $Y2=1.75
cc_278 VPB N_A_567_107#_c_1576_n 3.38114e-19 $X=0 $Y=3.955 $X2=2.59 $Y2=1.75
cc_279 N_VPB_c_124_p N_A_567_107#_c_1576_n 0.00328434f $X=19.44 $Y=4.07 $X2=2.59
+ $Y2=1.75
cc_280 N_VPB_M1022_b N_A_567_107#_c_1579_n 0.0136195f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_281 VPB N_A_567_107#_c_1579_n 6.59548e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_282 N_VPB_c_124_p N_A_567_107#_c_1579_n 0.00641695f $X=19.44 $Y=4.07 $X2=0
+ $Y2=0
cc_283 N_VPB_M1022_b N_A_2365_445#_c_1742_n 0.0344682f $X=-0.33 $Y=1.885
+ $X2=2.585 $Y2=2.075
cc_284 N_VPB_M1022_b N_A_2365_445#_c_1743_n 0.0336338f $X=-0.33 $Y=1.885
+ $X2=2.585 $Y2=0.745
cc_285 VPB N_A_2365_445#_c_1743_n 0.00750194f $X=0 $Y=3.955 $X2=2.585 $Y2=0.745
cc_286 N_VPB_c_124_p N_A_2365_445#_c_1743_n 0.146889f $X=19.44 $Y=4.07 $X2=2.585
+ $Y2=0.745
cc_287 N_VPB_M1022_b N_A_2365_445#_c_1746_n 0.00520177f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_288 VPB N_A_2365_445#_c_1746_n 0.00110147f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_289 N_VPB_c_124_p N_A_2365_445#_c_1746_n 0.0223208f $X=19.44 $Y=4.07 $X2=0
+ $Y2=0
cc_290 N_VPB_M1022_b N_A_2365_445#_c_1749_n 0.0178784f $X=-0.33 $Y=1.885
+ $X2=2.655 $Y2=3.505
cc_291 N_VPB_M1022_b N_Q_c_1783_n 0.00951539f $X=-0.33 $Y=1.885 $X2=2.585
+ $Y2=2.075
cc_292 N_VPB_M1022_b N_Q_c_1781_n 0.00534059f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_293 N_VPB_M1022_b N_Q_c_1785_n 0.0207182f $X=-0.33 $Y=1.885 $X2=2.425
+ $Y2=1.65
cc_294 N_VPB_M1022_b N_Q_N_c_1809_n 0.0667138f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_295 VPB N_Q_N_c_1809_n 0.00106225f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_296 N_VPB_c_124_p N_Q_N_c_1809_n 0.0175015f $X=19.44 $Y=4.07 $X2=0 $Y2=0
cc_297 N_SCE_M1022_g N_SCD_M1019_g 0.0100646f $X=0.665 $Y=2.785 $X2=0 $Y2=0
cc_298 N_SCE_M1028_g N_SCD_M1019_g 0.0756274f $X=1.095 $Y=0.745 $X2=0 $Y2=0
cc_299 N_SCE_M1020_g N_SCD_M1019_g 0.170505f $X=2.585 $Y=0.745 $X2=0 $Y2=0
cc_300 N_SCE_M1018_g N_SCD_M1019_g 0.036853f $X=2.655 $Y=3.505 $X2=0 $Y2=0
cc_301 N_SCE_c_314_p N_SCD_M1019_g 0.00473466f $X=2.59 $Y=2.26 $X2=0 $Y2=0
cc_302 N_SCE_c_302_n N_SCD_M1019_g 0.0328322f $X=2.425 $Y=1.65 $X2=0 $Y2=0
cc_303 N_SCE_M1022_g N_SCD_c_374_n 0.00343891f $X=0.665 $Y=2.785 $X2=0 $Y2=0
cc_304 N_SCE_M1020_g N_SCD_c_374_n 0.00161964f $X=2.585 $Y=0.745 $X2=0 $Y2=0
cc_305 N_SCE_c_301_n N_SCD_c_374_n 0.00406564f $X=0.73 $Y=1.715 $X2=0 $Y2=0
cc_306 N_SCE_c_314_p N_SCD_c_374_n 0.0176637f $X=2.59 $Y=2.26 $X2=0 $Y2=0
cc_307 N_SCE_c_302_n N_SCD_c_374_n 0.0298f $X=2.425 $Y=1.65 $X2=0 $Y2=0
cc_308 N_SCE_c_321_p N_SCD_c_374_n 0.00816368f $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_309 N_SCE_M1020_g N_A_30_515#_M1013_g 0.0148492f $X=2.585 $Y=0.745 $X2=0
+ $Y2=0
cc_310 N_SCE_M1020_g N_A_30_515#_c_399_n 0.0105883f $X=2.585 $Y=0.745 $X2=0
+ $Y2=0
cc_311 N_SCE_c_309_n N_A_30_515#_c_399_n 0.0294298f $X=2.59 $Y=2.26 $X2=0 $Y2=0
cc_312 N_SCE_c_314_p N_A_30_515#_c_399_n 0.00491742f $X=2.59 $Y=2.26 $X2=0 $Y2=0
cc_313 N_SCE_M1018_g N_A_30_515#_c_411_n 0.0294298f $X=2.655 $Y=3.505 $X2=0
+ $Y2=0
cc_314 N_SCE_c_301_n N_A_30_515#_c_400_n 0.0132841f $X=0.73 $Y=1.715 $X2=9.84
+ $Y2=0.057
cc_315 N_SCE_M1028_g N_A_30_515#_c_402_n 0.015895f $X=1.095 $Y=0.745 $X2=0 $Y2=0
cc_316 N_SCE_c_301_n N_A_30_515#_c_402_n 0.0174543f $X=0.73 $Y=1.715 $X2=0 $Y2=0
cc_317 N_SCE_M1020_g N_A_30_515#_c_404_n 0.032196f $X=2.585 $Y=0.745 $X2=0 $Y2=0
cc_318 SCE N_A_30_515#_c_404_n 0.0216226f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_319 N_SCE_c_301_n N_A_30_515#_c_404_n 0.0249442f $X=0.73 $Y=1.715 $X2=0 $Y2=0
cc_320 N_SCE_c_302_n N_A_30_515#_c_404_n 0.0941555f $X=2.425 $Y=1.65 $X2=0 $Y2=0
cc_321 N_SCE_c_334_p N_A_30_515#_c_404_n 0.00145487f $X=0.73 $Y=1.75 $X2=0 $Y2=0
cc_322 N_SCE_M1022_g N_A_30_515#_c_412_n 0.0128915f $X=0.665 $Y=2.785 $X2=0
+ $Y2=0
cc_323 N_SCE_c_301_n N_A_30_515#_c_405_n 0.0419427f $X=0.73 $Y=1.715 $X2=0 $Y2=0
cc_324 N_SCE_c_321_p N_A_30_515#_c_405_n 0.0239795f $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_325 N_SCE_c_334_p N_A_30_515#_c_405_n 0.0108273f $X=0.73 $Y=1.75 $X2=0 $Y2=0
cc_326 N_SCE_c_301_n N_A_30_515#_c_431_n 0.0113796f $X=0.73 $Y=1.715 $X2=0 $Y2=0
cc_327 N_SCE_c_334_p N_A_30_515#_c_431_n 0.0202678f $X=0.73 $Y=1.75 $X2=0 $Y2=0
cc_328 N_SCE_M1020_g N_A_30_515#_c_433_n 0.00258478f $X=2.585 $Y=0.745 $X2=0
+ $Y2=0
cc_329 SCE N_A_30_515#_c_433_n 0.00969702f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_330 N_SCE_c_314_p N_A_30_515#_c_433_n 0.00431225f $X=2.59 $Y=2.26 $X2=0 $Y2=0
cc_331 N_SCE_M1020_g N_A_30_515#_c_406_n 0.054187f $X=2.585 $Y=0.745 $X2=0 $Y2=0
cc_332 SCE N_A_30_515#_c_406_n 6.89294e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_333 N_SCE_c_314_p N_A_30_515#_c_406_n 4.5236e-19 $X=2.59 $Y=2.26 $X2=0 $Y2=0
cc_334 N_SCE_M1022_g N_VPWR_c_1343_n 0.0406668f $X=0.665 $Y=2.785 $X2=0 $Y2=0
cc_335 N_SCE_c_301_n N_VPWR_c_1343_n 0.010668f $X=0.73 $Y=1.715 $X2=0 $Y2=0
cc_336 N_SCE_c_321_p N_VPWR_c_1343_n 0.0108252f $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_337 N_SCE_M1018_g N_VPWR_c_1346_n 0.0226897f $X=2.655 $Y=3.505 $X2=0 $Y2=0
cc_338 N_SCE_M1022_g N_VPWR_c_1364_n 0.00623382f $X=0.665 $Y=2.785 $X2=0 $Y2=0
cc_339 N_SCE_M1018_g N_VPWR_c_1364_n 0.00436375f $X=2.655 $Y=3.505 $X2=0 $Y2=0
cc_340 N_SCE_M1018_g N_A_268_659#_c_1475_n 0.0348112f $X=2.655 $Y=3.505 $X2=0.24
+ $Y2=0
cc_341 N_SCE_c_309_n N_A_268_659#_c_1475_n 0.0030014f $X=2.59 $Y=2.26 $X2=0.24
+ $Y2=0
cc_342 N_SCE_c_314_p N_A_268_659#_c_1475_n 0.0238596f $X=2.59 $Y=2.26 $X2=0.24
+ $Y2=0
cc_343 N_SCE_M1022_g N_A_268_659#_c_1476_n 3.97663e-19 $X=0.665 $Y=2.785 $X2=0
+ $Y2=0
cc_344 N_SCE_M1018_g N_A_268_659#_c_1477_n 0.00542319f $X=2.655 $Y=3.505 $X2=0
+ $Y2=0
cc_345 N_SCE_M1018_g N_A_581_659#_c_1504_n 0.00738257f $X=2.655 $Y=3.505 $X2=0
+ $Y2=0
cc_346 N_SCE_M1018_g N_A_581_659#_c_1508_n 0.00418082f $X=2.655 $Y=3.505 $X2=0
+ $Y2=0
cc_347 N_SCE_M1020_g N_A_567_107#_c_1551_n 0.00154313f $X=2.585 $Y=0.745
+ $X2=19.44 $Y2=0
cc_348 N_SCE_c_309_n N_A_567_107#_c_1551_n 9.01204e-19 $X=2.59 $Y=2.26 $X2=19.44
+ $Y2=0
cc_349 N_SCE_c_309_n N_A_567_107#_c_1584_n 5.89345e-19 $X=2.59 $Y=2.26 $X2=0
+ $Y2=0
cc_350 N_SCE_M1020_g N_A_567_107#_c_1559_n 0.0140663f $X=2.585 $Y=0.745 $X2=0
+ $Y2=0
cc_351 N_SCE_M1028_g N_VGND_c_1822_n 0.0358184f $X=1.095 $Y=0.745 $X2=0 $Y2=0
cc_352 N_SCE_M1020_g N_VGND_c_1822_n 0.00407355f $X=2.585 $Y=0.745 $X2=0 $Y2=0
cc_353 N_SCE_M1028_g N_VGND_c_1836_n 0.00644701f $X=1.095 $Y=0.745 $X2=0 $Y2=0
cc_354 N_SCE_M1020_g N_VGND_c_1836_n 0.0179728f $X=2.585 $Y=0.745 $X2=0 $Y2=0
cc_355 N_SCE_c_301_n N_VGND_c_1836_n 0.00335051f $X=0.73 $Y=1.715 $X2=0 $Y2=0
cc_356 N_SCD_M1019_g N_A_30_515#_c_404_n 0.0271407f $X=1.875 $Y=0.745 $X2=0
+ $Y2=0
cc_357 N_SCD_M1019_g N_VPWR_c_1343_n 0.00892352f $X=1.875 $Y=0.745 $X2=0 $Y2=0
cc_358 N_SCD_M1019_g N_VPWR_c_1346_n 0.0259397f $X=1.875 $Y=0.745 $X2=0 $Y2=0
cc_359 N_SCD_M1019_g N_VPWR_c_1364_n 0.00499547f $X=1.875 $Y=0.745 $X2=0 $Y2=0
cc_360 N_SCD_M1019_g N_A_268_659#_c_1472_n 0.010394f $X=1.875 $Y=0.745 $X2=0
+ $Y2=0
cc_361 N_SCD_M1019_g N_A_268_659#_c_1475_n 0.0361142f $X=1.875 $Y=0.745 $X2=0.24
+ $Y2=0
cc_362 N_SCD_c_374_n N_A_268_659#_c_1475_n 0.0132f $X=1.81 $Y=2.015 $X2=0.24
+ $Y2=0
cc_363 N_SCD_M1019_g N_A_567_107#_c_1559_n 0.0017125f $X=1.875 $Y=0.745 $X2=0
+ $Y2=0
cc_364 N_SCD_M1019_g N_VGND_c_1822_n 0.0445503f $X=1.875 $Y=0.745 $X2=0 $Y2=0
cc_365 N_SCD_M1019_g N_VGND_c_1836_n 0.00461913f $X=1.875 $Y=0.745 $X2=0 $Y2=0
cc_366 N_A_30_515#_M1013_g N_D_M1014_g 0.049085f $X=3.365 $Y=0.745 $X2=0 $Y2=0
cc_367 N_A_30_515#_c_411_n N_D_M1007_g 0.0407044f $X=3.985 $Y=2.61 $X2=0 $Y2=0
cc_368 N_A_30_515#_c_399_n D 0.00163075f $X=3.365 $Y=2.36 $X2=0 $Y2=0
cc_369 N_A_30_515#_c_411_n D 2.95881e-19 $X=3.985 $Y=2.61 $X2=0 $Y2=0
cc_370 N_A_30_515#_c_406_n D 5.09607e-19 $X=3.23 $Y=1.34 $X2=0 $Y2=0
cc_371 N_A_30_515#_c_411_n N_D_c_486_n 0.00880255f $X=3.985 $Y=2.61 $X2=0 $Y2=0
cc_372 N_A_30_515#_c_406_n N_D_c_486_n 0.049085f $X=3.23 $Y=1.34 $X2=0 $Y2=0
cc_373 N_A_30_515#_c_412_n N_VPWR_c_1343_n 0.0283751f $X=0.275 $Y=2.785 $X2=0
+ $Y2=0
cc_374 N_A_30_515#_M1016_g N_VPWR_c_1364_n 0.0139661f $X=3.985 $Y=3.2 $X2=0
+ $Y2=0
cc_375 N_A_30_515#_c_411_n N_VPWR_c_1364_n 0.00130243f $X=3.985 $Y=2.61 $X2=0
+ $Y2=0
cc_376 N_A_30_515#_c_412_n N_VPWR_c_1364_n 0.0142526f $X=0.275 $Y=2.785 $X2=0
+ $Y2=0
cc_377 N_A_30_515#_M1016_g N_A_268_659#_c_1475_n 0.00227932f $X=3.985 $Y=3.2
+ $X2=0.24 $Y2=0
cc_378 N_A_30_515#_c_411_n N_A_268_659#_c_1475_n 0.0246004f $X=3.985 $Y=2.61
+ $X2=0.24 $Y2=0
cc_379 N_A_30_515#_M1016_g N_A_268_659#_c_1477_n 9.43117e-19 $X=3.985 $Y=3.2
+ $X2=0 $Y2=0
cc_380 N_A_30_515#_M1016_g N_A_581_659#_c_1504_n 0.00159021f $X=3.985 $Y=3.2
+ $X2=0 $Y2=0
cc_381 N_A_30_515#_M1016_g N_A_581_659#_c_1505_n 0.00445056f $X=3.985 $Y=3.2
+ $X2=0.24 $Y2=0
cc_382 N_A_30_515#_M1016_g N_A_581_659#_c_1511_n 0.031384f $X=3.985 $Y=3.2 $X2=0
+ $Y2=0
cc_383 N_A_30_515#_c_411_n N_A_581_659#_c_1511_n 6.87965e-19 $X=3.985 $Y=2.61
+ $X2=0 $Y2=0
cc_384 N_A_30_515#_c_411_n N_A_581_659#_c_1512_n 0.0127791f $X=3.985 $Y=2.61
+ $X2=0 $Y2=0
cc_385 N_A_30_515#_c_411_n N_A_581_659#_c_1521_n 0.0140854f $X=3.985 $Y=2.61
+ $X2=19.44 $Y2=0
cc_386 N_A_30_515#_M1013_g N_A_567_107#_c_1550_n 0.0265218f $X=3.365 $Y=0.745
+ $X2=0 $Y2=0
cc_387 N_A_30_515#_c_433_n N_A_567_107#_c_1550_n 0.013285f $X=3.23 $Y=1.34 $X2=0
+ $Y2=0
cc_388 N_A_30_515#_M1013_g N_A_567_107#_c_1551_n 0.00291227f $X=3.365 $Y=0.745
+ $X2=19.44 $Y2=0
cc_389 N_A_30_515#_c_399_n N_A_567_107#_c_1551_n 0.0206619f $X=3.365 $Y=2.36
+ $X2=19.44 $Y2=0
cc_390 N_A_30_515#_c_433_n N_A_567_107#_c_1551_n 0.0458459f $X=3.23 $Y=1.34
+ $X2=19.44 $Y2=0
cc_391 N_A_30_515#_c_406_n N_A_567_107#_c_1551_n 0.0215989f $X=3.23 $Y=1.34
+ $X2=19.44 $Y2=0
cc_392 N_A_30_515#_c_411_n N_A_567_107#_c_1563_n 0.0272648f $X=3.985 $Y=2.61
+ $X2=19.44 $Y2=0
cc_393 N_A_30_515#_c_399_n N_A_567_107#_c_1584_n 0.00165248f $X=3.365 $Y=2.36
+ $X2=0 $Y2=0
cc_394 N_A_30_515#_c_411_n N_A_567_107#_c_1584_n 0.0102529f $X=3.985 $Y=2.61
+ $X2=0 $Y2=0
cc_395 N_A_30_515#_M1016_g N_A_567_107#_c_1564_n 0.0104371f $X=3.985 $Y=3.2
+ $X2=9.84 $Y2=0
cc_396 N_A_30_515#_M1013_g N_A_567_107#_c_1559_n 0.010846f $X=3.365 $Y=0.745
+ $X2=0 $Y2=0
cc_397 N_A_30_515#_c_404_n N_A_567_107#_c_1559_n 0.0191696f $X=3.065 $Y=1.26
+ $X2=0 $Y2=0
cc_398 N_A_30_515#_c_433_n N_A_567_107#_c_1559_n 0.00585457f $X=3.23 $Y=1.34
+ $X2=0 $Y2=0
cc_399 N_A_30_515#_c_406_n N_A_567_107#_c_1559_n 0.00209008f $X=3.23 $Y=1.34
+ $X2=0 $Y2=0
cc_400 N_A_30_515#_c_402_n N_VGND_c_1822_n 0.0360627f $X=0.705 $Y=0.745 $X2=0
+ $Y2=0
cc_401 N_A_30_515#_c_404_n N_VGND_c_1822_n 0.0686854f $X=3.065 $Y=1.26 $X2=0
+ $Y2=0
cc_402 N_A_30_515#_M1013_g N_VGND_c_1824_n 0.00394291f $X=3.365 $Y=0.745 $X2=0
+ $Y2=0
cc_403 N_A_30_515#_M1013_g N_VGND_c_1836_n 0.0154688f $X=3.365 $Y=0.745 $X2=0
+ $Y2=0
cc_404 N_A_30_515#_c_400_n N_VGND_c_1836_n 0.00861761f $X=0.54 $Y=1.26 $X2=0
+ $Y2=0
cc_405 N_A_30_515#_c_401_n N_VGND_c_1836_n 0.00679505f $X=0.28 $Y=1.26 $X2=0
+ $Y2=0
cc_406 N_A_30_515#_c_402_n N_VGND_c_1836_n 0.025902f $X=0.705 $Y=0.745 $X2=0
+ $Y2=0
cc_407 N_A_30_515#_c_404_n N_VGND_c_1836_n 0.0330809f $X=3.065 $Y=1.26 $X2=0
+ $Y2=0
cc_408 N_A_30_515#_c_433_n N_VGND_c_1836_n 6.24171e-19 $X=3.23 $Y=1.34 $X2=0
+ $Y2=0
cc_409 N_D_c_486_n N_A_1124_81#_c_526_n 0.00965342f $X=4.765 $Y=1.475 $X2=0
+ $Y2=0
cc_410 N_D_M1007_g N_A_1124_81#_c_528_n 0.00965342f $X=4.765 $Y=3.2 $X2=0.24
+ $Y2=0
cc_411 N_D_c_486_n N_A_1067_107#_c_619_n 0.00168404f $X=4.765 $Y=1.475 $X2=0
+ $Y2=0
cc_412 N_D_c_486_n N_A_1067_107#_c_622_n 6.20443e-19 $X=4.765 $Y=1.475 $X2=0
+ $Y2=0
cc_413 N_D_M1007_g N_A_1067_107#_c_625_n 0.0076562f $X=4.765 $Y=3.2 $X2=0 $Y2=0
cc_414 N_D_c_486_n N_A_1067_107#_c_625_n 0.00259017f $X=4.765 $Y=1.475 $X2=0
+ $Y2=0
cc_415 N_D_M1007_g N_VPWR_c_1364_n 0.0163577f $X=4.765 $Y=3.2 $X2=0 $Y2=0
cc_416 N_D_M1007_g N_A_581_659#_c_1511_n 0.00101205f $X=4.765 $Y=3.2 $X2=0 $Y2=0
cc_417 N_D_M1007_g N_A_581_659#_c_1512_n 0.0313041f $X=4.765 $Y=3.2 $X2=0 $Y2=0
cc_418 N_D_M1007_g N_A_581_659#_c_1513_n 0.0223196f $X=4.765 $Y=3.2 $X2=0 $Y2=0
cc_419 N_D_M1014_g N_A_567_107#_c_1550_n 0.00114434f $X=4.075 $Y=0.745 $X2=0
+ $Y2=0
cc_420 N_D_M1014_g N_A_567_107#_c_1551_n 0.0105134f $X=4.075 $Y=0.745 $X2=19.44
+ $Y2=0
cc_421 D N_A_567_107#_c_1551_n 0.0356085f $X=4.475 $Y=1.21 $X2=19.44 $Y2=0
cc_422 N_D_M1007_g N_A_567_107#_c_1563_n 0.0344777f $X=4.765 $Y=3.2 $X2=19.44
+ $Y2=0
cc_423 D N_A_567_107#_c_1563_n 0.0398703f $X=4.475 $Y=1.21 $X2=19.44 $Y2=0
cc_424 N_D_c_486_n N_A_567_107#_c_1563_n 0.00708377f $X=4.765 $Y=1.475 $X2=19.44
+ $Y2=0
cc_425 N_D_M1007_g N_A_567_107#_c_1564_n 0.0161287f $X=4.765 $Y=3.2 $X2=9.84
+ $Y2=0
cc_426 N_D_M1007_g N_A_567_107#_c_1565_n 0.0159131f $X=4.765 $Y=3.2 $X2=9.84
+ $Y2=0.057
cc_427 N_D_M1014_g N_A_567_107#_c_1552_n 0.00295602f $X=4.075 $Y=0.745 $X2=0
+ $Y2=0
cc_428 N_D_M1007_g N_A_567_107#_c_1552_n 0.0203797f $X=4.765 $Y=3.2 $X2=0 $Y2=0
cc_429 D N_A_567_107#_c_1552_n 0.0470271f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_430 N_D_c_486_n N_A_567_107#_c_1552_n 0.0309296f $X=4.765 $Y=1.475 $X2=0
+ $Y2=0
cc_431 N_D_M1014_g N_A_567_107#_c_1559_n 0.00119732f $X=4.075 $Y=0.745 $X2=0
+ $Y2=0
cc_432 N_D_M1014_g N_VGND_c_1824_n 0.0628197f $X=4.075 $Y=0.745 $X2=0 $Y2=0
cc_433 D N_VGND_c_1824_n 0.0410075f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_434 N_D_c_486_n N_VGND_c_1824_n 0.0162034f $X=4.765 $Y=1.475 $X2=0 $Y2=0
cc_435 N_D_M1014_g N_VGND_c_1836_n 0.00309573f $X=4.075 $Y=0.745 $X2=0 $Y2=0
cc_436 D N_VGND_c_1836_n 0.00185728f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_437 N_D_c_486_n N_VGND_c_1836_n 0.00483963f $X=4.765 $Y=1.475 $X2=0 $Y2=0
cc_438 N_A_1124_81#_c_526_n N_A_1067_107#_c_618_n 0.0105049f $X=5.87 $Y=1.395
+ $X2=0 $Y2=0
cc_439 N_A_1124_81#_c_528_n N_A_1067_107#_M1001_g 0.0149116f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_440 N_A_1124_81#_c_534_n N_A_1067_107#_M1001_g 0.0424288f $X=7.74 $Y=2.43
+ $X2=0 $Y2=0
cc_441 N_A_1124_81#_c_537_n N_A_1067_107#_M1001_g 0.00724356f $X=7.91 $Y=2.98
+ $X2=0 $Y2=0
cc_442 N_A_1124_81#_c_540_n N_A_1067_107#_M1001_g 0.0110704f $X=7.825 $Y=2.22
+ $X2=0 $Y2=0
cc_443 N_A_1124_81#_c_526_n N_A_1067_107#_c_619_n 0.0162418f $X=5.87 $Y=1.395
+ $X2=0 $Y2=0
cc_444 N_A_1124_81#_c_528_n N_A_1067_107#_c_619_n 0.0127901f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_445 N_A_1124_81#_c_528_n N_A_1067_107#_c_620_n 0.0351046f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_446 N_A_1124_81#_c_528_n N_A_1067_107#_c_622_n 0.012965f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_447 N_A_1124_81#_M1002_d N_A_1067_107#_c_632_n 0.00132575f $X=8.35 $Y=2.895
+ $X2=0 $Y2=0
cc_448 N_A_1124_81#_c_528_n N_A_1067_107#_c_632_n 0.0232136f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_449 N_A_1124_81#_c_534_n N_A_1067_107#_c_632_n 0.0292887f $X=7.74 $Y=2.43
+ $X2=0 $Y2=0
cc_450 N_A_1124_81#_c_537_n N_A_1067_107#_c_632_n 0.0115624f $X=7.91 $Y=2.98
+ $X2=0 $Y2=0
cc_451 N_A_1124_81#_c_538_n N_A_1067_107#_c_632_n 0.0240122f $X=8.49 $Y=3.02
+ $X2=0 $Y2=0
cc_452 N_A_1124_81#_c_528_n N_A_1067_107#_c_624_n 0.0184114f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_453 N_A_1124_81#_c_528_n N_A_1067_107#_c_625_n 0.051011f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_454 N_A_1124_81#_c_529_n N_A_1570_457#_c_784_n 0.00214405f $X=8.7 $Y=2.135
+ $X2=0 $Y2=0
cc_455 N_A_1124_81#_c_530_n N_A_1570_457#_c_784_n 0.0119057f $X=8.78 $Y=1.11
+ $X2=0 $Y2=0
cc_456 N_A_1124_81#_c_536_n N_A_1570_457#_c_785_n 0.00777751f $X=8.615 $Y=2.22
+ $X2=0 $Y2=0
cc_457 N_A_1124_81#_c_529_n N_A_1570_457#_c_785_n 0.027316f $X=8.7 $Y=2.135
+ $X2=0 $Y2=0
cc_458 N_A_1124_81#_c_536_n N_A_1570_457#_c_798_n 0.0483258f $X=8.615 $Y=2.22
+ $X2=0 $Y2=0
cc_459 N_A_1124_81#_c_538_n N_A_1570_457#_c_798_n 0.0377283f $X=8.49 $Y=3.02
+ $X2=0 $Y2=0
cc_460 N_A_1124_81#_c_540_n N_A_1570_457#_c_798_n 0.0136431f $X=7.825 $Y=2.22
+ $X2=0 $Y2=0
cc_461 N_A_1124_81#_c_534_n N_A_1570_457#_c_799_n 2.50651e-19 $X=7.74 $Y=2.43
+ $X2=0 $Y2=0
cc_462 N_A_1124_81#_c_535_n N_A_1570_457#_c_799_n 0.00862831f $X=7.825 $Y=2.855
+ $X2=0 $Y2=0
cc_463 N_A_1124_81#_c_536_n N_A_1570_457#_c_799_n 0.0105349f $X=8.615 $Y=2.22
+ $X2=0 $Y2=0
cc_464 N_A_1124_81#_c_538_n N_A_1570_457#_c_799_n 0.00210336f $X=8.49 $Y=3.02
+ $X2=0 $Y2=0
cc_465 N_A_1124_81#_c_540_n N_A_1570_457#_c_799_n 0.0124065f $X=7.825 $Y=2.22
+ $X2=0 $Y2=0
cc_466 N_A_1124_81#_c_538_n N_A_1570_457#_c_820_n 0.00465552f $X=8.49 $Y=3.02
+ $X2=0 $Y2=0
cc_467 N_A_1124_81#_c_536_n N_A_1570_457#_c_805_n 0.0317233f $X=8.615 $Y=2.22
+ $X2=0 $Y2=0
cc_468 N_A_1124_81#_c_529_n N_A_1570_457#_c_805_n 0.00485086f $X=8.7 $Y=2.135
+ $X2=0 $Y2=0
cc_469 N_A_1124_81#_c_540_n N_A_1570_457#_c_805_n 6.26767e-19 $X=7.825 $Y=2.22
+ $X2=0 $Y2=0
cc_470 N_A_1124_81#_c_535_n N_A_1570_457#_c_806_n 0.00349903f $X=7.825 $Y=2.855
+ $X2=0 $Y2=0
cc_471 N_A_1124_81#_c_537_n N_A_1570_457#_c_806_n 0.00303619f $X=7.91 $Y=2.98
+ $X2=0 $Y2=0
cc_472 N_A_1124_81#_c_538_n N_A_1570_457#_c_806_n 0.0224614f $X=8.49 $Y=3.02
+ $X2=0 $Y2=0
cc_473 N_A_1124_81#_c_538_n N_A_1726_453#_M1027_g 0.010612f $X=8.49 $Y=3.02
+ $X2=0 $Y2=0
cc_474 N_A_1124_81#_c_536_n N_A_1726_453#_c_980_n 0.00903928f $X=8.615 $Y=2.22
+ $X2=0 $Y2=0
cc_475 N_A_1124_81#_c_536_n N_A_1726_453#_c_987_n 0.00458974f $X=8.615 $Y=2.22
+ $X2=0 $Y2=0
cc_476 N_A_1124_81#_c_529_n N_A_1726_453#_c_987_n 0.0306062f $X=8.7 $Y=2.135
+ $X2=0 $Y2=0
cc_477 N_A_1124_81#_c_536_n N_A_1726_453#_M1030_g 0.0026729f $X=8.615 $Y=2.22
+ $X2=0 $Y2=0
cc_478 N_A_1124_81#_c_529_n N_A_1726_453#_M1030_g 0.00979056f $X=8.7 $Y=2.135
+ $X2=0 $Y2=0
cc_479 N_A_1124_81#_c_530_n N_A_1726_453#_M1030_g 0.0130847f $X=8.78 $Y=1.11
+ $X2=0 $Y2=0
cc_480 N_A_1124_81#_c_528_n N_VPWR_c_1349_n 0.00417692f $X=6.095 $Y=2.605 $X2=0
+ $Y2=0
cc_481 N_A_1124_81#_c_528_n N_VPWR_c_1364_n 0.00751493f $X=6.095 $Y=2.605 $X2=0
+ $Y2=0
cc_482 N_A_1124_81#_c_538_n N_VPWR_c_1364_n 9.41913e-19 $X=8.49 $Y=3.02 $X2=0
+ $Y2=0
cc_483 N_A_1124_81#_c_528_n N_A_567_107#_c_1563_n 5.86391e-19 $X=6.095 $Y=2.605
+ $X2=19.44 $Y2=0
cc_484 N_A_1124_81#_c_528_n N_A_567_107#_c_1565_n 0.0144051f $X=6.095 $Y=2.605
+ $X2=9.84 $Y2=0.057
cc_485 N_A_1124_81#_c_526_n N_A_567_107#_c_1552_n 0.00578629f $X=5.87 $Y=1.395
+ $X2=0 $Y2=0
cc_486 N_A_1124_81#_c_526_n N_A_567_107#_c_1553_n 0.0127945f $X=5.87 $Y=1.395
+ $X2=0 $Y2=0
cc_487 N_A_1124_81#_c_526_n N_A_567_107#_c_1618_n 0.0372316f $X=5.87 $Y=1.395
+ $X2=0 $Y2=0
cc_488 N_A_1124_81#_c_528_n N_A_567_107#_c_1619_n 0.0589471f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_489 N_A_1124_81#_c_534_n N_A_567_107#_c_1619_n 0.0180402f $X=7.74 $Y=2.43
+ $X2=0 $Y2=0
cc_490 N_A_1124_81#_c_528_n N_A_567_107#_c_1621_n 0.0183722f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_491 N_A_1124_81#_c_526_n N_A_567_107#_c_1557_n 0.00991594f $X=5.87 $Y=1.395
+ $X2=0 $Y2=0
cc_492 N_A_1124_81#_c_528_n N_A_567_107#_c_1557_n 0.0101996f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_493 N_A_1124_81#_c_526_n N_A_567_107#_c_1624_n 0.00430069f $X=5.87 $Y=1.395
+ $X2=0 $Y2=0
cc_494 N_A_1124_81#_c_528_n N_A_567_107#_c_1624_n 0.00346669f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_495 N_A_1124_81#_c_528_n N_A_567_107#_c_1572_n 0.0292473f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_496 N_A_1124_81#_c_534_n N_A_567_107#_c_1572_n 0.0816365f $X=7.74 $Y=2.43
+ $X2=0 $Y2=0
cc_497 N_A_1124_81#_c_528_n N_A_567_107#_c_1628_n 0.00779832f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_498 N_A_1124_81#_c_528_n N_A_567_107#_c_1629_n 0.0208502f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_499 N_A_1124_81#_c_534_n N_A_567_107#_c_1629_n 0.0170247f $X=7.74 $Y=2.43
+ $X2=0 $Y2=0
cc_500 N_A_1124_81#_M1002_d N_A_567_107#_c_1573_n 0.00158821f $X=8.35 $Y=2.895
+ $X2=0 $Y2=0
cc_501 N_A_1124_81#_c_537_n N_A_567_107#_c_1573_n 0.00751529f $X=7.91 $Y=2.98
+ $X2=0 $Y2=0
cc_502 N_A_1124_81#_c_538_n N_A_567_107#_c_1573_n 0.0374343f $X=8.49 $Y=3.02
+ $X2=0 $Y2=0
cc_503 N_A_1124_81#_c_528_n N_A_567_107#_c_1634_n 0.0038041f $X=6.095 $Y=2.605
+ $X2=0 $Y2=0
cc_504 N_A_1124_81#_c_534_n N_A_567_107#_c_1576_n 0.0023352f $X=7.74 $Y=2.43
+ $X2=0 $Y2=0
cc_505 N_A_1124_81#_c_530_n N_A_567_107#_c_1561_n 0.0164174f $X=8.78 $Y=1.11
+ $X2=0 $Y2=0
cc_506 N_A_1124_81#_c_537_n A_1528_579# 0.00315232f $X=7.91 $Y=2.98 $X2=0 $Y2=0
cc_507 N_A_1124_81#_c_526_n N_VGND_c_1826_n 0.0112479f $X=5.87 $Y=1.395 $X2=0
+ $Y2=0
cc_508 N_A_1124_81#_c_528_n N_VGND_c_1826_n 9.41844e-19 $X=6.095 $Y=2.605 $X2=0
+ $Y2=0
cc_509 N_A_1124_81#_c_526_n N_VGND_c_1836_n 0.0204687f $X=5.87 $Y=1.395 $X2=0
+ $Y2=0
cc_510 N_A_1124_81#_c_530_n N_VGND_c_1836_n 0.00192581f $X=8.78 $Y=1.11 $X2=0
+ $Y2=0
cc_511 N_A_1124_81#_c_530_n N_A_1454_173#_c_1935_n 0.0193329f $X=8.78 $Y=1.11
+ $X2=0 $Y2=0
cc_512 N_A_1124_81#_c_530_n N_A_1454_173#_c_1937_n 0.0143234f $X=8.78 $Y=1.11
+ $X2=0.24 $Y2=0
cc_513 N_A_1067_107#_c_632_n N_A_1570_457#_M1008_d 6.97726e-19 $X=13.535
+ $Y=3.145 $X2=0 $Y2=0
cc_514 N_A_1067_107#_c_621_n N_A_1570_457#_c_796_n 0.00336688f $X=12.395
+ $Y=3.285 $X2=0 $Y2=0
cc_515 N_A_1067_107#_c_630_n N_A_1570_457#_c_796_n 0.0212392f $X=13.44 $Y=3.37
+ $X2=0 $Y2=0
cc_516 N_A_1067_107#_c_632_n N_A_1570_457#_c_796_n 0.0218542f $X=13.535 $Y=3.145
+ $X2=0 $Y2=0
cc_517 N_A_1067_107#_c_637_n N_A_1570_457#_c_796_n 0.0294443f $X=13.605 $Y=2.35
+ $X2=0 $Y2=0
cc_518 N_A_1067_107#_c_624_n N_A_1570_457#_c_784_n 7.39135e-19 $X=7.39 $Y=1.645
+ $X2=0 $Y2=0
cc_519 N_A_1067_107#_c_624_n N_A_1570_457#_c_785_n 0.0235115f $X=7.39 $Y=1.645
+ $X2=0 $Y2=0
cc_520 N_A_1067_107#_c_632_n N_A_1570_457#_c_798_n 0.00603917f $X=13.535
+ $Y=3.145 $X2=0 $Y2=0
cc_521 N_A_1067_107#_M1001_g N_A_1570_457#_c_799_n 0.0763549f $X=7.39 $Y=3.105
+ $X2=0 $Y2=0
cc_522 N_A_1067_107#_c_632_n N_A_1570_457#_c_800_n 0.0516061f $X=13.535 $Y=3.145
+ $X2=0 $Y2=0
cc_523 N_A_1067_107#_c_632_n N_A_1570_457#_c_801_n 0.0112137f $X=13.535 $Y=3.145
+ $X2=0 $Y2=0
cc_524 N_A_1067_107#_c_621_n N_A_1570_457#_c_786_n 8.31928e-19 $X=12.395
+ $Y=3.285 $X2=0 $Y2=0
cc_525 N_A_1067_107#_c_623_n N_A_1570_457#_c_786_n 0.00948375f $X=12.315
+ $Y=1.075 $X2=0 $Y2=0
cc_526 N_A_1067_107#_c_632_n N_A_1570_457#_c_802_n 0.0210328f $X=13.535 $Y=3.145
+ $X2=0 $Y2=0
cc_527 N_A_1067_107#_c_623_n N_A_1570_457#_c_787_n 0.0157359f $X=12.315 $Y=1.075
+ $X2=0 $Y2=0
cc_528 N_A_1067_107#_c_623_n N_A_1570_457#_c_788_n 0.0232604f $X=12.315 $Y=1.075
+ $X2=0 $Y2=0
cc_529 N_A_1067_107#_c_632_n N_A_1570_457#_c_820_n 0.00422089f $X=13.535
+ $Y=3.145 $X2=0 $Y2=0
cc_530 N_A_1067_107#_c_632_n N_A_1570_457#_c_793_n 0.0135797f $X=13.535 $Y=3.145
+ $X2=0 $Y2=0
cc_531 N_A_1067_107#_c_621_n N_A_1570_457#_c_795_n 5.62589e-19 $X=12.395
+ $Y=3.285 $X2=0 $Y2=0
cc_532 N_A_1067_107#_c_637_n N_A_1570_457#_c_795_n 0.00626464f $X=13.605 $Y=2.35
+ $X2=0 $Y2=0
cc_533 N_A_1067_107#_M1001_g N_A_1570_457#_c_805_n 0.0235115f $X=7.39 $Y=3.105
+ $X2=0 $Y2=0
cc_534 N_A_1067_107#_c_632_n N_A_1570_457#_c_806_n 0.00378428f $X=13.535
+ $Y=3.145 $X2=0 $Y2=0
cc_535 N_A_1067_107#_c_632_n N_A_1726_453#_M1024_s 0.00210346f $X=13.535
+ $Y=3.145 $X2=0 $Y2=0
cc_536 N_A_1067_107#_c_632_n N_A_1726_453#_M1027_g 0.00918884f $X=13.535
+ $Y=3.145 $X2=0 $Y2=0
cc_537 N_A_1067_107#_c_621_n N_A_1726_453#_M1034_g 0.0331583f $X=12.395 $Y=3.285
+ $X2=0 $Y2=0
cc_538 N_A_1067_107#_c_630_n N_A_1726_453#_M1034_g 0.0031855f $X=13.44 $Y=3.37
+ $X2=0 $Y2=0
cc_539 N_A_1067_107#_c_632_n N_A_1726_453#_M1034_g 0.00794742f $X=13.535
+ $Y=3.145 $X2=0 $Y2=0
cc_540 N_A_1067_107#_c_621_n N_A_1726_453#_c_968_n 0.00540301f $X=12.395
+ $Y=3.285 $X2=0 $Y2=0
cc_541 N_A_1067_107#_c_623_n N_A_1726_453#_c_968_n 0.010812f $X=12.315 $Y=1.075
+ $X2=0 $Y2=0
cc_542 N_A_1067_107#_c_621_n N_A_1726_453#_c_999_n 0.0395636f $X=12.395 $Y=3.285
+ $X2=0 $Y2=0
cc_543 N_A_1067_107#_c_621_n N_A_1726_453#_c_976_n 0.0380527f $X=12.395 $Y=3.285
+ $X2=0 $Y2=0
cc_544 N_A_1067_107#_c_623_n N_A_1726_453#_c_976_n 0.00740688f $X=12.315
+ $Y=1.075 $X2=0 $Y2=0
cc_545 N_A_1067_107#_c_632_n N_CLK_c_1076_n 0.00473331f $X=13.535 $Y=3.145 $X2=0
+ $Y2=0
cc_546 N_A_1067_107#_c_623_n N_CLK_M1026_g 0.00110492f $X=12.315 $Y=1.075 $X2=0
+ $Y2=0
cc_547 N_A_1067_107#_c_637_n N_A_2789_147#_c_1122_n 0.00384577f $X=13.605
+ $Y=2.35 $X2=0.24 $Y2=0
cc_548 N_A_1067_107#_c_637_n N_A_2789_147#_c_1127_n 0.00724778f $X=13.605
+ $Y=2.35 $X2=0 $Y2=0
cc_549 N_A_1067_107#_c_637_n N_A_2789_147#_c_1128_n 0.00678093f $X=13.605
+ $Y=2.35 $X2=0 $Y2=0
cc_550 N_A_1067_107#_c_632_n N_A_2518_445#_M1034_d 0.0012879f $X=13.535 $Y=3.145
+ $X2=0 $Y2=0
cc_551 N_A_1067_107#_c_621_n N_A_2518_445#_c_1231_n 0.025095f $X=12.395 $Y=3.285
+ $X2=19.44 $Y2=0
cc_552 N_A_1067_107#_c_637_n N_A_2518_445#_c_1231_n 0.00360947f $X=13.605
+ $Y=2.35 $X2=19.44 $Y2=0
cc_553 N_A_1067_107#_c_621_n N_A_2518_445#_c_1232_n 0.0537025f $X=12.395
+ $Y=3.285 $X2=0 $Y2=0
cc_554 N_A_1067_107#_c_630_n N_A_2518_445#_c_1232_n 0.0191164f $X=13.44 $Y=3.37
+ $X2=0 $Y2=0
cc_555 N_A_1067_107#_c_632_n N_A_2518_445#_c_1232_n 0.0214005f $X=13.535
+ $Y=3.145 $X2=0 $Y2=0
cc_556 N_A_1067_107#_c_634_n N_A_2518_445#_c_1232_n 2.42664e-19 $X=13.68
+ $Y=3.145 $X2=0 $Y2=0
cc_557 N_A_1067_107#_c_637_n N_A_2518_445#_c_1232_n 0.0244604f $X=13.605 $Y=2.35
+ $X2=0 $Y2=0
cc_558 N_A_1067_107#_c_621_n N_A_2518_445#_c_1225_n 0.023895f $X=12.395 $Y=3.285
+ $X2=9.84 $Y2=0
cc_559 N_A_1067_107#_c_637_n N_A_2518_445#_c_1234_n 0.0245542f $X=13.605 $Y=2.35
+ $X2=0 $Y2=0
cc_560 N_A_1067_107#_c_623_n N_A_2518_445#_c_1226_n 0.0218007f $X=12.315
+ $Y=1.075 $X2=0 $Y2=0
cc_561 N_A_1067_107#_c_632_n N_VPWR_M1035_d 0.00956677f $X=13.535 $Y=3.145 $X2=0
+ $Y2=0
cc_562 N_A_1067_107#_c_632_n N_VPWR_M1024_d 6.97726e-19 $X=13.535 $Y=3.145 $X2=0
+ $Y2=0
cc_563 N_A_1067_107#_M1001_g N_VPWR_c_1349_n 0.00169299f $X=7.39 $Y=3.105 $X2=0
+ $Y2=0
cc_564 N_A_1067_107#_c_632_n N_VPWR_c_1349_n 9.45631e-19 $X=13.535 $Y=3.145
+ $X2=0 $Y2=0
cc_565 N_A_1067_107#_c_632_n N_VPWR_c_1352_n 0.0386721f $X=13.535 $Y=3.145 $X2=0
+ $Y2=0
cc_566 N_A_1067_107#_M1035_s N_VPWR_c_1364_n 5.0983e-19 $X=5.58 $Y=2.715 $X2=0
+ $Y2=0
cc_567 N_A_1067_107#_M1001_g N_VPWR_c_1364_n 0.00561012f $X=7.39 $Y=3.105 $X2=0
+ $Y2=0
cc_568 N_A_1067_107#_c_630_n N_VPWR_c_1364_n 0.0323894f $X=13.44 $Y=3.37 $X2=0
+ $Y2=0
cc_569 N_A_1067_107#_c_631_n N_VPWR_c_1364_n 0.00508063f $X=12.48 $Y=3.37 $X2=0
+ $Y2=0
cc_570 N_A_1067_107#_c_632_n N_VPWR_c_1364_n 0.60918f $X=13.535 $Y=3.145 $X2=0
+ $Y2=0
cc_571 N_A_1067_107#_c_633_n N_VPWR_c_1364_n 0.0247788f $X=5.665 $Y=3.145 $X2=0
+ $Y2=0
cc_572 N_A_1067_107#_c_634_n N_VPWR_c_1364_n 0.0246036f $X=13.68 $Y=3.145 $X2=0
+ $Y2=0
cc_573 N_A_1067_107#_c_625_n N_VPWR_c_1364_n 0.0105705f $X=5.705 $Y=2.86 $X2=0
+ $Y2=0
cc_574 N_A_1067_107#_c_625_n N_A_581_659#_c_1512_n 0.0145597f $X=5.705 $Y=2.86
+ $X2=0 $Y2=0
cc_575 N_A_1067_107#_c_633_n N_A_581_659#_c_1513_n 0.00761388f $X=5.665 $Y=3.145
+ $X2=0 $Y2=0
cc_576 N_A_1067_107#_c_625_n N_A_581_659#_c_1513_n 0.0418107f $X=5.705 $Y=2.86
+ $X2=0 $Y2=0
cc_577 N_A_1067_107#_c_632_n N_A_567_107#_M1027_d 0.00220834f $X=13.535 $Y=3.145
+ $X2=0 $Y2=0
cc_578 N_A_1067_107#_c_625_n N_A_567_107#_c_1563_n 0.0105721f $X=5.705 $Y=2.86
+ $X2=19.44 $Y2=0
cc_579 N_A_1067_107#_M1035_s N_A_567_107#_c_1565_n 0.00141003f $X=5.58 $Y=2.715
+ $X2=9.84 $Y2=0.057
cc_580 N_A_1067_107#_c_632_n N_A_567_107#_c_1565_n 0.00164704f $X=13.535
+ $Y=3.145 $X2=9.84 $Y2=0.057
cc_581 N_A_1067_107#_c_633_n N_A_567_107#_c_1565_n 3.87376e-19 $X=5.665 $Y=3.145
+ $X2=9.84 $Y2=0.057
cc_582 N_A_1067_107#_c_625_n N_A_567_107#_c_1565_n 0.0246936f $X=5.705 $Y=2.86
+ $X2=9.84 $Y2=0.057
cc_583 N_A_1067_107#_c_619_n N_A_567_107#_c_1552_n 0.0752607f $X=5.48 $Y=0.7
+ $X2=0 $Y2=0
cc_584 N_A_1067_107#_c_622_n N_A_567_107#_c_1552_n 0.0137864f $X=5.552 $Y=1.69
+ $X2=0 $Y2=0
cc_585 N_A_1067_107#_c_625_n N_A_567_107#_c_1552_n 0.0309611f $X=5.705 $Y=2.86
+ $X2=0 $Y2=0
cc_586 N_A_1067_107#_c_619_n N_A_567_107#_c_1553_n 0.0209781f $X=5.48 $Y=0.7
+ $X2=0 $Y2=0
cc_587 N_A_1067_107#_c_619_n N_A_567_107#_c_1618_n 0.0435526f $X=5.48 $Y=0.7
+ $X2=0 $Y2=0
cc_588 N_A_1067_107#_c_632_n N_A_567_107#_c_1619_n 0.0111301f $X=13.535 $Y=3.145
+ $X2=0 $Y2=0
cc_589 N_A_1067_107#_c_633_n N_A_567_107#_c_1619_n 2.2981e-19 $X=5.665 $Y=3.145
+ $X2=0 $Y2=0
cc_590 N_A_1067_107#_c_625_n N_A_567_107#_c_1619_n 0.0542782f $X=5.705 $Y=2.86
+ $X2=0 $Y2=0
cc_591 N_A_1067_107#_c_625_n N_A_567_107#_c_1621_n 0.00562232f $X=5.705 $Y=2.86
+ $X2=0 $Y2=0
cc_592 N_A_1067_107#_c_618_n N_A_567_107#_c_1557_n 0.0245956f $X=7.02 $Y=1.395
+ $X2=0 $Y2=0
cc_593 N_A_1067_107#_c_620_n N_A_567_107#_c_1557_n 0.0760275f $X=6.955 $Y=1.69
+ $X2=0 $Y2=0
cc_594 N_A_1067_107#_c_624_n N_A_567_107#_c_1557_n 0.0117538f $X=7.39 $Y=1.645
+ $X2=0 $Y2=0
cc_595 N_A_1067_107#_c_619_n N_A_567_107#_c_1624_n 0.0128825f $X=5.48 $Y=0.7
+ $X2=0 $Y2=0
cc_596 N_A_1067_107#_c_620_n N_A_567_107#_c_1624_n 0.0123662f $X=6.955 $Y=1.69
+ $X2=0 $Y2=0
cc_597 N_A_1067_107#_M1001_g N_A_567_107#_c_1572_n 0.0211101f $X=7.39 $Y=3.105
+ $X2=0 $Y2=0
cc_598 N_A_1067_107#_c_620_n N_A_567_107#_c_1572_n 0.0679553f $X=6.955 $Y=1.69
+ $X2=0 $Y2=0
cc_599 N_A_1067_107#_c_624_n N_A_567_107#_c_1572_n 0.0112411f $X=7.39 $Y=1.645
+ $X2=0 $Y2=0
cc_600 N_A_1067_107#_c_620_n N_A_567_107#_c_1628_n 0.0123662f $X=6.955 $Y=1.69
+ $X2=0 $Y2=0
cc_601 N_A_1067_107#_c_625_n N_A_567_107#_c_1628_n 0.0130668f $X=5.705 $Y=2.86
+ $X2=0 $Y2=0
cc_602 N_A_1067_107#_M1001_g N_A_567_107#_c_1629_n 0.0162911f $X=7.39 $Y=3.105
+ $X2=0 $Y2=0
cc_603 N_A_1067_107#_c_632_n N_A_567_107#_c_1629_n 0.0378847f $X=13.535 $Y=3.145
+ $X2=0 $Y2=0
cc_604 N_A_1067_107#_M1001_g N_A_567_107#_c_1664_n 0.00406461f $X=7.39 $Y=3.105
+ $X2=0 $Y2=0
cc_605 N_A_1067_107#_c_620_n N_A_567_107#_c_1664_n 0.0122207f $X=6.955 $Y=1.69
+ $X2=0 $Y2=0
cc_606 N_A_1067_107#_c_624_n N_A_567_107#_c_1664_n 0.0297358f $X=7.39 $Y=1.645
+ $X2=0 $Y2=0
cc_607 N_A_1067_107#_c_624_n N_A_567_107#_c_1558_n 0.0111782f $X=7.39 $Y=1.645
+ $X2=0 $Y2=0
cc_608 N_A_1067_107#_M1001_g N_A_567_107#_c_1573_n 0.00590842f $X=7.39 $Y=3.105
+ $X2=0 $Y2=0
cc_609 N_A_1067_107#_c_632_n N_A_567_107#_c_1573_n 0.0168809f $X=13.535 $Y=3.145
+ $X2=0 $Y2=0
cc_610 N_A_1067_107#_c_632_n N_A_567_107#_c_1634_n 0.00579547f $X=13.535
+ $Y=3.145 $X2=0 $Y2=0
cc_611 N_A_1067_107#_c_633_n N_A_567_107#_c_1634_n 2.61257e-19 $X=5.665 $Y=3.145
+ $X2=0 $Y2=0
cc_612 N_A_1067_107#_c_625_n N_A_567_107#_c_1634_n 0.00736036f $X=5.705 $Y=2.86
+ $X2=0 $Y2=0
cc_613 N_A_1067_107#_c_624_n N_A_567_107#_c_1673_n 0.00339519f $X=7.39 $Y=1.645
+ $X2=0 $Y2=0
cc_614 N_A_1067_107#_M1001_g N_A_567_107#_c_1576_n 0.0205362f $X=7.39 $Y=3.105
+ $X2=0 $Y2=0
cc_615 N_A_1067_107#_c_632_n N_A_567_107#_c_1576_n 0.00912186f $X=13.535
+ $Y=3.145 $X2=0 $Y2=0
cc_616 N_A_1067_107#_c_618_n N_A_567_107#_c_1561_n 0.00374869f $X=7.02 $Y=1.395
+ $X2=0 $Y2=0
cc_617 N_A_1067_107#_c_632_n N_A_567_107#_c_1579_n 0.0175368f $X=13.535 $Y=3.145
+ $X2=0 $Y2=0
cc_618 N_A_1067_107#_c_632_n A_1528_579# 0.00220483f $X=13.535 $Y=3.145 $X2=0
+ $Y2=0
cc_619 N_A_1067_107#_c_621_n N_A_2365_445#_c_1742_n 0.0717884f $X=12.395
+ $Y=3.285 $X2=0 $Y2=0
cc_620 N_A_1067_107#_c_631_n N_A_2365_445#_c_1742_n 0.013485f $X=12.48 $Y=3.37
+ $X2=0 $Y2=0
cc_621 N_A_1067_107#_c_632_n N_A_2365_445#_c_1742_n 0.0324006f $X=13.535
+ $Y=3.145 $X2=0 $Y2=0
cc_622 N_A_1067_107#_c_630_n N_A_2365_445#_c_1743_n 0.0882194f $X=13.44 $Y=3.37
+ $X2=0.24 $Y2=0
cc_623 N_A_1067_107#_c_631_n N_A_2365_445#_c_1743_n 0.0116447f $X=12.48 $Y=3.37
+ $X2=0.24 $Y2=0
cc_624 N_A_1067_107#_c_632_n N_A_2365_445#_c_1743_n 0.00140155f $X=13.535
+ $Y=3.145 $X2=0.24 $Y2=0
cc_625 N_A_1067_107#_c_634_n N_A_2365_445#_c_1743_n 3.17804e-19 $X=13.68
+ $Y=3.145 $X2=0.24 $Y2=0
cc_626 N_A_1067_107#_c_630_n N_A_2365_445#_c_1749_n 0.0125778f $X=13.44 $Y=3.37
+ $X2=0 $Y2=0
cc_627 N_A_1067_107#_c_634_n N_A_2365_445#_c_1749_n 0.00738404f $X=13.68
+ $Y=3.145 $X2=0 $Y2=0
cc_628 N_A_1067_107#_c_637_n N_A_2365_445#_c_1749_n 0.0381323f $X=13.605 $Y=2.35
+ $X2=0 $Y2=0
cc_629 N_A_1067_107#_c_618_n N_VGND_c_1826_n 0.0317577f $X=7.02 $Y=1.395 $X2=0
+ $Y2=0
cc_630 N_A_1067_107#_c_618_n N_VGND_c_1836_n 0.00594485f $X=7.02 $Y=1.395 $X2=0
+ $Y2=0
cc_631 N_A_1067_107#_c_619_n N_VGND_c_1836_n 0.0227758f $X=5.48 $Y=0.7 $X2=0
+ $Y2=0
cc_632 N_A_1067_107#_c_623_n N_VGND_c_1836_n 0.00254021f $X=12.315 $Y=1.075
+ $X2=0 $Y2=0
cc_633 N_A_1067_107#_c_624_n N_A_1454_173#_c_1935_n 2.80466e-19 $X=7.39 $Y=1.645
+ $X2=0 $Y2=0
cc_634 N_A_1067_107#_c_618_n N_A_1454_173#_c_1938_n 0.00903914f $X=7.02 $Y=1.395
+ $X2=0 $Y2=0
cc_635 N_A_1067_107#_c_624_n N_A_1454_173#_c_1938_n 0.00154549f $X=7.39 $Y=1.645
+ $X2=0 $Y2=0
cc_636 N_A_1570_457#_c_800_n N_A_1726_453#_M1024_s 0.00571434f $X=10.185
+ $Y=2.835 $X2=0 $Y2=0
cc_637 N_A_1570_457#_c_799_n N_A_1726_453#_M1027_g 0.0191251f $X=8.255 $Y=2.57
+ $X2=0 $Y2=0
cc_638 N_A_1570_457#_c_800_n N_A_1726_453#_M1027_g 0.00860407f $X=10.185
+ $Y=2.835 $X2=0 $Y2=0
cc_639 N_A_1570_457#_c_820_n N_A_1726_453#_M1027_g 0.00860546f $X=8.92 $Y=2.58
+ $X2=0 $Y2=0
cc_640 N_A_1570_457#_c_806_n N_A_1726_453#_M1027_g 0.0172753f $X=8.135 $Y=2.785
+ $X2=0 $Y2=0
cc_641 N_A_1570_457#_c_796_n N_A_1726_453#_M1034_g 0.010922f $X=13.215 $Y=2.115
+ $X2=0 $Y2=0
cc_642 N_A_1570_457#_c_802_n N_A_1726_453#_M1034_g 7.96352e-19 $X=11.4 $Y=2.485
+ $X2=0 $Y2=0
cc_643 N_A_1570_457#_c_783_n N_A_1726_453#_c_968_n 0.0131639f $X=13.485 $Y=1.395
+ $X2=0 $Y2=0
cc_644 N_A_1570_457#_c_787_n N_A_1726_453#_c_968_n 0.00300768f $X=11.71 $Y=0.745
+ $X2=0 $Y2=0
cc_645 N_A_1570_457#_c_788_n N_A_1726_453#_c_968_n 0.0200643f $X=13.44 $Y=0.56
+ $X2=0 $Y2=0
cc_646 N_A_1570_457#_c_792_n N_A_1726_453#_c_968_n 7.62905e-19 $X=13.525
+ $Y=1.505 $X2=0 $Y2=0
cc_647 N_A_1570_457#_c_785_n N_A_1726_453#_c_980_n 3.61945e-19 $X=8.28 $Y=1.93
+ $X2=0 $Y2=0
cc_648 N_A_1570_457#_c_798_n N_A_1726_453#_c_980_n 0.0157738f $X=8.835 $Y=2.58
+ $X2=0 $Y2=0
cc_649 N_A_1570_457#_c_800_n N_A_1726_453#_c_980_n 0.0182245f $X=10.185 $Y=2.835
+ $X2=0 $Y2=0
cc_650 N_A_1570_457#_c_820_n N_A_1726_453#_c_980_n 0.0238277f $X=8.92 $Y=2.58
+ $X2=0 $Y2=0
cc_651 N_A_1570_457#_c_793_n N_A_1726_453#_c_980_n 0.0132648f $X=10.19 $Y=2.015
+ $X2=0 $Y2=0
cc_652 N_A_1570_457#_c_805_n N_A_1726_453#_c_980_n 0.0191251f $X=8.135 $Y=2.285
+ $X2=0 $Y2=0
cc_653 N_A_1570_457#_c_781_n N_A_1726_453#_c_970_n 0.0169725f $X=10.54 $Y=1.065
+ $X2=0 $Y2=0
cc_654 N_A_1570_457#_c_794_n N_A_1726_453#_c_970_n 0.041671f $X=10.66 $Y=1.25
+ $X2=0 $Y2=0
cc_655 N_A_1570_457#_c_868_p N_A_1726_453#_c_970_n 0.0200141f $X=10.825 $Y=1.23
+ $X2=0 $Y2=0
cc_656 N_A_1570_457#_c_801_n N_A_1726_453#_c_972_n 0.0149686f $X=11.315 $Y=2.385
+ $X2=0 $Y2=0
cc_657 N_A_1570_457#_c_786_n N_A_1726_453#_c_972_n 0.0489463f $X=11.625 $Y=1.18
+ $X2=0 $Y2=0
cc_658 N_A_1570_457#_c_793_n N_A_1726_453#_c_972_n 0.0170339f $X=10.19 $Y=2.015
+ $X2=0 $Y2=0
cc_659 N_A_1570_457#_c_794_n N_A_1726_453#_c_972_n 0.010069f $X=10.66 $Y=1.25
+ $X2=0 $Y2=0
cc_660 N_A_1570_457#_c_868_p N_A_1726_453#_c_972_n 0.0233935f $X=10.825 $Y=1.23
+ $X2=0 $Y2=0
cc_661 N_A_1570_457#_c_793_n N_A_1726_453#_c_973_n 0.015443f $X=10.19 $Y=2.015
+ $X2=0 $Y2=0
cc_662 N_A_1570_457#_c_875_p N_A_1726_453#_c_973_n 0.0219502f $X=10.27 $Y=2.017
+ $X2=0 $Y2=0
cc_663 N_A_1570_457#_c_800_n N_A_1726_453#_c_987_n 0.00972495f $X=10.185
+ $Y=2.835 $X2=0 $Y2=0
cc_664 N_A_1570_457#_c_800_n N_A_1726_453#_c_981_n 0.0196118f $X=10.185 $Y=2.835
+ $X2=0 $Y2=0
cc_665 N_A_1570_457#_c_878_p N_A_1726_453#_c_981_n 0.00678895f $X=10.27 $Y=2.75
+ $X2=0 $Y2=0
cc_666 N_A_1570_457#_c_820_n N_A_1726_453#_c_981_n 0.00225693f $X=8.92 $Y=2.58
+ $X2=0 $Y2=0
cc_667 N_A_1570_457#_c_793_n N_A_1726_453#_c_981_n 0.00541352f $X=10.19 $Y=2.015
+ $X2=0 $Y2=0
cc_668 N_A_1570_457#_c_881_p N_A_1726_453#_c_981_n 0.0114341f $X=10.27 $Y=2.385
+ $X2=0 $Y2=0
cc_669 N_A_1570_457#_c_882_p N_A_1726_453#_c_974_n 0.00680987f $X=10.27 $Y=2.3
+ $X2=0 $Y2=0
cc_670 N_A_1570_457#_c_793_n N_A_1726_453#_c_974_n 0.00977826f $X=10.19 $Y=2.015
+ $X2=0 $Y2=0
cc_671 N_A_1570_457#_c_875_p N_A_1726_453#_c_974_n 0.0175736f $X=10.27 $Y=2.017
+ $X2=0 $Y2=0
cc_672 N_A_1570_457#_c_881_p N_A_1726_453#_c_974_n 9.24685e-19 $X=10.27 $Y=2.385
+ $X2=0 $Y2=0
cc_673 N_A_1570_457#_c_786_n N_A_1726_453#_c_999_n 0.00624485f $X=11.625 $Y=1.18
+ $X2=0 $Y2=0
cc_674 N_A_1570_457#_c_784_n N_A_1726_453#_M1030_g 0.0365593f $X=8.28 $Y=1.43
+ $X2=0 $Y2=0
cc_675 N_A_1570_457#_c_794_n N_A_1726_453#_M1030_g 0.0132648f $X=10.66 $Y=1.25
+ $X2=0 $Y2=0
cc_676 N_A_1570_457#_c_805_n N_A_1726_453#_M1030_g 0.00608726f $X=8.135 $Y=2.285
+ $X2=0 $Y2=0
cc_677 N_A_1570_457#_c_786_n N_A_1726_453#_c_976_n 0.00277034f $X=11.625 $Y=1.18
+ $X2=0 $Y2=0
cc_678 N_A_1570_457#_c_795_n N_A_1726_453#_c_976_n 0.027942f $X=13.445 $Y=1.62
+ $X2=0 $Y2=0
cc_679 N_A_1570_457#_c_878_p N_CLK_c_1076_n 0.00105601f $X=10.27 $Y=2.75 $X2=0
+ $Y2=0
cc_680 N_A_1570_457#_c_801_n N_CLK_c_1076_n 0.0260888f $X=11.315 $Y=2.385 $X2=0
+ $Y2=0
cc_681 N_A_1570_457#_c_802_n N_CLK_c_1076_n 0.00222082f $X=11.4 $Y=2.485 $X2=0
+ $Y2=0
cc_682 N_A_1570_457#_c_882_p N_CLK_c_1073_n 9.13397e-19 $X=10.27 $Y=2.3 $X2=0
+ $Y2=0
cc_683 N_A_1570_457#_c_801_n N_CLK_c_1073_n 0.0105309f $X=11.315 $Y=2.385 $X2=0
+ $Y2=0
cc_684 N_A_1570_457#_c_793_n N_CLK_c_1073_n 0.0550573f $X=10.19 $Y=2.015 $X2=0
+ $Y2=0
cc_685 N_A_1570_457#_c_875_p N_CLK_c_1073_n 3.2947e-19 $X=10.27 $Y=2.017 $X2=0
+ $Y2=0
cc_686 N_A_1570_457#_c_794_n N_CLK_c_1073_n 0.00548119f $X=10.66 $Y=1.25 $X2=0
+ $Y2=0
cc_687 N_A_1570_457#_c_781_n N_CLK_M1026_g 0.0141968f $X=10.54 $Y=1.065 $X2=0
+ $Y2=0
cc_688 N_A_1570_457#_c_786_n N_CLK_M1026_g 0.0298245f $X=11.625 $Y=1.18 $X2=0
+ $Y2=0
cc_689 N_A_1570_457#_c_787_n N_CLK_M1026_g 0.0068721f $X=11.71 $Y=0.745 $X2=0
+ $Y2=0
cc_690 N_A_1570_457#_c_790_n N_CLK_M1026_g 0.00174579f $X=11.875 $Y=0.56 $X2=0
+ $Y2=0
cc_691 N_A_1570_457#_c_793_n N_CLK_M1026_g 0.00364643f $X=10.19 $Y=2.015 $X2=0
+ $Y2=0
cc_692 N_A_1570_457#_c_794_n N_CLK_M1026_g 0.033206f $X=10.66 $Y=1.25 $X2=0
+ $Y2=0
cc_693 N_A_1570_457#_c_868_p N_CLK_M1026_g 6.95325e-19 $X=10.825 $Y=1.23 $X2=0
+ $Y2=0
cc_694 N_A_1570_457#_c_801_n CLK 0.0487346f $X=11.315 $Y=2.385 $X2=0 $Y2=0
cc_695 N_A_1570_457#_c_793_n CLK 0.00206799f $X=10.19 $Y=2.015 $X2=0 $Y2=0
cc_696 N_A_1570_457#_c_875_p CLK 0.0115512f $X=10.27 $Y=2.017 $X2=0 $Y2=0
cc_697 N_A_1570_457#_c_783_n N_A_2789_147#_M1031_g 0.0812419f $X=13.485 $Y=1.395
+ $X2=0 $Y2=0
cc_698 N_A_1570_457#_c_792_n N_A_2789_147#_M1031_g 0.0016121f $X=13.525 $Y=1.505
+ $X2=0 $Y2=0
cc_699 N_A_1570_457#_c_795_n N_A_2789_147#_M1031_g 0.0124361f $X=13.445 $Y=1.62
+ $X2=0 $Y2=0
cc_700 N_A_1570_457#_c_913_p N_A_2789_147#_M1031_g 0.00128146f $X=13.525 $Y=1.62
+ $X2=0 $Y2=0
cc_701 N_A_1570_457#_c_796_n N_A_2789_147#_c_1128_n 0.00841341f $X=13.215
+ $Y=2.115 $X2=0 $Y2=0
cc_702 N_A_1570_457#_c_796_n N_A_2518_445#_c_1231_n 0.0105713f $X=13.215
+ $Y=2.115 $X2=19.44 $Y2=0
cc_703 N_A_1570_457#_c_795_n N_A_2518_445#_c_1231_n 0.00366213f $X=13.445
+ $Y=1.62 $X2=19.44 $Y2=0
cc_704 N_A_1570_457#_c_796_n N_A_2518_445#_c_1232_n 0.0228702f $X=13.215
+ $Y=2.115 $X2=0 $Y2=0
cc_705 N_A_1570_457#_c_783_n N_A_2518_445#_c_1225_n 5.7835e-19 $X=13.485
+ $Y=1.395 $X2=9.84 $Y2=0
cc_706 N_A_1570_457#_c_792_n N_A_2518_445#_c_1225_n 0.00619986f $X=13.525
+ $Y=1.505 $X2=9.84 $Y2=0
cc_707 N_A_1570_457#_c_795_n N_A_2518_445#_c_1225_n 0.0095851f $X=13.445 $Y=1.62
+ $X2=9.84 $Y2=0
cc_708 N_A_1570_457#_c_913_p N_A_2518_445#_c_1225_n 0.0115348f $X=13.525 $Y=1.62
+ $X2=9.84 $Y2=0
cc_709 N_A_1570_457#_c_795_n N_A_2518_445#_c_1234_n 0.0508801f $X=13.445 $Y=1.62
+ $X2=0 $Y2=0
cc_710 N_A_1570_457#_c_913_p N_A_2518_445#_c_1234_n 0.0218397f $X=13.525 $Y=1.62
+ $X2=0 $Y2=0
cc_711 N_A_1570_457#_c_783_n N_A_2518_445#_c_1226_n 0.0103904f $X=13.485
+ $Y=1.395 $X2=0 $Y2=0
cc_712 N_A_1570_457#_c_788_n N_A_2518_445#_c_1226_n 0.0304175f $X=13.44 $Y=0.56
+ $X2=0 $Y2=0
cc_713 N_A_1570_457#_c_792_n N_A_2518_445#_c_1226_n 0.0349418f $X=13.525
+ $Y=1.505 $X2=0 $Y2=0
cc_714 N_A_1570_457#_c_795_n N_A_2518_445#_c_1226_n 0.00584656f $X=13.445
+ $Y=1.62 $X2=0 $Y2=0
cc_715 N_A_1570_457#_c_801_n N_VPWR_M1024_d 0.00178343f $X=11.315 $Y=2.385 $X2=0
+ $Y2=0
cc_716 N_A_1570_457#_c_801_n N_VPWR_c_1352_n 0.0384364f $X=11.315 $Y=2.385 $X2=0
+ $Y2=0
cc_717 N_A_1570_457#_c_802_n N_VPWR_c_1352_n 0.01782f $X=11.4 $Y=2.485 $X2=0
+ $Y2=0
cc_718 N_A_1570_457#_c_793_n N_VPWR_c_1352_n 0.00352629f $X=10.19 $Y=2.015 $X2=0
+ $Y2=0
cc_719 N_A_1570_457#_c_802_n N_VPWR_c_1364_n 0.00150701f $X=11.4 $Y=2.485 $X2=0
+ $Y2=0
cc_720 N_A_1570_457#_c_793_n N_VPWR_c_1364_n 0.0094923f $X=10.19 $Y=2.015 $X2=0
+ $Y2=0
cc_721 N_A_1570_457#_c_800_n N_A_567_107#_M1027_d 0.00224f $X=10.185 $Y=2.835
+ $X2=0 $Y2=0
cc_722 N_A_1570_457#_c_805_n N_A_567_107#_c_1572_n 8.64057e-19 $X=8.135 $Y=2.285
+ $X2=0 $Y2=0
cc_723 N_A_1570_457#_c_785_n N_A_567_107#_c_1664_n 0.00281759f $X=8.28 $Y=1.93
+ $X2=0 $Y2=0
cc_724 N_A_1570_457#_c_784_n N_A_567_107#_c_1558_n 3.30196e-19 $X=8.28 $Y=1.43
+ $X2=0 $Y2=0
cc_725 N_A_1570_457#_c_798_n N_A_567_107#_c_1573_n 0.00176082f $X=8.835 $Y=2.58
+ $X2=0 $Y2=0
cc_726 N_A_1570_457#_c_800_n N_A_567_107#_c_1573_n 0.00191701f $X=10.185
+ $Y=2.835 $X2=0 $Y2=0
cc_727 N_A_1570_457#_c_820_n N_A_567_107#_c_1573_n 0.00349056f $X=8.92 $Y=2.58
+ $X2=0 $Y2=0
cc_728 N_A_1570_457#_c_806_n N_A_567_107#_c_1573_n 0.0244699f $X=8.135 $Y=2.785
+ $X2=0 $Y2=0
cc_729 N_A_1570_457#_c_806_n N_A_567_107#_c_1576_n 0.00141958f $X=8.135 $Y=2.785
+ $X2=0 $Y2=0
cc_730 N_A_1570_457#_c_784_n N_A_567_107#_c_1561_n 0.016403f $X=8.28 $Y=1.43
+ $X2=0 $Y2=0
cc_731 N_A_1570_457#_c_785_n N_A_567_107#_c_1561_n 0.0122033f $X=8.28 $Y=1.93
+ $X2=0 $Y2=0
cc_732 N_A_1570_457#_c_800_n N_A_567_107#_c_1579_n 0.0173768f $X=10.185 $Y=2.835
+ $X2=0 $Y2=0
cc_733 N_A_1570_457#_c_793_n N_A_567_107#_c_1579_n 0.00195f $X=10.19 $Y=2.015
+ $X2=0 $Y2=0
cc_734 N_A_1570_457#_c_801_n N_A_2365_445#_c_1742_n 0.0125436f $X=11.315
+ $Y=2.385 $X2=0 $Y2=0
cc_735 N_A_1570_457#_c_802_n N_A_2365_445#_c_1742_n 0.0431128f $X=11.4 $Y=2.485
+ $X2=0 $Y2=0
cc_736 N_A_1570_457#_c_796_n N_A_2365_445#_c_1743_n 0.00244394f $X=13.215
+ $Y=2.115 $X2=0.24 $Y2=0
cc_737 N_A_1570_457#_c_796_n N_A_2365_445#_c_1749_n 0.00134212f $X=13.215
+ $Y=2.115 $X2=0 $Y2=0
cc_738 N_A_1570_457#_c_781_n N_VGND_c_1828_n 0.0317136f $X=10.54 $Y=1.065 $X2=0
+ $Y2=0
cc_739 N_A_1570_457#_c_790_n N_VGND_c_1828_n 0.00911032f $X=11.875 $Y=0.56 $X2=0
+ $Y2=0
cc_740 N_A_1570_457#_c_868_p N_VGND_c_1828_n 0.0623901f $X=10.825 $Y=1.23 $X2=0
+ $Y2=0
cc_741 N_A_1570_457#_c_783_n N_VGND_c_1830_n 0.00281258f $X=13.485 $Y=1.395
+ $X2=0 $Y2=0
cc_742 N_A_1570_457#_c_788_n N_VGND_c_1830_n 0.00747629f $X=13.44 $Y=0.56 $X2=0
+ $Y2=0
cc_743 N_A_1570_457#_c_792_n N_VGND_c_1830_n 0.0227465f $X=13.525 $Y=1.505 $X2=0
+ $Y2=0
cc_744 N_A_1570_457#_M1026_d N_VGND_c_1836_n 6.6074e-19 $X=11.57 $Y=0.535 $X2=0
+ $Y2=0
cc_745 N_A_1570_457#_c_781_n N_VGND_c_1836_n 0.0118525f $X=10.54 $Y=1.065 $X2=0
+ $Y2=0
cc_746 N_A_1570_457#_c_783_n N_VGND_c_1836_n 0.00411901f $X=13.485 $Y=1.395
+ $X2=0 $Y2=0
cc_747 N_A_1570_457#_c_786_n N_VGND_c_1836_n 0.00579828f $X=11.625 $Y=1.18 $X2=0
+ $Y2=0
cc_748 N_A_1570_457#_c_788_n N_VGND_c_1836_n 0.0942134f $X=13.44 $Y=0.56 $X2=0
+ $Y2=0
cc_749 N_A_1570_457#_c_790_n N_VGND_c_1836_n 0.0238047f $X=11.875 $Y=0.56 $X2=0
+ $Y2=0
cc_750 N_A_1570_457#_c_868_p N_VGND_c_1836_n 0.00360995f $X=10.825 $Y=1.23 $X2=0
+ $Y2=0
cc_751 N_A_1570_457#_c_784_n N_A_1454_173#_c_1935_n 0.0238873f $X=8.28 $Y=1.43
+ $X2=0 $Y2=0
cc_752 N_A_1570_457#_c_781_n N_A_1454_173#_c_1937_n 8.1256e-19 $X=10.54 $Y=1.065
+ $X2=0.24 $Y2=0
cc_753 N_A_1570_457#_c_794_n N_A_1454_173#_c_1937_n 0.0031168f $X=10.66 $Y=1.25
+ $X2=0.24 $Y2=0
cc_754 N_A_1570_457#_c_784_n N_A_1454_173#_c_1938_n 0.00441215f $X=8.28 $Y=1.43
+ $X2=0 $Y2=0
cc_755 N_A_1726_453#_M1034_g N_CLK_c_1073_n 0.00423485f $X=12.34 $Y=2.435 $X2=0
+ $Y2=0
cc_756 N_A_1726_453#_c_972_n N_CLK_c_1073_n 0.00761182f $X=11.8 $Y=1.63 $X2=0
+ $Y2=0
cc_757 N_A_1726_453#_c_972_n N_CLK_M1026_g 0.0306302f $X=11.8 $Y=1.63 $X2=0
+ $Y2=0
cc_758 N_A_1726_453#_c_999_n N_CLK_M1026_g 0.0026884f $X=11.965 $Y=1.56 $X2=0
+ $Y2=0
cc_759 N_A_1726_453#_c_976_n N_CLK_M1026_g 0.05099f $X=12.34 $Y=1.745 $X2=0
+ $Y2=0
cc_760 N_A_1726_453#_c_972_n CLK 0.0487261f $X=11.8 $Y=1.63 $X2=0 $Y2=0
cc_761 N_A_1726_453#_c_999_n CLK 0.00511755f $X=11.965 $Y=1.56 $X2=0 $Y2=0
cc_762 N_A_1726_453#_c_976_n CLK 7.66893e-19 $X=12.34 $Y=1.745 $X2=0 $Y2=0
cc_763 N_A_1726_453#_M1034_g N_A_2518_445#_c_1231_n 0.00168742f $X=12.34
+ $Y=2.435 $X2=19.44 $Y2=0
cc_764 N_A_1726_453#_c_976_n N_A_2518_445#_c_1231_n 0.00803058f $X=12.34
+ $Y=1.745 $X2=19.44 $Y2=0
cc_765 N_A_1726_453#_M1034_g N_A_2518_445#_c_1232_n 0.00413505f $X=12.34
+ $Y=2.435 $X2=0 $Y2=0
cc_766 N_A_1726_453#_c_968_n N_A_2518_445#_c_1225_n 0.00335489f $X=12.705
+ $Y=1.395 $X2=9.84 $Y2=0
cc_767 N_A_1726_453#_c_976_n N_A_2518_445#_c_1225_n 0.0154468f $X=12.34 $Y=1.745
+ $X2=9.84 $Y2=0
cc_768 N_A_1726_453#_c_968_n N_A_2518_445#_c_1226_n 0.0193819f $X=12.705
+ $Y=1.395 $X2=0 $Y2=0
cc_769 N_A_1726_453#_M1027_g N_A_567_107#_c_1573_n 0.0258356f $X=8.88 $Y=3.105
+ $X2=0 $Y2=0
cc_770 N_A_1726_453#_M1027_g N_A_567_107#_c_1579_n 0.0100958f $X=8.88 $Y=3.105
+ $X2=0 $Y2=0
cc_771 N_A_1726_453#_c_980_n N_A_567_107#_c_1579_n 0.00123276f $X=9.17 $Y=2.515
+ $X2=0 $Y2=0
cc_772 N_A_1726_453#_M1034_g N_A_2365_445#_c_1742_n 0.0143391f $X=12.34 $Y=2.435
+ $X2=0 $Y2=0
cc_773 N_A_1726_453#_c_972_n N_A_2365_445#_c_1742_n 5.11203e-19 $X=11.8 $Y=1.63
+ $X2=0 $Y2=0
cc_774 N_A_1726_453#_c_999_n N_A_2365_445#_c_1742_n 0.0263043f $X=11.965 $Y=1.56
+ $X2=0 $Y2=0
cc_775 N_A_1726_453#_c_976_n N_A_2365_445#_c_1742_n 0.00899001f $X=12.34
+ $Y=1.745 $X2=0 $Y2=0
cc_776 N_A_1726_453#_c_970_n N_VGND_c_1828_n 0.0299917f $X=10.15 $Y=0.745 $X2=0
+ $Y2=0
cc_777 N_A_1726_453#_c_970_n N_VGND_c_1836_n 0.0253282f $X=10.15 $Y=0.745 $X2=0
+ $Y2=0
cc_778 N_A_1726_453#_c_970_n N_A_1454_173#_c_1935_n 0.0105605f $X=10.15 $Y=0.745
+ $X2=0 $Y2=0
cc_779 N_A_1726_453#_M1030_g N_A_1454_173#_c_1935_n 0.0230492f $X=9.17 $Y=1.11
+ $X2=0 $Y2=0
cc_780 N_A_1726_453#_c_969_n N_A_1454_173#_c_1937_n 0.0255389f $X=9.675 $Y=1.63
+ $X2=0.24 $Y2=0
cc_781 N_A_1726_453#_c_970_n N_A_1454_173#_c_1937_n 0.0358803f $X=10.15 $Y=0.745
+ $X2=0.24 $Y2=0
cc_782 N_A_1726_453#_M1030_g N_A_1454_173#_c_1937_n 0.0235368f $X=9.17 $Y=1.11
+ $X2=0.24 $Y2=0
cc_783 N_CLK_c_1076_n N_VPWR_c_1352_n 0.0402935f $X=11.01 $Y=2.23 $X2=0 $Y2=0
cc_784 N_CLK_c_1076_n N_VPWR_c_1364_n 0.00258191f $X=11.01 $Y=2.23 $X2=0 $Y2=0
cc_785 N_CLK_c_1076_n N_A_2365_445#_c_1742_n 0.00472104f $X=11.01 $Y=2.23 $X2=0
+ $Y2=0
cc_786 N_CLK_c_1073_n N_A_2365_445#_c_1742_n 6.67653e-19 $X=11.32 $Y=1.755 $X2=0
+ $Y2=0
cc_787 N_CLK_M1026_g N_VGND_c_1828_n 0.0353098f $X=11.32 $Y=0.745 $X2=0 $Y2=0
cc_788 N_CLK_M1026_g N_VGND_c_1836_n 0.00548949f $X=11.32 $Y=0.745 $X2=0 $Y2=0
cc_789 N_A_2789_147#_M1031_g N_A_2518_445#_c_1223_n 0.0136601f $X=14.195
+ $Y=1.075 $X2=0 $Y2=0
cc_790 N_A_2789_147#_c_1118_n N_A_2518_445#_c_1223_n 0.0302658f $X=15.48 $Y=0.66
+ $X2=0 $Y2=0
cc_791 N_A_2789_147#_c_1127_n N_A_2518_445#_M1015_g 0.0141029f $X=15.315 $Y=2.39
+ $X2=0 $Y2=0
cc_792 N_A_2789_147#_c_1128_n N_A_2518_445#_M1015_g 0.031999f $X=14.63 $Y=2.39
+ $X2=0 $Y2=0
cc_793 N_A_2789_147#_c_1118_n N_A_2518_445#_M1015_g 0.0240848f $X=15.48 $Y=0.66
+ $X2=0 $Y2=0
cc_794 N_A_2789_147#_c_1130_n N_A_2518_445#_M1015_g 0.0154155f $X=15.83 $Y=3.57
+ $X2=0 $Y2=0
cc_795 N_A_2789_147#_c_1134_n N_A_2518_445#_M1015_g 0.00609808f $X=15.995
+ $Y=3.72 $X2=0 $Y2=0
cc_796 N_A_2789_147#_c_1137_n N_A_2518_445#_M1015_g 0.0237887f $X=15.545 $Y=2.39
+ $X2=0 $Y2=0
cc_797 N_A_2789_147#_c_1138_n N_A_2518_445#_M1015_g 0.00475975f $X=15.83 $Y=2.86
+ $X2=0 $Y2=0
cc_798 N_A_2789_147#_c_1139_n N_A_2518_445#_M1015_g 0.0115472f $X=15.8 $Y=2.695
+ $X2=0 $Y2=0
cc_799 N_A_2789_147#_c_1120_n N_A_2518_445#_M1015_g 0.00396436f $X=17.645
+ $Y=1.665 $X2=0 $Y2=0
cc_800 N_A_2789_147#_M1031_g N_A_2518_445#_c_1234_n 0.042931f $X=14.195 $Y=1.075
+ $X2=0 $Y2=0
cc_801 N_A_2789_147#_c_1127_n N_A_2518_445#_c_1234_n 0.0508731f $X=15.315
+ $Y=2.39 $X2=0 $Y2=0
cc_802 N_A_2789_147#_c_1128_n N_A_2518_445#_c_1234_n 0.0113513f $X=14.63 $Y=2.39
+ $X2=0 $Y2=0
cc_803 N_A_2789_147#_c_1118_n N_A_2518_445#_c_1234_n 0.0140491f $X=15.48 $Y=0.66
+ $X2=0 $Y2=0
cc_804 N_A_2789_147#_M1031_g N_A_2518_445#_c_1235_n 0.00300205f $X=14.195
+ $Y=1.075 $X2=0 $Y2=0
cc_805 N_A_2789_147#_c_1118_n N_A_2518_445#_c_1235_n 0.0272184f $X=15.48 $Y=0.66
+ $X2=0 $Y2=0
cc_806 N_A_2789_147#_M1031_g N_A_2518_445#_c_1227_n 0.0237094f $X=14.195
+ $Y=1.075 $X2=0 $Y2=0
cc_807 N_A_2789_147#_M1010_g N_A_2518_445#_c_1227_n 0.00396436f $X=16.51 $Y=0.91
+ $X2=0 $Y2=0
cc_808 N_A_2789_147#_c_1127_n N_A_2518_445#_c_1227_n 0.0034152f $X=15.315
+ $Y=2.39 $X2=0 $Y2=0
cc_809 N_A_2789_147#_c_1128_n N_A_2518_445#_c_1227_n 0.00193533f $X=14.63
+ $Y=2.39 $X2=0 $Y2=0
cc_810 N_A_2789_147#_c_1118_n N_A_2518_445#_c_1227_n 0.0439895f $X=15.48 $Y=0.66
+ $X2=0 $Y2=0
cc_811 N_A_2789_147#_M1032_g N_A_3531_107#_c_1305_n 0.0292934f $X=17.405
+ $Y=0.745 $X2=19.44 $Y2=0
cc_812 N_A_2789_147#_c_1120_n N_A_3531_107#_c_1305_n 0.0138642f $X=17.645
+ $Y=1.665 $X2=19.44 $Y2=0
cc_813 N_A_2789_147#_M1033_g N_A_3531_107#_c_1313_n 0.0176886f $X=17.645 $Y=2.42
+ $X2=9.84 $Y2=0
cc_814 N_A_2789_147#_c_1174_p N_A_3531_107#_c_1307_n 0.0049561f $X=16.89 $Y=1.67
+ $X2=0 $Y2=0
cc_815 N_A_2789_147#_c_1120_n N_A_3531_107#_c_1307_n 0.0333031f $X=17.645
+ $Y=1.665 $X2=0 $Y2=0
cc_816 N_A_2789_147#_c_1120_n N_A_3531_107#_c_1317_n 0.00791153f $X=17.645
+ $Y=1.665 $X2=0 $Y2=0
cc_817 N_A_2789_147#_c_1122_n N_VPWR_c_1355_n 0.0437496f $X=14.565 $Y=2.605
+ $X2=0 $Y2=0
cc_818 N_A_2789_147#_c_1127_n N_VPWR_c_1355_n 0.062512f $X=15.315 $Y=2.39 $X2=0
+ $Y2=0
cc_819 N_A_2789_147#_c_1134_n N_VPWR_c_1355_n 0.00619827f $X=15.995 $Y=3.72
+ $X2=0 $Y2=0
cc_820 N_A_2789_147#_c_1137_n N_VPWR_c_1355_n 0.00876829f $X=15.545 $Y=2.39
+ $X2=0 $Y2=0
cc_821 N_A_2789_147#_c_1138_n N_VPWR_c_1355_n 0.0692219f $X=15.83 $Y=2.86 $X2=0
+ $Y2=0
cc_822 N_A_2789_147#_M1009_g N_VPWR_c_1358_n 0.00368676f $X=16.77 $Y=2.795 $X2=0
+ $Y2=0
cc_823 N_A_2789_147#_M1033_g N_VPWR_c_1358_n 0.071536f $X=17.645 $Y=2.42 $X2=0
+ $Y2=0
cc_824 N_A_2789_147#_c_1131_n N_VPWR_c_1358_n 0.00472818f $X=16.725 $Y=3.72
+ $X2=0 $Y2=0
cc_825 N_A_2789_147#_c_1185_p N_VPWR_c_1358_n 0.0573846f $X=16.81 $Y=3.635 $X2=0
+ $Y2=0
cc_826 N_A_2789_147#_c_1120_n N_VPWR_c_1358_n 0.0100705f $X=17.645 $Y=1.665
+ $X2=0 $Y2=0
cc_827 N_A_2789_147#_M1033_g N_VPWR_c_1361_n 0.00488892f $X=17.645 $Y=2.42 $X2=0
+ $Y2=0
cc_828 N_A_2789_147#_c_1122_n N_VPWR_c_1364_n 0.00570379f $X=14.565 $Y=2.605
+ $X2=0 $Y2=0
cc_829 N_A_2789_147#_M1009_g N_VPWR_c_1364_n 0.0187486f $X=16.77 $Y=2.795 $X2=0
+ $Y2=0
cc_830 N_A_2789_147#_M1033_g N_VPWR_c_1364_n 0.00593183f $X=17.645 $Y=2.42 $X2=0
+ $Y2=0
cc_831 N_A_2789_147#_c_1130_n N_VPWR_c_1364_n 0.0388577f $X=15.83 $Y=3.57 $X2=0
+ $Y2=0
cc_832 N_A_2789_147#_c_1131_n N_VPWR_c_1364_n 0.0354459f $X=16.725 $Y=3.72 $X2=0
+ $Y2=0
cc_833 N_A_2789_147#_c_1134_n N_VPWR_c_1364_n 0.0109965f $X=15.995 $Y=3.72 $X2=0
+ $Y2=0
cc_834 N_A_2789_147#_c_1185_p N_VPWR_c_1364_n 0.0199629f $X=16.81 $Y=3.635 $X2=0
+ $Y2=0
cc_835 N_A_2789_147#_c_1122_n N_A_2365_445#_c_1749_n 0.0144089f $X=14.565
+ $Y=2.605 $X2=0 $Y2=0
cc_836 N_A_2789_147#_c_1128_n N_A_2365_445#_c_1749_n 0.0112854f $X=14.63 $Y=2.39
+ $X2=0 $Y2=0
cc_837 N_A_2789_147#_M1009_g N_Q_c_1783_n 0.0160686f $X=16.77 $Y=2.795 $X2=0
+ $Y2=0
cc_838 N_A_2789_147#_c_1131_n N_Q_c_1783_n 0.0210086f $X=16.725 $Y=3.72 $X2=0
+ $Y2=0
cc_839 N_A_2789_147#_c_1185_p N_Q_c_1783_n 0.0640489f $X=16.81 $Y=3.635 $X2=0
+ $Y2=0
cc_840 N_A_2789_147#_c_1138_n N_Q_c_1783_n 0.0533362f $X=15.83 $Y=2.86 $X2=0
+ $Y2=0
cc_841 N_A_2789_147#_c_1139_n N_Q_c_1783_n 0.00735756f $X=15.8 $Y=2.695 $X2=0
+ $Y2=0
cc_842 N_A_2789_147#_M1010_g N_Q_c_1781_n 0.0228921f $X=16.51 $Y=0.91 $X2=0
+ $Y2=0
cc_843 N_A_2789_147#_M1009_g N_Q_c_1781_n 0.00283808f $X=16.77 $Y=2.795 $X2=0
+ $Y2=0
cc_844 N_A_2789_147#_c_1118_n N_Q_c_1781_n 0.123741f $X=15.48 $Y=0.66 $X2=0
+ $Y2=0
cc_845 N_A_2789_147#_c_1174_p N_Q_c_1781_n 0.0181781f $X=16.89 $Y=1.67 $X2=0
+ $Y2=0
cc_846 N_A_2789_147#_c_1120_n N_Q_c_1781_n 0.023345f $X=17.645 $Y=1.665 $X2=0
+ $Y2=0
cc_847 N_A_2789_147#_M1009_g N_Q_c_1785_n 0.0100836f $X=16.77 $Y=2.795 $X2=0
+ $Y2=0
cc_848 N_A_2789_147#_c_1118_n N_Q_c_1785_n 0.0205255f $X=15.48 $Y=0.66 $X2=0
+ $Y2=0
cc_849 N_A_2789_147#_c_1185_p N_Q_c_1785_n 0.0350788f $X=16.81 $Y=3.635 $X2=0
+ $Y2=0
cc_850 N_A_2789_147#_c_1137_n N_Q_c_1785_n 0.0221591f $X=15.545 $Y=2.39 $X2=0
+ $Y2=0
cc_851 N_A_2789_147#_c_1138_n N_Q_c_1785_n 0.00336671f $X=15.83 $Y=2.86 $X2=0
+ $Y2=0
cc_852 N_A_2789_147#_c_1120_n N_Q_c_1785_n 0.011804f $X=17.645 $Y=1.665 $X2=0
+ $Y2=0
cc_853 N_A_2789_147#_M1031_g N_VGND_c_1830_n 0.0631194f $X=14.195 $Y=1.075 $X2=0
+ $Y2=0
cc_854 N_A_2789_147#_c_1118_n N_VGND_c_1830_n 0.0283426f $X=15.48 $Y=0.66 $X2=0
+ $Y2=0
cc_855 N_A_2789_147#_M1010_g N_VGND_c_1832_n 0.0613206f $X=16.51 $Y=0.91 $X2=0
+ $Y2=0
cc_856 N_A_2789_147#_M1032_g N_VGND_c_1832_n 0.0683116f $X=17.405 $Y=0.745 $X2=0
+ $Y2=0
cc_857 N_A_2789_147#_c_1174_p N_VGND_c_1832_n 0.0271745f $X=16.89 $Y=1.67 $X2=0
+ $Y2=0
cc_858 N_A_2789_147#_c_1120_n N_VGND_c_1832_n 0.00673191f $X=17.645 $Y=1.665
+ $X2=0 $Y2=0
cc_859 N_A_2789_147#_M1032_g N_VGND_c_1834_n 0.00405414f $X=17.405 $Y=0.745
+ $X2=0 $Y2=0
cc_860 N_A_2789_147#_M1010_g N_VGND_c_1836_n 0.0118525f $X=16.51 $Y=0.91 $X2=0
+ $Y2=0
cc_861 N_A_2789_147#_M1032_g N_VGND_c_1836_n 0.0139641f $X=17.405 $Y=0.745 $X2=0
+ $Y2=0
cc_862 N_A_2789_147#_c_1118_n N_VGND_c_1836_n 0.0439682f $X=15.48 $Y=0.66 $X2=0
+ $Y2=0
cc_863 N_A_2518_445#_M1015_g N_VPWR_c_1355_n 0.0418602f $X=15.44 $Y=3.215 $X2=0
+ $Y2=0
cc_864 N_A_2518_445#_M1015_g N_VPWR_c_1364_n 0.0108618f $X=15.44 $Y=3.215 $X2=0
+ $Y2=0
cc_865 N_A_2518_445#_c_1232_n N_VPWR_c_1364_n 2.62923e-19 $X=12.825 $Y=3.02
+ $X2=0 $Y2=0
cc_866 N_A_2518_445#_c_1234_n N_A_2365_445#_c_1749_n 0.00993334f $X=14.805 $Y=2
+ $X2=0 $Y2=0
cc_867 N_A_2518_445#_M1015_g N_Q_c_1783_n 0.00230901f $X=15.44 $Y=3.215 $X2=0
+ $Y2=0
cc_868 N_A_2518_445#_c_1223_n N_Q_c_1781_n 0.001497f $X=15.09 $Y=1.395 $X2=0
+ $Y2=0
cc_869 N_A_2518_445#_c_1227_n N_Q_c_1781_n 0.0024456f $X=15.44 $Y=1.645 $X2=0
+ $Y2=0
cc_870 N_A_2518_445#_M1015_g N_Q_c_1785_n 0.00304658f $X=15.44 $Y=3.215 $X2=0
+ $Y2=0
cc_871 N_A_2518_445#_c_1223_n N_VGND_c_1830_n 0.029921f $X=15.09 $Y=1.395 $X2=0
+ $Y2=0
cc_872 N_A_2518_445#_c_1234_n N_VGND_c_1830_n 0.0273594f $X=14.805 $Y=2 $X2=0
+ $Y2=0
cc_873 N_A_2518_445#_c_1235_n N_VGND_c_1830_n 0.00407489f $X=14.97 $Y=1.71 $X2=0
+ $Y2=0
cc_874 N_A_2518_445#_c_1227_n N_VGND_c_1830_n 0.00176993f $X=15.44 $Y=1.645
+ $X2=0 $Y2=0
cc_875 N_A_2518_445#_c_1223_n N_VGND_c_1836_n 0.0293328f $X=15.09 $Y=1.395 $X2=0
+ $Y2=0
cc_876 N_A_2518_445#_c_1226_n N_VGND_c_1836_n 0.0033145f $X=13.095 $Y=1.075
+ $X2=0 $Y2=0
cc_877 N_A_3531_107#_c_1313_n N_VPWR_c_1358_n 0.0533757f $X=18.035 $Y=2.19 $X2=0
+ $Y2=0
cc_878 N_A_3531_107#_c_1307_n N_VPWR_c_1358_n 0.00158136f $X=18.2 $Y=1.67 $X2=0
+ $Y2=0
cc_879 N_A_3531_107#_M1021_g N_VPWR_c_1361_n 0.0682136f $X=18.995 $Y=2.965 $X2=0
+ $Y2=0
cc_880 N_A_3531_107#_c_1313_n N_VPWR_c_1361_n 0.0534954f $X=18.035 $Y=2.19 $X2=0
+ $Y2=0
cc_881 N_A_3531_107#_c_1308_n N_VPWR_c_1361_n 0.0298882f $X=18.875 $Y=1.67 $X2=0
+ $Y2=0
cc_882 N_A_3531_107#_c_1309_n N_VPWR_c_1361_n 0.00179471f $X=18.875 $Y=1.67
+ $X2=0 $Y2=0
cc_883 N_A_3531_107#_M1021_g N_VPWR_c_1364_n 0.0151867f $X=18.995 $Y=2.965 $X2=0
+ $Y2=0
cc_884 N_A_3531_107#_M1011_g N_Q_N_c_1809_n 0.0230149f $X=18.995 $Y=0.91 $X2=0
+ $Y2=0
cc_885 N_A_3531_107#_M1021_g N_Q_N_c_1809_n 0.0381317f $X=18.995 $Y=2.965 $X2=0
+ $Y2=0
cc_886 N_A_3531_107#_c_1308_n N_Q_N_c_1809_n 0.0250299f $X=18.875 $Y=1.67 $X2=0
+ $Y2=0
cc_887 N_A_3531_107#_c_1309_n N_Q_N_c_1809_n 0.0353277f $X=18.875 $Y=1.67 $X2=0
+ $Y2=0
cc_888 N_A_3531_107#_c_1305_n N_VGND_c_1832_n 0.0526461f $X=17.795 $Y=0.745
+ $X2=0 $Y2=0
cc_889 N_A_3531_107#_M1011_g N_VGND_c_1834_n 0.053985f $X=18.995 $Y=0.91 $X2=0
+ $Y2=0
cc_890 N_A_3531_107#_c_1305_n N_VGND_c_1834_n 0.068177f $X=17.795 $Y=0.745 $X2=0
+ $Y2=0
cc_891 N_A_3531_107#_c_1307_n N_VGND_c_1834_n 0.00530721f $X=18.2 $Y=1.67 $X2=0
+ $Y2=0
cc_892 N_A_3531_107#_c_1308_n N_VGND_c_1834_n 0.0684373f $X=18.875 $Y=1.67 $X2=0
+ $Y2=0
cc_893 N_A_3531_107#_c_1309_n N_VGND_c_1834_n 0.00163586f $X=18.875 $Y=1.67
+ $X2=0 $Y2=0
cc_894 N_A_3531_107#_M1011_g N_VGND_c_1836_n 0.0115807f $X=18.995 $Y=0.91 $X2=0
+ $Y2=0
cc_895 N_A_3531_107#_c_1305_n N_VGND_c_1836_n 0.0315421f $X=17.795 $Y=0.745
+ $X2=0 $Y2=0
cc_896 N_VPWR_c_1364_n N_A_268_659#_M1000_s 0.00311481f $X=18.855 $Y=3.59 $X2=0
+ $Y2=3.985
cc_897 N_VPWR_c_1343_n N_A_268_659#_c_1472_n 0.045143f $X=1.055 $Y=2.785
+ $X2=0.24 $Y2=4.07
cc_898 N_VPWR_c_1346_n N_A_268_659#_c_1472_n 0.0197671f $X=2.265 $Y=3.505
+ $X2=0.24 $Y2=4.07
cc_899 N_VPWR_c_1364_n N_A_268_659#_c_1472_n 0.0231871f $X=18.855 $Y=3.59
+ $X2=0.24 $Y2=4.07
cc_900 N_VPWR_c_1346_n N_A_268_659#_c_1475_n 0.0451328f $X=2.265 $Y=3.505 $X2=0
+ $Y2=0
cc_901 N_VPWR_c_1364_n N_A_268_659#_c_1475_n 0.0257489f $X=18.855 $Y=3.59 $X2=0
+ $Y2=0
cc_902 N_VPWR_c_1343_n N_A_268_659#_c_1476_n 0.0150665f $X=1.055 $Y=2.785
+ $X2=0.24 $Y2=4.07
cc_903 N_VPWR_c_1364_n N_A_268_659#_c_1477_n 0.00913626f $X=18.855 $Y=3.59
+ $X2=19.44 $Y2=4.07
cc_904 N_VPWR_c_1346_n N_A_581_659#_c_1504_n 0.0184508f $X=2.265 $Y=3.505
+ $X2=0.24 $Y2=4.07
cc_905 N_VPWR_c_1364_n N_A_581_659#_c_1504_n 0.0168135f $X=18.855 $Y=3.59
+ $X2=0.24 $Y2=4.07
cc_906 N_VPWR_c_1364_n N_A_581_659#_c_1505_n 0.0301678f $X=18.855 $Y=3.59 $X2=0
+ $Y2=0
cc_907 N_VPWR_c_1346_n N_A_581_659#_c_1508_n 0.0089875f $X=2.265 $Y=3.505
+ $X2=0.24 $Y2=4.07
cc_908 N_VPWR_c_1364_n N_A_581_659#_c_1508_n 0.00955363f $X=18.855 $Y=3.59
+ $X2=0.24 $Y2=4.07
cc_909 N_VPWR_c_1364_n N_A_581_659#_c_1511_n 0.0184183f $X=18.855 $Y=3.59
+ $X2=19.44 $Y2=4.07
cc_910 N_VPWR_c_1364_n N_A_581_659#_c_1512_n 0.0177877f $X=18.855 $Y=3.59
+ $X2=19.44 $Y2=4.07
cc_911 N_VPWR_c_1364_n N_A_581_659#_c_1513_n 0.00927265f $X=18.855 $Y=3.59 $X2=0
+ $Y2=0
cc_912 N_VPWR_c_1364_n N_A_567_107#_c_1564_n 0.0216587f $X=18.855 $Y=3.59 $X2=0
+ $Y2=0
cc_913 N_VPWR_c_1349_n N_A_567_107#_c_1565_n 0.00742195f $X=7.125 $Y=3.59 $X2=0
+ $Y2=0
cc_914 N_VPWR_c_1364_n N_A_567_107#_c_1565_n 0.0628619f $X=18.855 $Y=3.59 $X2=0
+ $Y2=0
cc_915 N_VPWR_c_1364_n N_A_567_107#_c_1568_n 0.00929118f $X=18.855 $Y=3.59 $X2=0
+ $Y2=0
cc_916 N_VPWR_c_1349_n N_A_567_107#_c_1621_n 0.0103845f $X=7.125 $Y=3.59 $X2=0
+ $Y2=0
cc_917 N_VPWR_c_1364_n N_A_567_107#_c_1621_n 0.0135697f $X=18.855 $Y=3.59 $X2=0
+ $Y2=0
cc_918 N_VPWR_M1035_d N_A_567_107#_c_1629_n 0.0189626f $X=6.345 $Y=2.715 $X2=0
+ $Y2=0
cc_919 N_VPWR_c_1349_n N_A_567_107#_c_1629_n 0.0499958f $X=7.125 $Y=3.59 $X2=0
+ $Y2=0
cc_920 N_VPWR_c_1364_n N_A_567_107#_c_1629_n 0.0151563f $X=18.855 $Y=3.59 $X2=0
+ $Y2=0
cc_921 N_VPWR_c_1364_n N_A_567_107#_c_1573_n 0.0511721f $X=18.855 $Y=3.59 $X2=0
+ $Y2=0
cc_922 N_VPWR_c_1364_n N_A_567_107#_c_1576_n 0.00683296f $X=18.855 $Y=3.59 $X2=0
+ $Y2=0
cc_923 N_VPWR_c_1364_n N_A_567_107#_c_1579_n 0.0128366f $X=18.855 $Y=3.59 $X2=0
+ $Y2=0
cc_924 N_VPWR_c_1352_n N_A_2365_445#_c_1742_n 0.0118751f $X=10.62 $Y=2.89
+ $X2=0.24 $Y2=4.07
cc_925 N_VPWR_c_1364_n N_A_2365_445#_c_1742_n 0.0239292f $X=18.855 $Y=3.59
+ $X2=0.24 $Y2=4.07
cc_926 N_VPWR_c_1355_n N_A_2365_445#_c_1743_n 0.00699923f $X=15.05 $Y=2.86 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1364_n N_A_2365_445#_c_1743_n 0.0764229f $X=18.855 $Y=3.59 $X2=0
+ $Y2=0
cc_928 N_VPWR_c_1352_n N_A_2365_445#_c_1746_n 0.00107828f $X=10.62 $Y=2.89
+ $X2=0.24 $Y2=4.07
cc_929 N_VPWR_c_1364_n N_A_2365_445#_c_1746_n 0.0121864f $X=18.855 $Y=3.59
+ $X2=0.24 $Y2=4.07
cc_930 N_VPWR_c_1355_n N_A_2365_445#_c_1749_n 0.0715294f $X=15.05 $Y=2.86
+ $X2=19.44 $Y2=4.07
cc_931 N_VPWR_c_1364_n N_A_2365_445#_c_1749_n 0.0335382f $X=18.855 $Y=3.59
+ $X2=19.44 $Y2=4.07
cc_932 N_VPWR_c_1364_n N_Q_c_1783_n 0.0228057f $X=18.855 $Y=3.59 $X2=0.24
+ $Y2=4.07
cc_933 N_VPWR_c_1361_n N_Q_N_c_1809_n 0.0865233f $X=18.605 $Y=2.34 $X2=9.84
+ $Y2=4.07
cc_934 N_VPWR_c_1364_n N_Q_N_c_1809_n 0.0444416f $X=18.855 $Y=3.59 $X2=9.84
+ $Y2=4.07
cc_935 N_A_268_659#_c_1475_n N_A_581_659#_c_1504_n 0.0242126f $X=3.43 $Y=3.01
+ $X2=0.24 $Y2=4.07
cc_936 N_A_268_659#_c_1477_n N_A_581_659#_c_1504_n 0.0105547f $X=3.595 $Y=3.2
+ $X2=0.24 $Y2=4.07
cc_937 N_A_268_659#_c_1475_n N_A_581_659#_c_1505_n 0.00429912f $X=3.43 $Y=3.01
+ $X2=0 $Y2=0
cc_938 N_A_268_659#_c_1477_n N_A_581_659#_c_1505_n 0.0163505f $X=3.595 $Y=3.2
+ $X2=0 $Y2=0
cc_939 N_A_268_659#_c_1475_n N_A_581_659#_c_1511_n 0.00839273f $X=3.43 $Y=3.01
+ $X2=19.44 $Y2=4.07
cc_940 N_A_268_659#_c_1477_n N_A_581_659#_c_1511_n 0.0115725f $X=3.595 $Y=3.2
+ $X2=19.44 $Y2=4.07
cc_941 N_A_268_659#_c_1475_n N_A_567_107#_c_1584_n 0.0073868f $X=3.43 $Y=3.01
+ $X2=0 $Y2=0
cc_942 N_A_581_659#_c_1512_n N_A_567_107#_c_1563_n 0.0771097f $X=4.99 $Y=2.765
+ $X2=0 $Y2=0
cc_943 N_A_581_659#_c_1521_n N_A_567_107#_c_1563_n 0.0123662f $X=4.03 $Y=2.765
+ $X2=0 $Y2=0
cc_944 N_A_581_659#_c_1505_n N_A_567_107#_c_1564_n 0.00169592f $X=3.86 $Y=3.695
+ $X2=0 $Y2=0
cc_945 N_A_581_659#_c_1511_n N_A_567_107#_c_1564_n 0.0387899f $X=3.945 $Y=3.61
+ $X2=0 $Y2=0
cc_946 N_A_581_659#_c_1512_n N_A_567_107#_c_1564_n 0.0200383f $X=4.99 $Y=2.765
+ $X2=0 $Y2=0
cc_947 N_A_581_659#_c_1513_n N_A_567_107#_c_1564_n 0.0133572f $X=5.155 $Y=3.2
+ $X2=0 $Y2=0
cc_948 N_A_581_659#_c_1513_n N_A_567_107#_c_1565_n 0.0144411f $X=5.155 $Y=3.2
+ $X2=0 $Y2=0
cc_949 N_A_581_659#_c_1505_n N_A_567_107#_c_1568_n 0.0102055f $X=3.86 $Y=3.695
+ $X2=0 $Y2=0
cc_950 N_A_567_107#_c_1573_n A_1528_579# 0.00102794f $X=9.105 $Y=3.37 $X2=0
+ $Y2=0
cc_951 N_A_567_107#_c_1557_n N_VGND_M1003_d 0.00594047f $X=7.3 $Y=1.34 $X2=0
+ $Y2=0
cc_952 N_A_567_107#_c_1550_n N_VGND_c_1824_n 0.0139735f $X=3.51 $Y=0.91 $X2=0
+ $Y2=0
cc_953 N_A_567_107#_c_1552_n N_VGND_c_1824_n 0.0428011f $X=5.05 $Y=2.33 $X2=0
+ $Y2=0
cc_954 N_A_567_107#_c_1555_n N_VGND_c_1824_n 0.00489946f $X=5.135 $Y=0.35 $X2=0
+ $Y2=0
cc_955 N_A_567_107#_c_1553_n N_VGND_c_1826_n 0.00477932f $X=5.825 $Y=0.35 $X2=0
+ $Y2=0
cc_956 N_A_567_107#_c_1618_n N_VGND_c_1826_n 0.0253511f $X=5.91 $Y=1.255 $X2=0
+ $Y2=0
cc_957 N_A_567_107#_c_1557_n N_VGND_c_1826_n 0.0633953f $X=7.3 $Y=1.34 $X2=0
+ $Y2=0
cc_958 N_A_567_107#_c_1550_n N_VGND_c_1836_n 0.0237358f $X=3.51 $Y=0.91 $X2=0
+ $Y2=0
cc_959 N_A_567_107#_c_1552_n N_VGND_c_1836_n 0.0201148f $X=5.05 $Y=2.33 $X2=0
+ $Y2=0
cc_960 N_A_567_107#_c_1553_n N_VGND_c_1836_n 0.0335185f $X=5.825 $Y=0.35 $X2=0
+ $Y2=0
cc_961 N_A_567_107#_c_1555_n N_VGND_c_1836_n 0.00777234f $X=5.135 $Y=0.35 $X2=0
+ $Y2=0
cc_962 N_A_567_107#_c_1618_n N_VGND_c_1836_n 0.0199629f $X=5.91 $Y=1.255 $X2=0
+ $Y2=0
cc_963 N_A_567_107#_c_1559_n N_VGND_c_1836_n 0.0232655f $X=2.975 $Y=0.745 $X2=0
+ $Y2=0
cc_964 N_A_567_107#_c_1561_n N_VGND_c_1836_n 0.00192217f $X=8 $Y=1.11 $X2=0
+ $Y2=0
cc_965 N_A_567_107#_c_1550_n A_723_107# 0.00125759f $X=3.51 $Y=0.91 $X2=0 $Y2=0
cc_966 N_A_567_107#_c_1558_n N_A_1454_173#_M1012_d 9.14618e-19 $X=7.835 $Y=1.34
+ $X2=0 $Y2=0
cc_967 N_A_567_107#_c_1673_n N_A_1454_173#_M1012_d 0.00162126f $X=7.385 $Y=1.34
+ $X2=0 $Y2=0
cc_968 N_A_567_107#_c_1558_n N_A_1454_173#_c_1935_n 0.00934732f $X=7.835 $Y=1.34
+ $X2=0 $Y2=0
cc_969 N_A_567_107#_c_1561_n N_A_1454_173#_c_1935_n 0.0213165f $X=8 $Y=1.11
+ $X2=0 $Y2=0
cc_970 N_A_567_107#_c_1557_n N_A_1454_173#_c_1938_n 0.00165922f $X=7.3 $Y=1.34
+ $X2=0 $Y2=0
cc_971 N_A_567_107#_c_1558_n N_A_1454_173#_c_1938_n 0.00791107f $X=7.835 $Y=1.34
+ $X2=0 $Y2=0
cc_972 N_A_567_107#_c_1673_n N_A_1454_173#_c_1938_n 0.0120483f $X=7.385 $Y=1.34
+ $X2=0 $Y2=0
cc_973 N_A_567_107#_c_1561_n N_A_1454_173#_c_1938_n 0.0083639f $X=8 $Y=1.11
+ $X2=0 $Y2=0
cc_974 N_Q_c_1781_n N_VGND_c_1832_n 0.0611058f $X=16.12 $Y=0.66 $X2=0 $Y2=0
cc_975 N_Q_c_1781_n N_VGND_c_1836_n 0.0313203f $X=16.12 $Y=0.66 $X2=0 $Y2=0
cc_976 N_Q_N_c_1809_n N_VGND_c_1834_n 0.0611641f $X=19.385 $Y=0.66 $X2=0 $Y2=0
cc_977 N_Q_N_c_1809_n N_VGND_c_1836_n 0.0336637f $X=19.385 $Y=0.66 $X2=0 $Y2=0
cc_978 N_VGND_c_1836_n A_425_107# 0.00286287f $X=18.95 $Y=0.48 $X2=0 $Y2=0
cc_979 N_VGND_c_1836_n A_723_107# 0.006628f $X=18.95 $Y=0.48 $X2=0 $Y2=0
cc_980 N_VGND_c_1836_n N_A_1454_173#_c_1935_n 0.110924f $X=18.95 $Y=0.48 $X2=0
+ $Y2=0
cc_981 N_VGND_c_1826_n N_A_1454_173#_c_1938_n 0.0375185f $X=6.26 $Y=0.48 $X2=0
+ $Y2=0
cc_982 N_VGND_c_1836_n N_A_1454_173#_c_1938_n 0.0244721f $X=18.95 $Y=0.48 $X2=0
+ $Y2=0
