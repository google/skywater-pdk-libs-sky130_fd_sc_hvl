* File: sky130_fd_sc_hvl__probec_p_8.pxi.spice
* Created: Fri Aug 28 09:39:15 2020
* 
x_PM_SKY130_FD_SC_HVL__PROBEC_P_8%VNB N_VNB_M1003_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__PROBEC_P_8%VNB
x_PM_SKY130_FD_SC_HVL__PROBEC_P_8%VPB N_VPB_M1006_b VPB N_VPB_c_52_p VPB
+ PM_SKY130_FD_SC_HVL__PROBEC_P_8%VPB
x_PM_SKY130_FD_SC_HVL__PROBEC_P_8%A N_A_M1006_g N_A_c_141_n N_A_M1003_g
+ N_A_c_143_n N_A_c_144_n N_A_M1008_g N_A_M1007_g N_A_c_145_n N_A_M1015_g
+ N_A_M1019_g N_A_c_146_n A A A A N_A_c_147_n PM_SKY130_FD_SC_HVL__PROBEC_P_8%A
x_PM_SKY130_FD_SC_HVL__PROBEC_P_8%A_45_443# N_A_45_443#_M1003_d
+ N_A_45_443#_M1008_d N_A_45_443#_M1006_s N_A_45_443#_M1007_s
+ N_A_45_443#_M1001_g N_A_45_443#_c_238_n N_A_45_443#_M1000_g
+ N_A_45_443#_M1002_g N_A_45_443#_c_241_n N_A_45_443#_M1004_g
+ N_A_45_443#_M1009_g N_A_45_443#_c_244_n N_A_45_443#_M1005_g
+ N_A_45_443#_M1013_g N_A_45_443#_c_247_n N_A_45_443#_M1010_g
+ N_A_45_443#_M1014_g N_A_45_443#_c_250_n N_A_45_443#_M1011_g
+ N_A_45_443#_M1018_g N_A_45_443#_c_253_n N_A_45_443#_M1012_g
+ N_A_45_443#_M1020_g N_A_45_443#_c_256_n N_A_45_443#_M1016_g
+ N_A_45_443#_M1021_g N_A_45_443#_c_259_n N_A_45_443#_M1017_g
+ N_A_45_443#_c_272_n N_A_45_443#_c_234_n N_A_45_443#_c_263_n
+ N_A_45_443#_c_265_n N_A_45_443#_c_280_n N_A_45_443#_c_417_p
+ N_A_45_443#_c_282_n N_A_45_443#_c_286_n N_A_45_443#_c_235_n
+ N_A_45_443#_c_236_n N_A_45_443#_c_267_n N_A_45_443#_c_268_n
+ N_A_45_443#_c_294_n N_A_45_443#_c_297_n N_A_45_443#_c_237_n
+ PM_SKY130_FD_SC_HVL__PROBEC_P_8%A_45_443#
x_PM_SKY130_FD_SC_HVL__PROBEC_P_8%VPWR N_VPWR_M1006_d N_VPWR_M1019_d
+ N_VPWR_M1004_s N_VPWR_M1010_s N_VPWR_M1012_s N_VPWR_M1017_s N_VPWR_c_487_n
+ N_VPWR_c_490_n N_VPWR_c_493_n N_VPWR_c_496_n N_VPWR_c_499_n N_VPWR_c_500_n
+ N_VPWR_c_501_n N_VPWR_c_504_n N_VPWR_c_507_n N_VPWR_c_510_n VPWR
+ N_VPWR_c_530_n N_VPWR_c_560_n N_VPWR_c_565_n N_VPWR_c_570_n N_VPWR_c_514_n
+ N_VPWR_c_517_n N_VPWR_c_520_n N_VPWR_c_486_n N_VPWR_c_524_n VPWR
+ PM_SKY130_FD_SC_HVL__PROBEC_P_8%VPWR
x_PM_SKY130_FD_SC_HVL__PROBEC_P_8%noxref_6 N_noxref_6_M1001_d N_noxref_6_M1009_d
+ N_noxref_6_M1014_d N_noxref_6_M1020_d N_noxref_6_M1000_d N_noxref_6_M1005_d
+ N_noxref_6_M1011_d N_noxref_6_M1016_d N_noxref_6_c_657_n N_noxref_6_c_645_n
+ N_noxref_6_c_652_n N_noxref_6_c_665_n N_noxref_6_c_646_n N_noxref_6_c_670_n
+ N_noxref_6_c_647_n N_noxref_6_c_653_n N_noxref_6_c_678_n N_noxref_6_c_680_n
+ N_noxref_6_c_648_n N_noxref_6_c_685_n N_noxref_6_c_689_n N_noxref_6_c_654_n
+ N_noxref_6_c_695_n N_noxref_6_c_698_n N_noxref_6_c_649_n N_noxref_6_c_753_n
+ N_noxref_6_R23_noxref_neg N_noxref_6_c_758_n N_noxref_6_c_759_n
+ PM_SKY130_FD_SC_HVL__PROBEC_P_8%noxref_6
x_PM_SKY130_FD_SC_HVL__PROBEC_P_8%VGND N_VGND_M1003_s N_VGND_M1015_s
+ N_VGND_M1002_s N_VGND_M1013_s N_VGND_M1018_s N_VGND_M1021_s N_VGND_c_804_n
+ N_VGND_c_805_n VGND N_VGND_c_807_n N_VGND_c_809_n N_VGND_c_811_n
+ N_VGND_c_813_n N_VGND_c_814_n N_VGND_c_815_n N_VGND_c_816_n N_VGND_c_817_n
+ N_VGND_c_818_n N_VGND_c_819_n N_VGND_c_820_n N_VGND_c_821_n N_VGND_c_823_n
+ VGND PM_SKY130_FD_SC_HVL__PROBEC_P_8%VGND
x_PM_SKY130_FD_SC_HVL__PROBEC_P_8%X X N_X_c_930_n N_X_c_928_n N_X_R23_noxref_pos
+ PM_SKY130_FD_SC_HVL__PROBEC_P_8%X
cc_1 N_VNB_M1003_b N_A_c_141_n 0.0456634f $X=-0.33 $Y=-0.365 $X2=0.78 $Y2=1.565
cc_2 N_VNB_c_2_p N_A_c_141_n 5.58874e-19 $X=0.24 $Y=0 $X2=0.78 $Y2=1.565
cc_3 N_VNB_M1003_b N_A_c_143_n 0.0274014f $X=-0.33 $Y=-0.365 $X2=1.57 $Y2=1.815
cc_4 N_VNB_M1003_b N_A_c_144_n 0.0391903f $X=-0.33 $Y=-0.365 $X2=1.82 $Y2=1.565
cc_5 N_VNB_M1003_b N_A_c_145_n 0.0372172f $X=-0.33 $Y=-0.365 $X2=2.6 $Y2=1.565
cc_6 N_VNB_M1003_b N_A_c_146_n 0.0267973f $X=-0.33 $Y=-0.365 $X2=0.77 $Y2=1.815
cc_7 N_VNB_M1003_b N_A_c_147_n 0.0504375f $X=-0.33 $Y=-0.365 $X2=2.6 $Y2=1.815
cc_8 N_VNB_M1003_b N_A_45_443#_M1001_g 0.0402362f $X=-0.33 $Y=-0.365 $X2=1.82
+ $Y2=2.965
cc_9 N_VNB_M1003_b N_A_45_443#_M1002_g 0.0400604f $X=-0.33 $Y=-0.365 $X2=2.6
+ $Y2=2.965
cc_10 N_VNB_M1003_b N_A_45_443#_M1009_g 0.0398303f $X=-0.33 $Y=-0.365 $X2=0
+ $Y2=0
cc_11 N_VNB_M1003_b N_A_45_443#_M1013_g 0.0397623f $X=-0.33 $Y=-0.365 $X2=1.82
+ $Y2=1.815
cc_12 N_VNB_M1003_b N_A_45_443#_M1014_g 0.0403249f $X=-0.33 $Y=-0.365 $X2=0
+ $Y2=0
cc_13 N_VNB_M1003_b N_A_45_443#_M1018_g 0.0406374f $X=-0.33 $Y=-0.365 $X2=0
+ $Y2=0
cc_14 N_VNB_M1003_b N_A_45_443#_M1020_g 0.03984f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_15 N_VNB_M1003_b N_A_45_443#_M1021_g 0.0484728f $X=-0.33 $Y=-0.365 $X2=0
+ $Y2=0
cc_16 N_VNB_M1003_b N_A_45_443#_c_234_n 0.0201484f $X=-0.33 $Y=-0.365 $X2=0
+ $Y2=0
cc_17 N_VNB_M1003_b N_A_45_443#_c_235_n 0.00170227f $X=-0.33 $Y=-0.365 $X2=0
+ $Y2=0
cc_18 N_VNB_M1003_b N_A_45_443#_c_236_n 0.00131963f $X=-0.33 $Y=-0.365 $X2=0
+ $Y2=0
cc_19 N_VNB_M1003_b N_A_45_443#_c_237_n 0.219442f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_20 N_VNB_M1003_b N_VPWR_c_486_n 0.110666f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_21 N_VNB_M1003_b N_noxref_6_c_645_n 0.00865581f $X=-0.33 $Y=-0.365 $X2=1.735
+ $Y2=1.815
cc_22 N_VNB_M1003_b N_noxref_6_c_646_n 0.00805267f $X=-0.33 $Y=-0.365 $X2=0
+ $Y2=0
cc_23 N_VNB_M1003_b N_noxref_6_c_647_n 0.00270308f $X=-0.33 $Y=-0.365 $X2=0
+ $Y2=0
cc_24 N_VNB_M1003_b N_noxref_6_c_648_n 0.00157904f $X=-0.33 $Y=-0.365 $X2=0
+ $Y2=0
cc_25 N_VNB_M1003_b N_noxref_6_c_649_n 0.00159871f $X=-0.33 $Y=-0.365 $X2=0
+ $Y2=0
cc_26 N_VNB_M1003_b N_noxref_6_R23_noxref_neg 0.0803921f $X=-0.33 $Y=-0.365
+ $X2=0 $Y2=0
cc_27 N_VNB_c_2_p N_noxref_6_R23_noxref_neg 0.0282792f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_28 N_VNB_M1003_b N_VGND_c_804_n 0.0113819f $X=-0.33 $Y=-0.365 $X2=2.6
+ $Y2=1.08
cc_29 N_VNB_M1003_b N_VGND_c_805_n 0.0377886f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_30 N_VNB_M1003_b VGND 0.00539689f $X=-0.33 $Y=-0.365 $X2=1.735 $Y2=1.815
cc_31 N_VNB_M1003_b N_VGND_c_807_n 0.090476f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_32 N_VNB_c_2_p N_VGND_c_807_n 0.00538291f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_33 N_VNB_M1003_b N_VGND_c_809_n 0.0421797f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_34 N_VNB_c_2_p N_VGND_c_809_n 0.00247336f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_35 N_VNB_M1003_b N_VGND_c_811_n 0.251098f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_36 N_VNB_c_2_p N_VGND_c_811_n 0.0166628f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_37 N_VNB_M1003_b N_VGND_c_813_n 0.00648157f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_38 N_VNB_M1003_b N_VGND_c_814_n 0.00846255f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_39 N_VNB_M1003_b N_VGND_c_815_n 0.00648157f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_40 N_VNB_M1003_b N_VGND_c_816_n 0.00846255f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_41 N_VNB_M1003_b N_VGND_c_817_n 0.00659769f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_42 N_VNB_M1003_b N_VGND_c_818_n 0.0125653f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_43 N_VNB_M1003_b N_VGND_c_819_n 0.00867017f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_44 N_VNB_M1003_b N_VGND_c_820_n 0.0133169f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_45 N_VNB_M1003_b N_VGND_c_821_n 0.223127f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_46 N_VNB_c_2_p N_VGND_c_821_n 0.035463f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_47 N_VNB_M1003_b N_VGND_c_823_n 0.142767f $X=-0.33 $Y=-0.365 $X2=0 $Y2=0
cc_48 N_VNB_c_2_p N_VGND_c_823_n 1.02751f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_49 N_VNB_M1003_b N_X_R23_noxref_pos 0.00262201f $X=-0.33 $Y=-0.365 $X2=1.82
+ $Y2=1.565
cc_50 N_VPB_M1006_b N_A_M1006_g 0.0429652f $X=-0.33 $Y=1.885 $X2=0.76 $Y2=2.965
cc_51 VPB N_A_M1006_g 0.00970178f $X=0 $Y=3.955 $X2=0.76 $Y2=2.965
cc_52 N_VPB_c_52_p N_A_M1006_g 0.0148199f $X=9.36 $Y=4.07 $X2=0.76 $Y2=2.965
cc_53 N_VPB_M1006_b N_A_c_143_n 0.0193995f $X=-0.33 $Y=1.885 $X2=1.57 $Y2=1.815
cc_54 N_VPB_M1006_b N_A_M1007_g 0.0378158f $X=-0.33 $Y=1.885 $X2=1.82 $Y2=2.965
cc_55 VPB N_A_M1007_g 0.00970178f $X=0 $Y=3.955 $X2=1.82 $Y2=2.965
cc_56 N_VPB_c_52_p N_A_M1007_g 0.013528f $X=9.36 $Y=4.07 $X2=1.82 $Y2=2.965
cc_57 N_VPB_M1006_b N_A_M1019_g 0.0357299f $X=-0.33 $Y=1.885 $X2=2.6 $Y2=2.965
cc_58 VPB N_A_M1019_g 0.00970178f $X=0 $Y=3.955 $X2=2.6 $Y2=2.965
cc_59 N_VPB_c_52_p N_A_M1019_g 0.0135178f $X=9.36 $Y=4.07 $X2=2.6 $Y2=2.965
cc_60 N_VPB_M1006_b N_A_c_146_n 0.0144517f $X=-0.33 $Y=1.885 $X2=0.77 $Y2=1.815
cc_61 N_VPB_M1006_b N_A_c_147_n 0.0294867f $X=-0.33 $Y=1.885 $X2=2.6 $Y2=1.815
cc_62 N_VPB_M1006_b N_A_45_443#_c_238_n 0.0324045f $X=-0.33 $Y=1.885 $X2=2.6
+ $Y2=1.565
cc_63 VPB N_A_45_443#_c_238_n 0.00970178f $X=0 $Y=3.955 $X2=2.6 $Y2=1.565
cc_64 N_VPB_c_52_p N_A_45_443#_c_238_n 0.0135156f $X=9.36 $Y=4.07 $X2=2.6
+ $Y2=1.565
cc_65 N_VPB_M1006_b N_A_45_443#_c_241_n 0.0320824f $X=-0.33 $Y=1.885 $X2=0.77
+ $Y2=1.815
cc_66 VPB N_A_45_443#_c_241_n 0.00970178f $X=0 $Y=3.955 $X2=0.77 $Y2=1.815
cc_67 N_VPB_c_52_p N_A_45_443#_c_241_n 0.0135156f $X=9.36 $Y=4.07 $X2=0.77
+ $Y2=1.815
cc_68 N_VPB_M1006_b N_A_45_443#_c_244_n 0.0424935f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_69 VPB N_A_45_443#_c_244_n 0.00917643f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_70 N_VPB_c_52_p N_A_45_443#_c_244_n 0.0130128f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_71 N_VPB_M1006_b N_A_45_443#_c_247_n 0.042862f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_72 VPB N_A_45_443#_c_247_n 0.00915454f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_73 N_VPB_c_52_p N_A_45_443#_c_247_n 0.0129919f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_74 N_VPB_M1006_b N_A_45_443#_c_250_n 0.0332756f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_75 VPB N_A_45_443#_c_250_n 0.00963611f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_76 N_VPB_c_52_p N_A_45_443#_c_250_n 0.0134528f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_77 N_VPB_M1006_b N_A_45_443#_c_253_n 0.0321055f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_78 VPB N_A_45_443#_c_253_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_79 N_VPB_c_52_p N_A_45_443#_c_253_n 0.0135156f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_80 N_VPB_M1006_b N_A_45_443#_c_256_n 0.0407709f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_81 VPB N_A_45_443#_c_256_n 0.00926399f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_82 N_VPB_c_52_p N_A_45_443#_c_256_n 0.0130966f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_83 N_VPB_M1006_b N_A_45_443#_c_259_n 0.0495025f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_84 VPB N_A_45_443#_c_259_n 0.00910227f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_85 N_VPB_c_52_p N_A_45_443#_c_259_n 0.0129494f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_86 N_VPB_M1006_b N_A_45_443#_c_234_n 0.00998322f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_87 VPB N_A_45_443#_c_263_n 4.22267e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_88 N_VPB_c_52_p N_A_45_443#_c_263_n 0.00452125f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_89 N_VPB_M1006_b N_A_45_443#_c_265_n 0.00764217f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_90 N_VPB_M1006_b N_A_45_443#_c_235_n 0.00244843f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_91 N_VPB_M1006_b N_A_45_443#_c_267_n 0.00526456f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_92 N_VPB_M1006_b N_A_45_443#_c_268_n 0.00486023f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_93 N_VPB_M1006_b N_A_45_443#_c_237_n 0.174554f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_94 N_VPB_M1006_b N_VPWR_c_487_n 0.0010569f $X=-0.33 $Y=1.885 $X2=2.6 $Y2=1.08
cc_95 VPB N_VPWR_c_487_n 0.00362936f $X=0 $Y=3.955 $X2=2.6 $Y2=1.08
cc_96 N_VPB_c_52_p N_VPWR_c_487_n 0.054215f $X=9.36 $Y=4.07 $X2=2.6 $Y2=1.08
cc_97 N_VPB_M1006_b N_VPWR_c_490_n 0.0010569f $X=-0.33 $Y=1.885 $X2=2.6
+ $Y2=2.965
cc_98 VPB N_VPWR_c_490_n 0.00262607f $X=0 $Y=3.955 $X2=2.6 $Y2=2.965
cc_99 N_VPB_c_52_p N_VPWR_c_490_n 0.0405322f $X=9.36 $Y=4.07 $X2=2.6 $Y2=2.965
cc_100 N_VPB_M1006_b N_VPWR_c_493_n 0.0010569f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_493_n 0.00260627f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_102 N_VPB_c_52_p N_VPWR_c_493_n 0.0405322f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_103 N_VPB_M1006_b N_VPWR_c_496_n 0.0010569f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_104 VPB N_VPWR_c_496_n 0.00262607f $X=0 $Y=3.955 $X2=0.635 $Y2=1.58
cc_105 N_VPB_c_52_p N_VPWR_c_496_n 0.0405322f $X=9.36 $Y=4.07 $X2=0.635 $Y2=1.58
cc_106 N_VPB_M1006_b N_VPWR_c_499_n 0.0076911f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_107 N_VPB_M1006_b N_VPWR_c_500_n 0.0467833f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_108 N_VPB_M1006_b N_VPWR_c_501_n 0.00105831f $X=-0.33 $Y=1.885 $X2=1.82
+ $Y2=1.815
cc_109 VPB N_VPWR_c_501_n 0.00279423f $X=0 $Y=3.955 $X2=1.82 $Y2=1.815
cc_110 N_VPB_c_52_p N_VPWR_c_501_n 0.0413412f $X=9.36 $Y=4.07 $X2=1.82 $Y2=1.815
cc_111 N_VPB_M1006_b N_VPWR_c_504_n 0.00105831f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_504_n 0.0038448f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_113 N_VPB_c_52_p N_VPWR_c_504_n 0.0545489f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_114 N_VPB_M1006_b N_VPWR_c_507_n 0.00105831f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_507_n 0.00383421f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_116 N_VPB_c_52_p N_VPWR_c_507_n 0.0545489f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_117 N_VPB_M1006_b N_VPWR_c_510_n 0.00105831f $X=-0.33 $Y=1.885 $X2=1.2
+ $Y2=1.697
cc_118 VPB N_VPWR_c_510_n 0.00384715f $X=0 $Y=3.955 $X2=1.2 $Y2=1.697
cc_119 N_VPB_c_52_p N_VPWR_c_510_n 0.0545489f $X=9.36 $Y=4.07 $X2=1.2 $Y2=1.697
cc_120 N_VPB_M1006_b VPWR 0.0052729f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_121 N_VPB_M1006_b N_VPWR_c_514_n 0.00270841f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_514_n 0.00513943f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_123 N_VPB_c_52_p N_VPWR_c_514_n 0.0771568f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_124 N_VPB_M1006_b N_VPWR_c_517_n 0.0010569f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_517_n 0.00530115f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_126 N_VPB_c_52_p N_VPWR_c_517_n 0.0847725f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_127 N_VPB_M1006_b N_VPWR_c_520_n 0.0133169f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_128 N_VPB_M1006_b N_VPWR_c_486_n 0.111007f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_486_n 0.035463f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_130 N_VPB_c_52_p N_VPWR_c_486_n 8.1781e-19 $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_131 N_VPB_M1006_b N_VPWR_c_524_n 0.0403869f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_524_n 1.01754f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_133 N_VPB_c_52_p N_VPWR_c_524_n 0.0332942f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_134 N_VPB_M1006_b N_noxref_6_c_652_n 0.00186667f $X=-0.33 $Y=1.885 $X2=1.735
+ $Y2=1.73
cc_135 N_VPB_M1006_b N_noxref_6_c_653_n 0.00267366f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_136 N_VPB_M1006_b N_noxref_6_c_654_n 0.0017141f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_137 N_VPB_M1006_b N_noxref_6_R23_noxref_neg 0.0789898f $X=-0.33 $Y=1.885
+ $X2=0 $Y2=0
cc_138 VPB N_noxref_6_R23_noxref_neg 0.0282792f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_139 N_VPB_M1006_b N_X_c_928_n 0.00341864f $X=-0.33 $Y=1.885 $X2=1.57
+ $Y2=1.815
cc_140 N_VPB_M1006_b N_X_R23_noxref_pos 7.17606e-19 $X=-0.33 $Y=1.885 $X2=1.82
+ $Y2=1.565
cc_141 N_A_c_145_n N_A_45_443#_M1001_g 0.0209951f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_142 N_A_M1019_g N_A_45_443#_c_238_n 0.0209951f $X=2.6 $Y=2.965 $X2=9.36 $Y2=0
cc_143 N_A_c_141_n N_A_45_443#_c_272_n 0.00436519f $X=0.78 $Y=1.565 $X2=0 $Y2=0
cc_144 N_A_c_141_n N_A_45_443#_c_234_n 0.00386514f $X=0.78 $Y=1.565 $X2=0 $Y2=0
cc_145 N_A_c_146_n N_A_45_443#_c_234_n 0.0206904f $X=0.77 $Y=1.815 $X2=0 $Y2=0
cc_146 A N_A_45_443#_c_234_n 0.0165919f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_147 N_A_M1006_g N_A_45_443#_c_265_n 0.0358157f $X=0.76 $Y=2.965 $X2=0 $Y2=0
cc_148 N_A_c_143_n N_A_45_443#_c_265_n 0.011632f $X=1.57 $Y=1.815 $X2=0 $Y2=0
cc_149 N_A_M1007_g N_A_45_443#_c_265_n 0.0313016f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_150 A N_A_45_443#_c_265_n 0.0678558f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A_M1007_g N_A_45_443#_c_280_n 0.0260651f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_152 N_A_M1019_g N_A_45_443#_c_280_n 0.0467838f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_153 N_A_c_144_n N_A_45_443#_c_282_n 0.00182905f $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_154 N_A_c_145_n N_A_45_443#_c_282_n 0.0126752f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_155 A N_A_45_443#_c_282_n 0.00323676f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_156 N_A_c_147_n N_A_45_443#_c_282_n 0.00406669f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_157 N_A_M1007_g N_A_45_443#_c_286_n 3.42237e-19 $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_158 N_A_M1019_g N_A_45_443#_c_286_n 0.00228752f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_159 N_A_c_147_n N_A_45_443#_c_286_n 0.00975529f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_160 N_A_c_147_n N_A_45_443#_c_235_n 0.0281224f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_161 N_A_M1007_g N_A_45_443#_c_268_n 0.00229199f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_162 N_A_M1019_g N_A_45_443#_c_268_n 0.0148913f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_163 A N_A_45_443#_c_268_n 0.0112571f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A_c_147_n N_A_45_443#_c_268_n 0.00355898f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_165 N_A_c_145_n N_A_45_443#_c_294_n 0.0148072f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_166 A N_A_45_443#_c_294_n 0.00887026f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_167 N_A_c_147_n N_A_45_443#_c_294_n 0.00269586f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_168 A N_A_45_443#_c_297_n 0.0150286f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A_c_147_n N_A_45_443#_c_297_n 0.0133111f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_170 N_A_c_147_n N_A_45_443#_c_237_n 0.0209951f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_171 N_A_M1007_g N_VPWR_c_487_n 0.0103088f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_172 N_A_M1019_g N_VPWR_c_487_n 0.0156302f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_173 N_A_M1019_g N_VPWR_c_501_n 0.00249815f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_174 N_A_M1007_g N_VPWR_c_530_n 7.78697e-19 $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_175 N_A_M1019_g N_VPWR_c_530_n 0.0291392f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_176 N_A_M1006_g N_VPWR_c_514_n 0.0716973f $X=0.76 $Y=2.965 $X2=0 $Y2=0
cc_177 N_A_M1007_g N_VPWR_c_514_n 0.0862897f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_178 N_A_M1019_g N_VPWR_c_514_n 0.00121482f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_179 N_A_M1006_g N_VPWR_c_524_n 0.00951892f $X=0.76 $Y=2.965 $X2=0 $Y2=0
cc_180 N_A_M1007_g N_VPWR_c_524_n 0.010513f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_181 N_A_M1019_g N_VPWR_c_524_n 0.00989232f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_182 N_A_c_144_n N_VGND_c_804_n 0.00367492f $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_183 N_A_c_145_n N_VGND_c_804_n 0.00793008f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_184 N_A_c_141_n N_VGND_c_807_n 0.0572185f $X=0.78 $Y=1.565 $X2=0 $Y2=0
cc_185 N_A_c_143_n N_VGND_c_807_n 0.00914385f $X=1.57 $Y=1.815 $X2=0 $Y2=0
cc_186 N_A_c_144_n N_VGND_c_807_n 0.0624373f $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_187 N_A_c_145_n N_VGND_c_807_n 6.48731e-19 $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_188 A N_VGND_c_807_n 0.0836537f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A_c_144_n N_VGND_c_809_n 4.13084e-19 $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_190 N_A_c_145_n N_VGND_c_809_n 0.0397279f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_191 N_A_c_141_n N_VGND_c_823_n 0.00915616f $X=0.78 $Y=1.565 $X2=0 $Y2=0
cc_192 N_A_c_144_n N_VGND_c_823_n 0.00865748f $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_193 N_A_c_145_n N_VGND_c_823_n 0.00754101f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_194 N_A_c_144_n N_X_c_930_n 5.53867e-19 $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_195 N_A_c_145_n N_X_c_930_n 0.0036162f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_196 N_A_M1019_g N_X_c_930_n 0.00272405f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_197 A N_X_c_930_n 0.00154727f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_198 N_A_c_147_n N_X_c_930_n 0.00612932f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_199 N_A_M1019_g N_X_c_928_n 0.00251614f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_200 N_A_c_147_n N_X_c_928_n 0.00208709f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_201 N_A_c_144_n N_X_R23_noxref_pos 0.00135324f $X=1.82 $Y=1.565 $X2=0.24
+ $Y2=0
cc_202 N_A_M1007_g N_X_R23_noxref_pos 2.48235e-19 $X=1.82 $Y=2.965 $X2=0.24
+ $Y2=0
cc_203 N_A_c_145_n N_X_R23_noxref_pos 0.00243628f $X=2.6 $Y=1.565 $X2=0.24 $Y2=0
cc_204 N_A_M1019_g N_X_R23_noxref_pos 0.00253449f $X=2.6 $Y=2.965 $X2=0.24 $Y2=0
cc_205 A N_X_R23_noxref_pos 0.00218633f $X=2.075 $Y=1.58 $X2=0.24 $Y2=0
cc_206 N_A_c_147_n N_X_R23_noxref_pos 0.0116291f $X=2.6 $Y=1.815 $X2=0.24 $Y2=0
cc_207 N_A_45_443#_c_265_n N_VPWR_M1006_d 0.00539862f $X=2.045 $Y=2.18 $X2=0
+ $Y2=0
cc_208 N_A_45_443#_M1007_s N_VPWR_c_487_n 8.13713e-19 $X=2.07 $Y=2.215 $X2=0
+ $Y2=0
cc_209 N_A_45_443#_c_280_n N_VPWR_c_487_n 0.0314378f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_210 N_A_45_443#_c_238_n N_VPWR_c_490_n 0.00981852f $X=3.38 $Y=2.105 $X2=4.8
+ $Y2=0
cc_211 N_A_45_443#_c_241_n N_VPWR_c_490_n 0.00984257f $X=4.16 $Y=2.105 $X2=4.8
+ $Y2=0
cc_212 N_A_45_443#_c_244_n N_VPWR_c_493_n 0.00984257f $X=4.94 $Y=2.105 $X2=4.8
+ $Y2=0.057
cc_213 N_A_45_443#_c_247_n N_VPWR_c_493_n 0.00984257f $X=5.72 $Y=2.105 $X2=4.8
+ $Y2=0.057
cc_214 N_A_45_443#_c_250_n N_VPWR_c_496_n 0.00984257f $X=6.5 $Y=2.105 $X2=4.8
+ $Y2=0.058
cc_215 N_A_45_443#_c_253_n N_VPWR_c_496_n 0.00984257f $X=7.28 $Y=2.105 $X2=4.8
+ $Y2=0.058
cc_216 N_A_45_443#_c_256_n N_VPWR_c_499_n 7.80614e-19 $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_217 N_A_45_443#_c_259_n N_VPWR_c_499_n 0.014504f $X=8.84 $Y=2.105 $X2=0 $Y2=0
cc_218 N_A_45_443#_c_238_n N_VPWR_c_501_n 0.00656115f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_219 N_A_45_443#_c_241_n N_VPWR_c_504_n 0.00656544f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_220 N_A_45_443#_c_244_n N_VPWR_c_504_n 0.00656544f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_221 N_A_45_443#_c_247_n N_VPWR_c_507_n 0.00656544f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_222 N_A_45_443#_c_250_n N_VPWR_c_507_n 0.00656544f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_223 N_A_45_443#_c_253_n N_VPWR_c_510_n 0.00656544f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_224 N_A_45_443#_c_256_n N_VPWR_c_510_n 0.00656544f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_225 N_A_45_443#_c_238_n N_VPWR_c_530_n 0.0586252f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_226 N_A_45_443#_c_241_n N_VPWR_c_530_n 4.52391e-19 $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_227 N_A_45_443#_c_280_n N_VPWR_c_530_n 0.0866648f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_228 N_A_45_443#_c_235_n N_VPWR_c_530_n 0.0220882f $X=3.295 $Y=1.79 $X2=0
+ $Y2=0
cc_229 N_A_45_443#_c_238_n N_VPWR_c_560_n 4.54877e-19 $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_230 N_A_45_443#_c_241_n N_VPWR_c_560_n 0.0555877f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_231 N_A_45_443#_c_244_n N_VPWR_c_560_n 0.054087f $X=4.94 $Y=2.105 $X2=0 $Y2=0
cc_232 N_A_45_443#_c_247_n N_VPWR_c_560_n 4.54877e-19 $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_233 N_A_45_443#_c_237_n N_VPWR_c_560_n 5.99646e-19 $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_234 N_A_45_443#_c_244_n N_VPWR_c_565_n 4.54877e-19 $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_235 N_A_45_443#_c_247_n N_VPWR_c_565_n 0.0536603f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_236 N_A_45_443#_c_250_n N_VPWR_c_565_n 0.0568798f $X=6.5 $Y=2.105 $X2=0 $Y2=0
cc_237 N_A_45_443#_c_253_n N_VPWR_c_565_n 4.54877e-19 $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_238 N_A_45_443#_c_237_n N_VPWR_c_565_n 5.92537e-19 $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_239 N_A_45_443#_c_250_n N_VPWR_c_570_n 4.54877e-19 $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_240 N_A_45_443#_c_253_n N_VPWR_c_570_n 0.0570434f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_241 N_A_45_443#_c_256_n N_VPWR_c_570_n 0.0569076f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_242 N_A_45_443#_c_259_n N_VPWR_c_570_n 0.0011619f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_243 N_A_45_443#_c_237_n N_VPWR_c_570_n 6.12604e-19 $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_244 N_A_45_443#_c_263_n N_VPWR_c_514_n 0.0817667f $X=0.35 $Y=2.36 $X2=0 $Y2=0
cc_245 N_A_45_443#_c_265_n N_VPWR_c_514_n 0.0847738f $X=2.045 $Y=2.18 $X2=0
+ $Y2=0
cc_246 N_A_45_443#_c_280_n N_VPWR_c_514_n 0.0787997f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_247 N_A_45_443#_c_256_n N_VPWR_c_517_n 0.0098265f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_248 N_A_45_443#_c_259_n N_VPWR_c_517_n 0.0115186f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_249 N_A_45_443#_c_256_n N_VPWR_c_486_n 0.00267747f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_250 N_A_45_443#_c_259_n N_VPWR_c_486_n 0.00803402f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_251 N_A_45_443#_M1006_s N_VPWR_c_524_n 0.00425071f $X=0.225 $Y=2.215 $X2=0
+ $Y2=0
cc_252 N_A_45_443#_c_238_n N_VPWR_c_524_n 0.00914786f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_253 N_A_45_443#_c_241_n N_VPWR_c_524_n 0.00966853f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_254 N_A_45_443#_c_244_n N_VPWR_c_524_n 0.00804425f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_255 N_A_45_443#_c_247_n N_VPWR_c_524_n 0.00803501f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_256 N_A_45_443#_c_250_n N_VPWR_c_524_n 0.00991229f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_257 N_A_45_443#_c_253_n N_VPWR_c_524_n 0.00994001f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_258 N_A_45_443#_c_256_n N_VPWR_c_524_n 0.00804598f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_259 N_A_45_443#_c_259_n N_VPWR_c_524_n 0.014756f $X=8.84 $Y=2.105 $X2=0 $Y2=0
cc_260 N_A_45_443#_c_263_n N_VPWR_c_524_n 0.0196936f $X=0.35 $Y=2.36 $X2=0 $Y2=0
cc_261 N_A_45_443#_c_280_n N_VPWR_c_524_n 0.0205648f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_262 N_A_45_443#_c_238_n N_noxref_6_c_657_n 0.0239099f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_263 N_A_45_443#_c_241_n N_noxref_6_c_657_n 0.0239099f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_264 N_A_45_443#_M1001_g N_noxref_6_c_645_n 0.00442853f $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_265 N_A_45_443#_M1002_g N_noxref_6_c_645_n 0.0044376f $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_266 N_A_45_443#_c_237_n N_noxref_6_c_645_n 0.00438476f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_267 N_A_45_443#_c_241_n N_noxref_6_c_652_n 0.0169508f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_268 N_A_45_443#_c_244_n N_noxref_6_c_652_n 0.0163241f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_269 N_A_45_443#_c_237_n N_noxref_6_c_652_n 0.0780335f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_270 N_A_45_443#_c_244_n N_noxref_6_c_665_n 0.0219493f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_271 N_A_45_443#_c_247_n N_noxref_6_c_665_n 0.0219493f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_272 N_A_45_443#_M1009_g N_noxref_6_c_646_n 0.00506746f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_273 N_A_45_443#_M1013_g N_noxref_6_c_646_n 0.00506746f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_274 N_A_45_443#_c_237_n N_noxref_6_c_646_n 0.00437511f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_275 N_A_45_443#_c_250_n N_noxref_6_c_670_n 0.0256649f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_276 N_A_45_443#_c_253_n N_noxref_6_c_670_n 0.0259143f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_277 N_A_45_443#_M1014_g N_noxref_6_c_647_n 0.00400399f $X=6.5 $Y=1.08 $X2=0
+ $Y2=0
cc_278 N_A_45_443#_M1018_g N_noxref_6_c_647_n 0.00400399f $X=7.28 $Y=1.08 $X2=0
+ $Y2=0
cc_279 N_A_45_443#_c_237_n N_noxref_6_c_647_n 0.00455707f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_280 N_A_45_443#_c_253_n N_noxref_6_c_653_n 0.018715f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_281 N_A_45_443#_c_256_n N_noxref_6_c_653_n 0.0186574f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_282 N_A_45_443#_c_237_n N_noxref_6_c_653_n 0.0821832f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_283 N_A_45_443#_c_256_n N_noxref_6_c_678_n 0.00796164f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_284 N_A_45_443#_c_259_n N_noxref_6_c_678_n 0.0261864f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_285 N_A_45_443#_c_256_n N_noxref_6_c_680_n 0.0174543f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_286 N_A_45_443#_c_259_n N_noxref_6_c_680_n 0.0363022f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_287 N_A_45_443#_M1020_g N_noxref_6_c_648_n 0.00569856f $X=8.06 $Y=1.08 $X2=0
+ $Y2=0
cc_288 N_A_45_443#_M1021_g N_noxref_6_c_648_n 0.045504f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_289 N_A_45_443#_c_237_n N_noxref_6_c_648_n 0.00541261f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_290 N_A_45_443#_c_238_n N_noxref_6_c_685_n 0.00494888f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_291 N_A_45_443#_c_241_n N_noxref_6_c_685_n 0.00141551f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_292 N_A_45_443#_c_235_n N_noxref_6_c_685_n 0.0173736f $X=3.295 $Y=1.79 $X2=0
+ $Y2=0
cc_293 N_A_45_443#_c_237_n N_noxref_6_c_685_n 0.0312834f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_294 N_A_45_443#_c_244_n N_noxref_6_c_689_n 0.00141551f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_295 N_A_45_443#_c_247_n N_noxref_6_c_689_n 0.00141551f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_296 N_A_45_443#_c_237_n N_noxref_6_c_689_n 0.0224144f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_297 N_A_45_443#_c_247_n N_noxref_6_c_654_n 0.0160507f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_298 N_A_45_443#_c_250_n N_noxref_6_c_654_n 0.0185061f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_299 N_A_45_443#_c_237_n N_noxref_6_c_654_n 0.0789792f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_300 N_A_45_443#_c_250_n N_noxref_6_c_695_n 0.00141551f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_301 N_A_45_443#_c_253_n N_noxref_6_c_695_n 0.00141551f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_302 N_A_45_443#_c_237_n N_noxref_6_c_695_n 0.0236345f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_303 N_A_45_443#_c_256_n N_noxref_6_c_698_n 0.00141551f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_304 N_A_45_443#_c_259_n N_noxref_6_c_698_n 0.00911503f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_305 N_A_45_443#_c_237_n N_noxref_6_c_698_n 0.0578292f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_306 N_A_45_443#_M1002_g N_noxref_6_c_649_n 6.18587e-19 $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_307 N_A_45_443#_c_241_n N_noxref_6_c_649_n 6.9098e-19 $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_308 N_A_45_443#_M1009_g N_noxref_6_c_649_n 0.0040183f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_309 N_A_45_443#_c_244_n N_noxref_6_c_649_n 0.00648623f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_310 N_A_45_443#_M1013_g N_noxref_6_c_649_n 0.00583477f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_311 N_A_45_443#_c_247_n N_noxref_6_c_649_n 0.00206235f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_312 N_A_45_443#_M1014_g N_noxref_6_c_649_n 9.74028e-19 $X=6.5 $Y=1.08 $X2=0
+ $Y2=0
cc_313 N_A_45_443#_c_250_n N_noxref_6_c_649_n 0.00108806f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_314 N_A_45_443#_c_237_n N_noxref_6_c_649_n 7.46635e-19 $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_315 N_A_45_443#_M1002_g N_noxref_6_R23_noxref_neg 2.08344e-19 $X=4.16 $Y=1.08
+ $X2=0 $Y2=0
cc_316 N_A_45_443#_c_241_n N_noxref_6_R23_noxref_neg 3.03057e-19 $X=4.16
+ $Y=2.105 $X2=0 $Y2=0
cc_317 N_A_45_443#_M1009_g N_noxref_6_R23_noxref_neg 4.18085e-19 $X=4.94 $Y=1.08
+ $X2=0 $Y2=0
cc_318 N_A_45_443#_c_244_n N_noxref_6_R23_noxref_neg 0.00178224f $X=4.94
+ $Y=2.105 $X2=0 $Y2=0
cc_319 N_A_45_443#_M1013_g N_noxref_6_R23_noxref_neg 2.09742e-19 $X=5.72 $Y=1.08
+ $X2=0 $Y2=0
cc_320 N_A_45_443#_c_247_n N_noxref_6_R23_noxref_neg 0.00118463f $X=5.72
+ $Y=2.105 $X2=0 $Y2=0
cc_321 N_A_45_443#_M1014_g N_noxref_6_R23_noxref_neg 0.00271381f $X=6.5 $Y=1.08
+ $X2=0 $Y2=0
cc_322 N_A_45_443#_c_250_n N_noxref_6_R23_noxref_neg 0.00340122f $X=6.5 $Y=2.105
+ $X2=0 $Y2=0
cc_323 N_A_45_443#_c_237_n N_noxref_6_R23_noxref_neg 5.74971e-19 $X=8.84
+ $Y=1.855 $X2=0 $Y2=0
cc_324 N_A_45_443#_c_417_p N_VGND_c_804_n 0.0122346f $X=2.21 $Y=0.895 $X2=0
+ $Y2=0
cc_325 N_A_45_443#_M1021_g N_VGND_c_805_n 0.00759687f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_326 N_A_45_443#_c_272_n N_VGND_c_807_n 0.0377885f $X=0.37 $Y=0.97 $X2=0 $Y2=0
cc_327 N_A_45_443#_M1001_g N_VGND_c_809_n 0.0545773f $X=3.38 $Y=1.08 $X2=0 $Y2=0
cc_328 N_A_45_443#_M1002_g N_VGND_c_809_n 0.00107285f $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_329 N_A_45_443#_c_282_n N_VGND_c_809_n 0.00345517f $X=2.51 $Y=1.625 $X2=0
+ $Y2=0
cc_330 N_A_45_443#_c_235_n N_VGND_c_809_n 0.0459241f $X=3.295 $Y=1.79 $X2=0
+ $Y2=0
cc_331 N_A_45_443#_c_294_n N_VGND_c_809_n 0.0137366f $X=2.51 $Y=1.315 $X2=0
+ $Y2=0
cc_332 N_A_45_443#_M1001_g N_VGND_c_811_n 0.00328808f $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_333 N_A_45_443#_M1002_g N_VGND_c_811_n 0.00328808f $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_334 N_A_45_443#_M1001_g N_VGND_c_813_n 0.00107181f $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_335 N_A_45_443#_M1002_g N_VGND_c_813_n 0.0516357f $X=4.16 $Y=1.08 $X2=0 $Y2=0
cc_336 N_A_45_443#_M1009_g N_VGND_c_813_n 0.0508722f $X=4.94 $Y=1.08 $X2=0 $Y2=0
cc_337 N_A_45_443#_M1013_g N_VGND_c_813_n 0.00177985f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_338 N_A_45_443#_c_237_n N_VGND_c_813_n 0.00249165f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_339 N_A_45_443#_M1009_g N_VGND_c_814_n 0.00328808f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_340 N_A_45_443#_M1013_g N_VGND_c_814_n 0.00328808f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_341 N_A_45_443#_M1009_g N_VGND_c_815_n 0.00177985f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_342 N_A_45_443#_M1013_g N_VGND_c_815_n 0.0508722f $X=5.72 $Y=1.08 $X2=0 $Y2=0
cc_343 N_A_45_443#_M1014_g N_VGND_c_815_n 0.052403f $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_344 N_A_45_443#_M1018_g N_VGND_c_815_n 9.10934e-19 $X=7.28 $Y=1.08 $X2=0
+ $Y2=0
cc_345 N_A_45_443#_c_237_n N_VGND_c_815_n 0.00244934f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_346 N_A_45_443#_M1014_g N_VGND_c_816_n 0.00328808f $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_347 N_A_45_443#_M1018_g N_VGND_c_816_n 0.00328808f $X=7.28 $Y=1.08 $X2=0
+ $Y2=0
cc_348 N_A_45_443#_M1014_g N_VGND_c_817_n 9.10934e-19 $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_349 N_A_45_443#_M1018_g N_VGND_c_817_n 0.0525668f $X=7.28 $Y=1.08 $X2=0 $Y2=0
cc_350 N_A_45_443#_M1020_g N_VGND_c_817_n 0.0564921f $X=8.06 $Y=1.08 $X2=0 $Y2=0
cc_351 N_A_45_443#_M1021_g N_VGND_c_817_n 0.00263084f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_352 N_A_45_443#_c_237_n N_VGND_c_817_n 0.00257674f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_353 N_A_45_443#_M1020_g N_VGND_c_818_n 0.00520463f $X=8.06 $Y=1.08 $X2=0
+ $Y2=0
cc_354 N_A_45_443#_M1021_g N_VGND_c_818_n 0.00966456f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_355 N_A_45_443#_M1021_g N_VGND_c_819_n 0.00617584f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_356 N_A_45_443#_M1020_g N_VGND_c_821_n 0.00209553f $X=8.06 $Y=1.08 $X2=0
+ $Y2=0
cc_357 N_A_45_443#_M1021_g N_VGND_c_821_n 0.00725856f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_358 N_A_45_443#_M1001_g N_VGND_c_823_n 0.00754797f $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_359 N_A_45_443#_M1002_g N_VGND_c_823_n 0.00786843f $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_360 N_A_45_443#_M1009_g N_VGND_c_823_n 0.00676762f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_361 N_A_45_443#_M1013_g N_VGND_c_823_n 0.00676762f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_362 N_A_45_443#_M1014_g N_VGND_c_823_n 0.00808151f $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_363 N_A_45_443#_M1018_g N_VGND_c_823_n 0.00808151f $X=7.28 $Y=1.08 $X2=0
+ $Y2=0
cc_364 N_A_45_443#_M1020_g N_VGND_c_823_n 0.00676762f $X=8.06 $Y=1.08 $X2=0
+ $Y2=0
cc_365 N_A_45_443#_M1021_g N_VGND_c_823_n 0.0228805f $X=8.84 $Y=1.08 $X2=0 $Y2=0
cc_366 N_A_45_443#_c_272_n N_VGND_c_823_n 0.0118041f $X=0.37 $Y=0.97 $X2=0 $Y2=0
cc_367 N_A_45_443#_c_417_p N_VGND_c_823_n 0.00689067f $X=2.21 $Y=0.895 $X2=0
+ $Y2=0
cc_368 N_A_45_443#_c_294_n N_VGND_c_823_n 0.00762664f $X=2.51 $Y=1.315 $X2=0
+ $Y2=0
cc_369 N_A_45_443#_M1001_g N_X_c_930_n 0.00310982f $X=3.38 $Y=1.08 $X2=0 $Y2=0
cc_370 N_A_45_443#_c_238_n N_X_c_930_n 0.00688764f $X=3.38 $Y=2.105 $X2=0 $Y2=0
cc_371 N_A_45_443#_c_280_n N_X_c_930_n 0.00748404f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_372 N_A_45_443#_c_282_n N_X_c_930_n 0.00319717f $X=2.51 $Y=1.625 $X2=0 $Y2=0
cc_373 N_A_45_443#_c_286_n N_X_c_930_n 0.00110944f $X=2.51 $Y=2.095 $X2=0 $Y2=0
cc_374 N_A_45_443#_c_235_n N_X_c_930_n 0.00256495f $X=3.295 $Y=1.79 $X2=0 $Y2=0
cc_375 N_A_45_443#_c_268_n N_X_c_930_n 0.00343251f $X=2.32 $Y=2.18 $X2=0 $Y2=0
cc_376 N_A_45_443#_c_294_n N_X_c_930_n 0.00102022f $X=2.51 $Y=1.315 $X2=0 $Y2=0
cc_377 N_A_45_443#_c_297_n N_X_c_930_n 3.57797e-19 $X=2.51 $Y=1.79 $X2=0 $Y2=0
cc_378 N_A_45_443#_c_237_n N_X_c_930_n 0.00328139f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_379 N_A_45_443#_c_238_n N_X_c_928_n 0.00775937f $X=3.38 $Y=2.105 $X2=0 $Y2=0
cc_380 N_A_45_443#_c_286_n N_X_c_928_n 0.00173712f $X=2.51 $Y=2.095 $X2=0 $Y2=0
cc_381 N_A_45_443#_c_235_n N_X_c_928_n 0.010945f $X=3.295 $Y=1.79 $X2=0 $Y2=0
cc_382 N_A_45_443#_c_268_n N_X_c_928_n 0.0015254f $X=2.32 $Y=2.18 $X2=0 $Y2=0
cc_383 N_A_45_443#_c_237_n N_X_c_928_n 0.00617226f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_384 N_A_45_443#_M1008_d N_X_R23_noxref_pos 0.00135986f $X=2.07 $Y=0.705
+ $X2=0.24 $Y2=0
cc_385 N_A_45_443#_M1001_g N_X_R23_noxref_pos 0.0021287f $X=3.38 $Y=1.08
+ $X2=0.24 $Y2=0
cc_386 N_A_45_443#_c_238_n N_X_R23_noxref_pos 0.00253449f $X=3.38 $Y=2.105
+ $X2=0.24 $Y2=0
cc_387 N_A_45_443#_M1002_g N_X_R23_noxref_pos 0.0021287f $X=4.16 $Y=1.08
+ $X2=0.24 $Y2=0
cc_388 N_A_45_443#_c_241_n N_X_R23_noxref_pos 0.00253449f $X=4.16 $Y=2.105
+ $X2=0.24 $Y2=0
cc_389 N_A_45_443#_c_280_n N_X_R23_noxref_pos 0.0142404f $X=2.21 $Y=2.34
+ $X2=0.24 $Y2=0
cc_390 N_A_45_443#_c_236_n N_X_R23_noxref_pos 8.95427e-19 $X=0.35 $Y=1.475
+ $X2=0.24 $Y2=0
cc_391 N_A_45_443#_c_268_n N_X_R23_noxref_pos 0.00420439f $X=2.32 $Y=2.18
+ $X2=0.24 $Y2=0
cc_392 N_A_45_443#_c_294_n N_X_R23_noxref_pos 0.00784726f $X=2.51 $Y=1.315
+ $X2=0.24 $Y2=0
cc_393 N_VPWR_c_490_n N_noxref_6_M1000_d 8.28689e-19 $X=4.105 $Y=3.71 $X2=-0.33
+ $Y2=-0.365
cc_394 N_VPWR_c_493_n N_noxref_6_M1005_d 8.28689e-19 $X=5.665 $Y=3.71 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_496_n N_noxref_6_M1011_d 8.28689e-19 $X=7.225 $Y=3.71 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_517_n N_noxref_6_M1016_d 8.28689e-19 $X=8.905 $Y=3.635 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_490_n N_noxref_6_c_657_n 0.0178796f $X=4.105 $Y=3.71 $X2=0 $Y2=0
cc_398 N_VPWR_c_530_n N_noxref_6_c_657_n 0.0838628f $X=2.99 $Y=2.55 $X2=0 $Y2=0
cc_399 N_VPWR_c_560_n N_noxref_6_c_657_n 0.0840852f $X=4.55 $Y=2.55 $X2=0 $Y2=0
cc_400 N_VPWR_c_524_n N_noxref_6_c_657_n 0.01238f $X=9.415 $Y=3.63 $X2=0 $Y2=0
cc_401 N_VPWR_c_560_n N_noxref_6_c_652_n 0.0692707f $X=4.55 $Y=2.55 $X2=0 $Y2=0
cc_402 N_VPWR_c_493_n N_noxref_6_c_665_n 0.0178796f $X=5.665 $Y=3.71 $X2=0 $Y2=0
cc_403 N_VPWR_c_560_n N_noxref_6_c_665_n 0.0839242f $X=4.55 $Y=2.55 $X2=0 $Y2=0
cc_404 N_VPWR_c_565_n N_noxref_6_c_665_n 0.0838049f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_405 N_VPWR_c_524_n N_noxref_6_c_665_n 0.0122121f $X=9.415 $Y=3.63 $X2=0 $Y2=0
cc_406 N_VPWR_c_496_n N_noxref_6_c_670_n 0.0178796f $X=7.225 $Y=3.71 $X2=0 $Y2=0
cc_407 N_VPWR_c_565_n N_noxref_6_c_670_n 0.0842143f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_408 N_VPWR_c_570_n N_noxref_6_c_670_n 0.0842143f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_409 N_VPWR_c_486_n N_noxref_6_c_670_n 0.0010411f $X=9.76 $Y=3.635 $X2=0 $Y2=0
cc_410 N_VPWR_c_524_n N_noxref_6_c_670_n 0.01238f $X=9.415 $Y=3.63 $X2=0 $Y2=0
cc_411 N_VPWR_c_570_n N_noxref_6_c_653_n 0.0676163f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_412 N_VPWR_c_486_n N_noxref_6_c_653_n 0.00189868f $X=9.76 $Y=3.635 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_499_n N_noxref_6_c_678_n 0.00310535f $X=9.32 $Y=3.475 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_500_n N_noxref_6_c_678_n 0.0279072f $X=9.23 $Y=2.55 $X2=0 $Y2=0
cc_415 N_VPWR_c_570_n N_noxref_6_c_678_n 0.045569f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_416 N_VPWR_c_517_n N_noxref_6_c_678_n 0.0308132f $X=8.905 $Y=3.635 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_486_n N_noxref_6_c_678_n 0.00468236f $X=9.76 $Y=3.635 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_524_n N_noxref_6_c_678_n 0.0228407f $X=9.415 $Y=3.63 $X2=0 $Y2=0
cc_419 N_VPWR_c_500_n N_noxref_6_c_680_n 0.0222528f $X=9.23 $Y=2.55 $X2=0 $Y2=0
cc_420 N_VPWR_c_570_n N_noxref_6_c_680_n 0.0422153f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_421 N_VPWR_c_486_n N_noxref_6_c_680_n 0.00765982f $X=9.76 $Y=3.635 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_565_n N_noxref_6_c_654_n 0.0689643f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_423 N_VPWR_M1010_s N_noxref_6_c_649_n 0.00192727f $X=5.97 $Y=2.215 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_560_n N_noxref_6_c_649_n 0.00162743f $X=4.55 $Y=2.55 $X2=0 $Y2=0
cc_425 N_VPWR_c_565_n N_noxref_6_c_649_n 0.0105841f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_426 N_VPWR_c_524_n N_noxref_6_c_649_n 0.0129114f $X=9.415 $Y=3.63 $X2=0 $Y2=0
cc_427 N_VPWR_c_565_n N_noxref_6_c_753_n 0.00364733f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_428 N_VPWR_c_560_n N_noxref_6_R23_noxref_neg 0.0198058f $X=4.55 $Y=2.55 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_565_n N_noxref_6_R23_noxref_neg 0.0122645f $X=6.11 $Y=2.55 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_486_n N_noxref_6_R23_noxref_neg 0.119287f $X=9.76 $Y=3.635 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_524_n N_noxref_6_R23_noxref_neg 0.0409695f $X=9.415 $Y=3.63
+ $X2=0 $Y2=0
cc_432 N_VPWR_c_565_n N_noxref_6_c_758_n 0.00779455f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_433 N_VPWR_c_565_n N_noxref_6_c_759_n 0.00483754f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_434 N_VPWR_c_486_n N_VGND_c_805_n 0.00250322f $X=9.76 $Y=3.635 $X2=0 $Y2=0
cc_435 N_VPWR_c_500_n N_VGND_c_821_n 0.00260627f $X=9.23 $Y=2.55 $X2=0 $Y2=0
cc_436 N_VPWR_c_486_n N_VGND_c_821_n 0.218481f $X=9.76 $Y=3.635 $X2=0 $Y2=0
cc_437 N_VPWR_c_530_n N_X_c_930_n 0.0108923f $X=2.99 $Y=2.55 $X2=0 $Y2=0
cc_438 N_VPWR_c_514_n N_X_c_930_n 9.22025e-19 $X=1.15 $Y=2.55 $X2=0 $Y2=0
cc_439 N_VPWR_c_524_n N_X_c_930_n 0.0162902f $X=9.415 $Y=3.63 $X2=0 $Y2=0
cc_440 N_VPWR_c_530_n N_X_c_928_n 0.00579934f $X=2.99 $Y=2.55 $X2=0 $Y2=0
cc_441 N_VPWR_c_530_n N_X_R23_noxref_pos 0.0110619f $X=2.99 $Y=2.55 $X2=0.24
+ $Y2=0
cc_442 N_VPWR_c_560_n N_X_R23_noxref_pos 0.00150025f $X=4.55 $Y=2.55 $X2=0.24
+ $Y2=0
cc_443 N_VPWR_c_514_n N_X_R23_noxref_pos 0.00127107f $X=1.15 $Y=2.55 $X2=0.24
+ $Y2=0
cc_444 N_VPWR_c_524_n N_X_R23_noxref_pos 0.0293367f $X=9.415 $Y=3.63 $X2=0.24
+ $Y2=0
cc_445 N_noxref_6_c_649_n N_VGND_M1013_s 0.00196128f $X=5.6 $Y=2.035 $X2=0 $Y2=0
cc_446 N_noxref_6_c_648_n N_VGND_c_805_n 0.0353446f $X=8.45 $Y=0.97 $X2=0 $Y2=0
cc_447 N_noxref_6_c_645_n N_VGND_c_809_n 0.0310184f $X=3.77 $Y=0.97 $X2=0 $Y2=0
cc_448 N_noxref_6_R23_noxref_neg N_VGND_c_809_n 6.9774e-19 $X=4.26 $Y=2.035
+ $X2=0 $Y2=0
cc_449 N_noxref_6_c_645_n N_VGND_c_811_n 0.0086879f $X=3.77 $Y=0.97 $X2=0 $Y2=0
cc_450 N_noxref_6_c_645_n N_VGND_c_813_n 0.030957f $X=3.77 $Y=0.97 $X2=0 $Y2=0
cc_451 N_noxref_6_c_652_n N_VGND_c_813_n 0.0772082f $X=5.165 $Y=1.915 $X2=0
+ $Y2=0
cc_452 N_noxref_6_c_646_n N_VGND_c_813_n 0.0392681f $X=5.33 $Y=0.97 $X2=0 $Y2=0
cc_453 N_noxref_6_c_649_n N_VGND_c_813_n 3.09146e-19 $X=5.6 $Y=2.035 $X2=0 $Y2=0
cc_454 N_noxref_6_R23_noxref_neg N_VGND_c_813_n 0.0197926f $X=4.26 $Y=2.035
+ $X2=0 $Y2=0
cc_455 N_noxref_6_c_646_n N_VGND_c_814_n 0.0110067f $X=5.33 $Y=0.97 $X2=0 $Y2=0
cc_456 N_noxref_6_c_646_n N_VGND_c_815_n 0.0392681f $X=5.33 $Y=0.97 $X2=0 $Y2=0
cc_457 N_noxref_6_c_654_n N_VGND_c_815_n 0.0772623f $X=6.725 $Y=1.915 $X2=0
+ $Y2=0
cc_458 N_noxref_6_c_649_n N_VGND_c_815_n 0.00438917f $X=5.6 $Y=2.035 $X2=0 $Y2=0
cc_459 N_noxref_6_c_753_n N_VGND_c_815_n 0.00355428f $X=6.025 $Y=2.035 $X2=0
+ $Y2=0
cc_460 N_noxref_6_R23_noxref_neg N_VGND_c_815_n 0.00946502f $X=4.26 $Y=2.035
+ $X2=0 $Y2=0
cc_461 N_noxref_6_c_758_n N_VGND_c_815_n 0.00580423f $X=6.05 $Y=2.035 $X2=0
+ $Y2=0
cc_462 N_noxref_6_c_759_n N_VGND_c_815_n 0.00431302f $X=6.025 $Y=2.035 $X2=0
+ $Y2=0
cc_463 N_noxref_6_c_647_n N_VGND_c_816_n 0.0086879f $X=6.89 $Y=0.97 $X2=0 $Y2=0
cc_464 N_noxref_6_c_653_n N_VGND_c_817_n 0.0757221f $X=8.285 $Y=1.915 $X2=0
+ $Y2=0
cc_465 N_noxref_6_c_648_n N_VGND_c_817_n 0.0363619f $X=8.45 $Y=0.97 $X2=0 $Y2=0
cc_466 N_noxref_6_R23_noxref_neg N_VGND_c_817_n 6.65414e-19 $X=4.26 $Y=2.035
+ $X2=0 $Y2=0
cc_467 N_noxref_6_c_648_n N_VGND_c_818_n 0.0324116f $X=8.45 $Y=0.97 $X2=0 $Y2=0
cc_468 N_noxref_6_M1020_d N_VGND_c_821_n 2.92037e-19 $X=8.31 $Y=0.705 $X2=0
+ $Y2=0
cc_469 N_noxref_6_c_647_n N_VGND_c_821_n 7.24629e-19 $X=6.89 $Y=0.97 $X2=0 $Y2=0
cc_470 N_noxref_6_c_653_n N_VGND_c_821_n 0.00163768f $X=8.285 $Y=1.915 $X2=0
+ $Y2=0
cc_471 N_noxref_6_c_648_n N_VGND_c_821_n 0.0108355f $X=8.45 $Y=0.97 $X2=0 $Y2=0
cc_472 N_noxref_6_c_698_n N_VGND_c_821_n 6.16682e-19 $X=8.625 $Y=1.915 $X2=0
+ $Y2=0
cc_473 N_noxref_6_R23_noxref_neg N_VGND_c_821_n 0.119314f $X=4.26 $Y=2.035 $X2=0
+ $Y2=0
cc_474 N_noxref_6_c_645_n N_VGND_c_823_n 0.00668507f $X=3.77 $Y=0.97 $X2=0 $Y2=0
cc_475 N_noxref_6_c_646_n N_VGND_c_823_n 0.00646874f $X=5.33 $Y=0.97 $X2=0 $Y2=0
cc_476 N_noxref_6_c_647_n N_VGND_c_823_n 0.00668507f $X=6.89 $Y=0.97 $X2=0 $Y2=0
cc_477 N_noxref_6_c_648_n N_VGND_c_823_n 0.0175488f $X=8.45 $Y=0.97 $X2=0 $Y2=0
cc_478 N_noxref_6_c_649_n N_VGND_c_823_n 0.0144641f $X=5.6 $Y=2.035 $X2=0 $Y2=0
cc_479 N_noxref_6_R23_noxref_neg N_VGND_c_823_n 0.0464145f $X=4.26 $Y=2.035
+ $X2=0 $Y2=0
cc_480 N_noxref_6_c_657_n N_X_c_930_n 0.00329012f $X=3.77 $Y=2.34 $X2=0 $Y2=0
cc_481 N_noxref_6_c_645_n N_X_c_930_n 0.00173013f $X=3.77 $Y=0.97 $X2=0 $Y2=0
cc_482 N_noxref_6_c_685_n N_X_c_930_n 0.00185251f $X=3.605 $Y=1.955 $X2=0 $Y2=0
cc_483 N_noxref_6_c_685_n N_X_c_928_n 0.00987178f $X=3.605 $Y=1.955 $X2=0 $Y2=0
cc_484 N_noxref_6_M1001_d N_X_R23_noxref_pos 0.00135817f $X=3.63 $Y=0.705
+ $X2=0.24 $Y2=0
cc_485 N_noxref_6_c_657_n N_X_R23_noxref_pos 0.00725409f $X=3.77 $Y=2.34
+ $X2=0.24 $Y2=0
cc_486 N_noxref_6_c_645_n N_X_R23_noxref_pos 0.00554638f $X=3.77 $Y=0.97
+ $X2=0.24 $Y2=0
cc_487 N_noxref_6_c_652_n N_X_R23_noxref_pos 8.93242e-19 $X=5.165 $Y=1.915
+ $X2=0.24 $Y2=0
cc_488 N_noxref_6_c_685_n N_X_R23_noxref_pos 9.90742e-19 $X=3.605 $Y=1.955
+ $X2=0.24 $Y2=0
cc_489 N_VGND_c_809_n N_X_c_930_n 0.00859918f $X=2.69 $Y=0.465 $X2=0 $Y2=0
cc_490 N_VGND_c_823_n N_X_c_930_n 0.01616f $X=9.415 $Y=0.44 $X2=0 $Y2=0
cc_491 N_VGND_c_809_n N_X_c_928_n 0.00441639f $X=2.69 $Y=0.465 $X2=0 $Y2=0
cc_492 N_VGND_c_807_n N_X_R23_noxref_pos 4.93623e-19 $X=1.925 $Y=0.882 $X2=0.24
+ $Y2=0
cc_493 N_VGND_c_809_n N_X_R23_noxref_pos 0.013732f $X=2.69 $Y=0.465 $X2=0.24
+ $Y2=0
cc_494 N_VGND_c_813_n N_X_R23_noxref_pos 0.00220478f $X=5.055 $Y=0.912 $X2=0.24
+ $Y2=0
cc_495 N_VGND_c_823_n N_X_R23_noxref_pos 0.0301598f $X=9.415 $Y=0.44 $X2=0.24
+ $Y2=0
