* File: sky130_fd_sc_hvl__a21oi_1.pxi.spice
* Created: Fri Aug 28 09:32:15 2020
* 
x_PM_SKY130_FD_SC_HVL__A21OI_1%VNB N_VNB_M1000_b VNB N_VNB_c_8_p VNB
+ PM_SKY130_FD_SC_HVL__A21OI_1%VNB
x_PM_SKY130_FD_SC_HVL__A21OI_1%VPB N_VPB_M1003_b VPB N_VPB_c_23_p VPB
+ PM_SKY130_FD_SC_HVL__A21OI_1%VPB
x_PM_SKY130_FD_SC_HVL__A21OI_1%A2 N_A2_M1003_g N_A2_M1000_g A2 A2 A2 N_A2_c_51_n
+ PM_SKY130_FD_SC_HVL__A21OI_1%A2
x_PM_SKY130_FD_SC_HVL__A21OI_1%A1 A1 N_A1_M1004_g N_A1_M1005_g
+ PM_SKY130_FD_SC_HVL__A21OI_1%A1
x_PM_SKY130_FD_SC_HVL__A21OI_1%B1 N_B1_M1001_g N_B1_M1002_g B1 B1 B1 B1
+ N_B1_c_98_n N_B1_c_107_n N_B1_c_99_n N_B1_c_102_n
+ PM_SKY130_FD_SC_HVL__A21OI_1%B1
x_PM_SKY130_FD_SC_HVL__A21OI_1%A_56_443# N_A_56_443#_M1003_s N_A_56_443#_M1005_d
+ N_A_56_443#_c_126_n N_A_56_443#_c_129_n N_A_56_443#_c_130_n
+ N_A_56_443#_c_131_n PM_SKY130_FD_SC_HVL__A21OI_1%A_56_443#
x_PM_SKY130_FD_SC_HVL__A21OI_1%VPWR N_VPWR_M1003_d VPWR N_VPWR_c_155_n
+ N_VPWR_c_158_n PM_SKY130_FD_SC_HVL__A21OI_1%VPWR
x_PM_SKY130_FD_SC_HVL__A21OI_1%Y N_Y_M1004_d N_Y_M1001_d N_Y_c_177_n N_Y_c_179_n
+ N_Y_c_180_n Y Y Y Y Y N_Y_c_181_n Y PM_SKY130_FD_SC_HVL__A21OI_1%Y
x_PM_SKY130_FD_SC_HVL__A21OI_1%VGND N_VGND_M1000_s N_VGND_M1002_d VGND
+ N_VGND_c_206_n N_VGND_c_208_n N_VGND_c_210_n PM_SKY130_FD_SC_HVL__A21OI_1%VGND
cc_1 N_VNB_M1000_b N_A2_M1000_g 0.0432009f $X=-0.33 $Y=-0.265 $X2=1.105 $Y2=0.91
cc_2 N_VNB_M1000_b A2 0.0295357f $X=-0.33 $Y=-0.265 $X2=1.115 $Y2=1.58
cc_3 N_VNB_M1000_b N_A2_c_51_n 0.074207f $X=-0.33 $Y=-0.265 $X2=1.105 $Y2=1.75
cc_4 N_VNB_M1000_b A1 0.00170292f $X=-0.33 $Y=-0.265 $X2=0.815 $Y2=2.085
cc_5 N_VNB_M1000_b N_A1_M1004_g 0.0800036f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_M1000_b N_B1_c_98_n 0.0567369f $X=-0.33 $Y=-0.265 $X2=0.75 $Y2=1.625
cc_7 N_VNB_M1000_b N_B1_c_99_n 0.0482022f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_8 N_VNB_c_8_p N_B1_c_99_n 0.00107521f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_9 N_VNB_M1000_b N_Y_c_177_n 0.010179f $X=-0.33 $Y=-0.265 $X2=0.155 $Y2=1.58
cc_10 N_VNB_c_8_p N_Y_c_177_n 6.32535e-19 $X=0.24 $Y=0 $X2=0.155 $Y2=1.58
cc_11 N_VNB_M1000_b N_Y_c_179_n 0.00148584f $X=-0.33 $Y=-0.265 $X2=1.115
+ $Y2=1.58
cc_12 N_VNB_M1000_b N_Y_c_180_n 0.00452301f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_13 N_VNB_M1000_b N_Y_c_181_n 0.0100524f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_14 N_VNB_M1000_b Y 0.0130024f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_15 N_VNB_M1000_b N_VGND_c_206_n 0.131643f $X=-0.33 $Y=-0.265 $X2=0.75
+ $Y2=1.625
cc_16 N_VNB_c_8_p N_VGND_c_206_n 0.00484573f $X=0.24 $Y=0 $X2=0.75 $Y2=1.625
cc_17 N_VNB_M1000_b N_VGND_c_208_n 0.0620116f $X=-0.33 $Y=-0.265 $X2=1.105
+ $Y2=1.75
cc_18 N_VNB_c_8_p N_VGND_c_208_n 0.00166879f $X=0.24 $Y=0 $X2=1.105 $Y2=1.75
cc_19 N_VNB_M1000_b N_VGND_c_210_n 0.0779957f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_20 N_VNB_c_8_p N_VGND_c_210_n 0.359258f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_21 N_VPB_M1003_b N_A2_M1003_g 0.0410315f $X=-0.33 $Y=1.885 $X2=0.815
+ $Y2=2.965
cc_22 VPB N_A2_M1003_g 0.00970178f $X=0 $Y=3.955 $X2=0.815 $Y2=2.965
cc_23 N_VPB_c_23_p N_A2_M1003_g 0.0152133f $X=3.12 $Y=4.07 $X2=0.815 $Y2=2.965
cc_24 N_VPB_M1003_b N_A2_c_51_n 0.0343323f $X=-0.33 $Y=1.885 $X2=1.105 $Y2=1.75
cc_25 N_VPB_M1003_b N_A1_M1004_g 0.0532918f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_26 VPB N_A1_M1004_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_27 N_VPB_c_23_p N_A1_M1004_g 0.0152133f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_28 N_VPB_M1003_b N_B1_c_98_n 0.0292346f $X=-0.33 $Y=1.885 $X2=0.75 $Y2=1.625
cc_29 N_VPB_M1003_b N_B1_c_102_n 0.0373173f $X=-0.33 $Y=1.885 $X2=0.815 $Y2=1.75
cc_30 VPB N_B1_c_102_n 0.00970178f $X=0 $Y=3.955 $X2=0.815 $Y2=1.75
cc_31 N_VPB_c_23_p N_B1_c_102_n 0.0196751f $X=3.12 $Y=4.07 $X2=0.815 $Y2=1.75
cc_32 N_VPB_M1003_b N_A_56_443#_c_126_n 0.0566623f $X=-0.33 $Y=1.885 $X2=0.155
+ $Y2=1.58
cc_33 VPB N_A_56_443#_c_126_n 7.60114e-19 $X=0 $Y=3.955 $X2=0.155 $Y2=1.58
cc_34 N_VPB_c_23_p N_A_56_443#_c_126_n 0.0131049f $X=3.12 $Y=4.07 $X2=0.155
+ $Y2=1.58
cc_35 N_VPB_M1003_b N_A_56_443#_c_129_n 0.0202971f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_36 N_VPB_M1003_b N_A_56_443#_c_130_n 0.0101035f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_37 N_VPB_M1003_b N_A_56_443#_c_131_n 0.00351534f $X=-0.33 $Y=1.885 $X2=0.75
+ $Y2=1.625
cc_38 VPB N_A_56_443#_c_131_n 5.14916e-19 $X=0 $Y=3.955 $X2=0.75 $Y2=1.625
cc_39 N_VPB_c_23_p N_A_56_443#_c_131_n 0.00887752f $X=3.12 $Y=4.07 $X2=0.75
+ $Y2=1.625
cc_40 N_VPB_M1003_b N_VPWR_c_155_n 0.00243985f $X=-0.33 $Y=1.885 $X2=1.105
+ $Y2=0.91
cc_41 VPB N_VPWR_c_155_n 0.00512219f $X=0 $Y=3.955 $X2=1.105 $Y2=0.91
cc_42 N_VPB_c_23_p N_VPWR_c_155_n 0.0629871f $X=3.12 $Y=4.07 $X2=1.105 $Y2=0.91
cc_43 N_VPB_M1003_b N_VPWR_c_158_n 0.0533288f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_158_n 0.356873f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_45 N_VPB_c_23_p N_VPWR_c_158_n 0.017378f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_46 N_VPB_M1003_b Y 0.0687178f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_47 VPB Y 7.75439e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_48 N_VPB_c_23_p Y 0.0133691f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_49 A2 A1 0.0143444f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_50 N_A2_c_51_n A1 0.00100828f $X=1.105 $Y=1.75 $X2=0 $Y2=0
cc_51 N_A2_M1003_g N_A1_M1004_g 0.0235148f $X=0.815 $Y=2.965 $X2=0 $Y2=0
cc_52 N_A2_M1000_g N_A1_M1004_g 0.11556f $X=1.105 $Y=0.91 $X2=0 $Y2=0
cc_53 A2 N_A1_M1004_g 2.84513e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_54 N_A2_M1003_g N_A_56_443#_c_126_n 0.00856321f $X=0.815 $Y=2.965 $X2=0 $Y2=0
cc_55 N_A2_M1003_g N_A_56_443#_c_129_n 0.0119376f $X=0.815 $Y=2.965 $X2=0 $Y2=0
cc_56 A2 N_A_56_443#_c_129_n 0.0540158f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_57 N_A2_c_51_n N_A_56_443#_c_129_n 0.0317378f $X=1.105 $Y=1.75 $X2=0 $Y2=0
cc_58 A2 N_A_56_443#_c_130_n 0.0207942f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_59 N_A2_M1003_g N_VPWR_c_155_n 0.0724558f $X=0.815 $Y=2.965 $X2=0 $Y2=0
cc_60 N_A2_c_51_n N_VPWR_c_155_n 0.00199241f $X=1.105 $Y=1.75 $X2=0 $Y2=0
cc_61 N_A2_M1003_g N_VPWR_c_158_n 0.00882348f $X=0.815 $Y=2.965 $X2=0 $Y2=0
cc_62 N_A2_M1000_g N_VGND_c_206_n 0.0733244f $X=1.105 $Y=0.91 $X2=3.12 $Y2=0
cc_63 A2 N_VGND_c_206_n 0.0765049f $X=1.115 $Y=1.58 $X2=3.12 $Y2=0
cc_64 N_A2_c_51_n N_VGND_c_206_n 0.00874501f $X=1.105 $Y=1.75 $X2=3.12 $Y2=0
cc_65 A1 N_B1_c_98_n 7.76131e-19 $X=1.595 $Y=1.58 $X2=3.12 $Y2=0
cc_66 N_A1_M1004_g N_B1_c_98_n 0.0502776f $X=1.815 $Y=0.91 $X2=3.12 $Y2=0
cc_67 N_A1_M1004_g N_B1_c_107_n 0.00117094f $X=1.815 $Y=0.91 $X2=3.12 $Y2=0
cc_68 N_A1_M1004_g N_B1_c_99_n 0.0202414f $X=1.815 $Y=0.91 $X2=0 $Y2=0
cc_69 A1 N_A_56_443#_c_129_n 0.0233149f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_70 N_A1_M1004_g N_A_56_443#_c_129_n 0.0313866f $X=1.815 $Y=0.91 $X2=0 $Y2=0
cc_71 N_A1_M1004_g N_A_56_443#_c_131_n 0.00390345f $X=1.815 $Y=0.91 $X2=3.12
+ $Y2=0
cc_72 N_A1_M1004_g N_VPWR_c_155_n 0.0966717f $X=1.815 $Y=0.91 $X2=0 $Y2=0
cc_73 N_A1_M1004_g N_VPWR_c_158_n 0.00803924f $X=1.815 $Y=0.91 $X2=0 $Y2=0
cc_74 N_A1_M1004_g N_Y_c_177_n 0.00994158f $X=1.815 $Y=0.91 $X2=0 $Y2=0
cc_75 A1 N_Y_c_180_n 0.00653648f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_76 N_A1_M1004_g N_Y_c_180_n 0.00265785f $X=1.815 $Y=0.91 $X2=0 $Y2=0
cc_77 A1 N_VGND_c_206_n 0.0260011f $X=1.595 $Y=1.58 $X2=3.12 $Y2=0
cc_78 N_A1_M1004_g N_VGND_c_206_n 0.0702762f $X=1.815 $Y=0.91 $X2=3.12 $Y2=0
cc_79 N_A1_M1004_g N_VGND_c_208_n 4.39341e-19 $X=1.815 $Y=0.91 $X2=0 $Y2=0
cc_80 N_A1_M1004_g N_VGND_c_210_n 0.00317792f $X=1.815 $Y=0.91 $X2=1.68 $Y2=0
cc_81 N_B1_c_98_n N_A_56_443#_c_129_n 0.0016752f $X=2.635 $Y=1.89 $X2=0 $Y2=0
cc_82 N_B1_c_107_n N_A_56_443#_c_129_n 0.0137302f $X=2.635 $Y=1.89 $X2=0 $Y2=0
cc_83 N_B1_c_98_n N_A_56_443#_c_131_n 0.00449023f $X=2.635 $Y=1.89 $X2=3.12
+ $Y2=0
cc_84 N_B1_c_107_n N_A_56_443#_c_131_n 0.0456233f $X=2.635 $Y=1.89 $X2=3.12
+ $Y2=0
cc_85 N_B1_c_107_n N_VPWR_c_158_n 0.0158931f $X=2.635 $Y=1.89 $X2=0 $Y2=0
cc_86 N_B1_c_102_n N_VPWR_c_158_n 0.0255147f $X=2.645 $Y=2.105 $X2=0 $Y2=0
cc_87 N_B1_c_98_n N_Y_c_177_n 0.00616299f $X=2.635 $Y=1.89 $X2=0 $Y2=0
cc_88 N_B1_c_99_n N_Y_c_177_n 0.0213616f $X=2.645 $Y=1.395 $X2=0 $Y2=0
cc_89 N_B1_c_98_n N_Y_c_179_n 0.0345087f $X=2.635 $Y=1.89 $X2=0.24 $Y2=0
cc_90 N_B1_c_107_n N_Y_c_179_n 0.0238596f $X=2.635 $Y=1.89 $X2=0.24 $Y2=0
cc_91 N_B1_c_98_n N_Y_c_180_n 0.00959201f $X=2.635 $Y=1.89 $X2=0 $Y2=0
cc_92 N_B1_c_98_n Y 0.0178508f $X=2.635 $Y=1.89 $X2=0 $Y2=0
cc_93 N_B1_c_107_n Y 0.106516f $X=2.635 $Y=1.89 $X2=0 $Y2=0
cc_94 N_B1_c_102_n Y 0.0476066f $X=2.645 $Y=2.105 $X2=0 $Y2=0
cc_95 N_B1_c_99_n N_VGND_c_206_n 8.13181e-19 $X=2.645 $Y=1.395 $X2=3.12 $Y2=0
cc_96 N_B1_c_99_n N_VGND_c_208_n 0.0458846f $X=2.645 $Y=1.395 $X2=0 $Y2=0
cc_97 N_B1_c_99_n N_VGND_c_210_n 0.0125521f $X=2.645 $Y=1.395 $X2=1.68 $Y2=0
cc_98 N_A_56_443#_c_126_n N_VPWR_c_155_n 0.0620876f $X=0.425 $Y=2.34 $X2=0 $Y2=0
cc_99 N_A_56_443#_c_129_n N_VPWR_c_155_n 0.0891231f $X=2.12 $Y=2.015 $X2=0 $Y2=0
cc_100 N_A_56_443#_c_131_n N_VPWR_c_155_n 0.0620165f $X=2.205 $Y=2.34 $X2=0
+ $Y2=0
cc_101 N_A_56_443#_M1003_s N_VPWR_c_158_n 0.00221032f $X=0.28 $Y=2.215 $X2=3.12
+ $Y2=4.07
cc_102 N_A_56_443#_M1005_d N_VPWR_c_158_n 0.00442064f $X=2.065 $Y=2.215 $X2=3.12
+ $Y2=4.07
cc_103 N_A_56_443#_c_126_n N_VPWR_c_158_n 0.0367512f $X=0.425 $Y=2.34 $X2=3.12
+ $Y2=4.07
cc_104 N_A_56_443#_c_131_n N_VPWR_c_158_n 0.0302124f $X=2.205 $Y=2.34 $X2=3.12
+ $Y2=4.07
cc_105 N_A_56_443#_c_129_n N_Y_c_180_n 0.00435725f $X=2.12 $Y=2.015 $X2=0.24
+ $Y2=4.07
cc_106 N_A_56_443#_c_129_n N_VGND_c_206_n 0.0116804f $X=2.12 $Y=2.015 $X2=3.12
+ $Y2=4.07
cc_107 N_VPWR_c_158_n N_Y_M1001_d 0.00567177f $X=1.855 $Y=3.59 $X2=0 $Y2=0
cc_108 N_VPWR_c_158_n Y 0.042328f $X=1.855 $Y=3.59 $X2=0 $Y2=0
cc_109 N_Y_c_177_n N_VGND_c_206_n 0.0623992f $X=2.305 $Y=0.66 $X2=3.12 $Y2=0
cc_110 N_Y_c_177_n N_VGND_c_208_n 0.0499691f $X=2.305 $Y=0.66 $X2=0 $Y2=0
cc_111 N_Y_c_179_n N_VGND_c_208_n 0.0207619f $X=2.98 $Y=1.54 $X2=0 $Y2=0
cc_112 N_Y_c_181_n N_VGND_c_208_n 0.0215754f $X=3.107 $Y=1.625 $X2=0 $Y2=0
cc_113 N_Y_M1004_d N_VGND_c_210_n 0.00650585f $X=2.065 $Y=0.535 $X2=1.68 $Y2=0
cc_114 N_Y_c_177_n N_VGND_c_210_n 0.0244142f $X=2.305 $Y=0.66 $X2=1.68 $Y2=0
