* File: sky130_fd_sc_hvl__and3_1.pxi.spice
* Created: Fri Aug 28 09:32:43 2020
* 
x_PM_SKY130_FD_SC_HVL__AND3_1%VNB N_VNB_M1002_b VNB N_VNB_c_8_p VNB
+ PM_SKY130_FD_SC_HVL__AND3_1%VNB
x_PM_SKY130_FD_SC_HVL__AND3_1%VPB N_VPB_M1007_b VPB N_VPB_c_29_p VPB
+ PM_SKY130_FD_SC_HVL__AND3_1%VPB
x_PM_SKY130_FD_SC_HVL__AND3_1%A N_A_M1007_g N_A_M1002_g A A N_A_c_50_n
+ N_A_c_51_n PM_SKY130_FD_SC_HVL__AND3_1%A
x_PM_SKY130_FD_SC_HVL__AND3_1%B B B N_B_M1003_g N_B_c_74_n N_B_M1000_g
+ PM_SKY130_FD_SC_HVL__AND3_1%B
x_PM_SKY130_FD_SC_HVL__AND3_1%C N_C_M1004_g N_C_M1006_g C C C N_C_c_95_n
+ N_C_c_96_n PM_SKY130_FD_SC_HVL__AND3_1%C
x_PM_SKY130_FD_SC_HVL__AND3_1%A_30_517# N_A_30_517#_M1002_s N_A_30_517#_M1007_s
+ N_A_30_517#_M1000_d N_A_30_517#_M1005_g N_A_30_517#_M1001_g
+ N_A_30_517#_c_131_n N_A_30_517#_c_140_n N_A_30_517#_c_132_n
+ N_A_30_517#_c_142_n N_A_30_517#_c_133_n N_A_30_517#_c_134_n
+ N_A_30_517#_c_135_n N_A_30_517#_c_170_n N_A_30_517#_c_136_n
+ PM_SKY130_FD_SC_HVL__AND3_1%A_30_517#
x_PM_SKY130_FD_SC_HVL__AND3_1%VPWR N_VPWR_M1007_d N_VPWR_M1006_d VPWR
+ N_VPWR_c_196_n N_VPWR_c_199_n N_VPWR_c_202_n PM_SKY130_FD_SC_HVL__AND3_1%VPWR
x_PM_SKY130_FD_SC_HVL__AND3_1%X N_X_M1001_d N_X_M1005_d X X X X X X X
+ N_X_c_226_n X PM_SKY130_FD_SC_HVL__AND3_1%X
x_PM_SKY130_FD_SC_HVL__AND3_1%VGND N_VGND_M1004_d VGND N_VGND_c_245_n
+ N_VGND_c_247_n PM_SKY130_FD_SC_HVL__AND3_1%VGND
cc_1 N_VNB_M1002_b N_A_c_50_n 0.0534941f $X=-0.33 $Y=-0.265 $X2=0.77 $Y2=1.56
cc_2 N_VNB_M1002_b N_A_c_51_n 0.0535845f $X=-0.33 $Y=-0.265 $X2=0.72 $Y2=1.395
cc_3 N_VNB_M1002_b N_B_M1003_g 0.0854757f $X=-0.33 $Y=-0.265 $X2=0.755 $Y2=1.075
cc_4 N_VNB_M1002_b C 0.00959842f $X=-0.33 $Y=-0.265 $X2=0.72 $Y2=1.56
cc_5 N_VNB_M1002_b N_C_c_95_n 0.0493889f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_M1002_b N_C_c_96_n 0.0504574f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_7 N_VNB_M1002_b N_A_30_517#_M1001_g 0.0493995f $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=1.895
cc_8 N_VNB_c_8_p N_A_30_517#_M1001_g 8.65757e-19 $X=0.24 $Y=0 $X2=0.72 $Y2=1.895
cc_9 N_VNB_M1002_b N_A_30_517#_c_131_n 0.0509202f $X=-0.33 $Y=-0.265 $X2=0.77
+ $Y2=1.295
cc_10 N_VNB_M1002_b N_A_30_517#_c_132_n 0.00553035f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1002_b N_A_30_517#_c_133_n 0.0057957f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1002_b N_A_30_517#_c_134_n 0.00272105f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1002_b N_A_30_517#_c_135_n 0.00148421f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_M1002_b N_A_30_517#_c_136_n 0.0519301f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_15 N_VNB_M1002_b N_X_c_226_n 0.0619021f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_16 N_VNB_c_8_p N_X_c_226_n 7.40038e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_17 N_VNB_M1002_b N_VGND_c_245_n 0.0602519f $X=-0.33 $Y=-0.265 $X2=0.755
+ $Y2=1.075
cc_18 N_VNB_c_8_p N_VGND_c_245_n 0.00227897f $X=0.24 $Y=0 $X2=0.755 $Y2=1.075
cc_19 N_VNB_M1002_b N_VGND_c_247_n 0.129686f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=0.84
cc_20 N_VNB_c_8_p N_VGND_c_247_n 0.410937f $X=0.24 $Y=0 $X2=0.635 $Y2=0.84
cc_21 N_VPB_M1007_b N_A_M1007_g 0.094578f $X=-0.33 $Y=1.885 $X2=0.685 $Y2=2.795
cc_22 N_VPB_M1007_b N_A_c_50_n 0.00298978f $X=-0.33 $Y=1.885 $X2=0.77 $Y2=1.56
cc_23 N_VPB_M1007_b N_B_M1003_g 0.0889222f $X=-0.33 $Y=1.885 $X2=0.755 $Y2=1.075
cc_24 N_VPB_M1007_b N_B_c_74_n 0.00509122f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_25 N_VPB_M1007_b N_C_M1006_g 0.0868724f $X=-0.33 $Y=1.885 $X2=0.755 $Y2=1.075
cc_26 N_VPB_M1007_b N_C_c_95_n 0.00287806f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_27 N_VPB_M1007_b N_A_30_517#_M1005_g 0.0421265f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=1.56
cc_28 VPB N_A_30_517#_M1005_g 0.00970178f $X=0 $Y=3.955 $X2=0.72 $Y2=1.56
cc_29 N_VPB_c_29_p N_A_30_517#_M1005_g 0.0162989f $X=3.6 $Y=4.07 $X2=0.72
+ $Y2=1.56
cc_30 N_VPB_M1007_b N_A_30_517#_c_140_n 0.0520466f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_31 N_VPB_M1007_b N_A_30_517#_c_132_n 0.00478659f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_32 N_VPB_M1007_b N_A_30_517#_c_142_n 0.00931153f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_33 N_VPB_M1007_b N_A_30_517#_c_133_n 0.0038334f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_34 N_VPB_M1007_b N_A_30_517#_c_134_n 0.00682132f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_35 N_VPB_M1007_b N_A_30_517#_c_136_n 0.0220634f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_36 N_VPB_M1007_b N_VPWR_c_196_n 0.0506373f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_196_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_38 N_VPB_c_29_p N_VPWR_c_196_n 0.0409968f $X=3.6 $Y=4.07 $X2=0 $Y2=0
cc_39 N_VPB_M1007_b N_VPWR_c_199_n 0.03028f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_199_n 0.00335473f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_41 N_VPB_c_29_p N_VPWR_c_199_n 0.0490696f $X=3.6 $Y=4.07 $X2=0 $Y2=0
cc_42 N_VPB_M1007_b N_VPWR_c_202_n 0.0787033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_202_n 0.40979f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_44 N_VPB_c_29_p N_VPWR_c_202_n 0.0202928f $X=3.6 $Y=4.07 $X2=0 $Y2=0
cc_45 N_VPB_M1007_b X 0.0071429f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_46 N_VPB_M1007_b N_X_c_226_n 0.0126954f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_47 N_VPB_M1007_b X 0.0486863f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_48 VPB X 0.00110823f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_49 N_VPB_c_29_p X 0.0182942f $X=3.6 $Y=4.07 $X2=0 $Y2=0
cc_50 N_A_M1007_g N_B_M1003_g 0.0437572f $X=0.685 $Y=2.795 $X2=0 $Y2=0
cc_51 A N_B_M1003_g 7.63528e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_52 N_A_c_51_n N_B_M1003_g 0.0785565f $X=0.72 $Y=1.395 $X2=0 $Y2=0
cc_53 N_A_M1007_g N_B_c_74_n 0.0263931f $X=0.685 $Y=2.795 $X2=0.24 $Y2=0
cc_54 N_A_c_50_n N_B_c_74_n 3.95025e-19 $X=0.77 $Y=1.56 $X2=0.24 $Y2=0
cc_55 A C 0.0665032f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_56 N_A_c_51_n C 0.00623468f $X=0.72 $Y=1.395 $X2=0 $Y2=0
cc_57 A N_A_30_517#_c_131_n 0.0609427f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_58 N_A_c_50_n N_A_30_517#_c_131_n 0.016851f $X=0.77 $Y=1.56 $X2=0 $Y2=0
cc_59 N_A_c_51_n N_A_30_517#_c_131_n 0.00618774f $X=0.72 $Y=1.395 $X2=0 $Y2=0
cc_60 N_A_M1007_g N_A_30_517#_c_140_n 0.023891f $X=0.685 $Y=2.795 $X2=1.92
+ $Y2=0.058
cc_61 N_A_M1007_g N_A_30_517#_c_132_n 0.0192586f $X=0.685 $Y=2.795 $X2=0 $Y2=0
cc_62 A N_A_30_517#_c_132_n 0.0238596f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_63 N_A_c_50_n N_A_30_517#_c_132_n 0.0219675f $X=0.77 $Y=1.56 $X2=0 $Y2=0
cc_64 N_A_M1007_g N_VPWR_c_196_n 0.0400939f $X=0.685 $Y=2.795 $X2=0.24 $Y2=0
cc_65 N_A_M1007_g N_VPWR_c_202_n 0.0036578f $X=0.685 $Y=2.795 $X2=0 $Y2=0
cc_66 A N_VGND_c_247_n 0.0171859f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_67 N_A_c_51_n N_VGND_c_247_n 0.016332f $X=0.72 $Y=1.395 $X2=0 $Y2=0
cc_68 N_B_M1003_g N_C_M1006_g 0.0379545f $X=1.465 $Y=1.075 $X2=0 $Y2=0
cc_69 N_B_c_74_n N_C_M1006_g 2.25959e-19 $X=1.4 $Y=2.26 $X2=0 $Y2=0
cc_70 N_B_M1003_g C 0.065831f $X=1.465 $Y=1.075 $X2=0 $Y2=0
cc_71 N_B_M1003_g N_C_c_96_n 0.0793101f $X=1.465 $Y=1.075 $X2=1.92 $Y2=0.057
cc_72 N_B_c_74_n N_A_30_517#_c_140_n 0.0208158f $X=1.4 $Y=2.26 $X2=1.92
+ $Y2=0.058
cc_73 N_B_M1003_g N_A_30_517#_c_132_n 0.0301404f $X=1.465 $Y=1.075 $X2=0 $Y2=0
cc_74 N_B_c_74_n N_A_30_517#_c_132_n 0.0674562f $X=1.4 $Y=2.26 $X2=0 $Y2=0
cc_75 N_B_M1003_g N_A_30_517#_c_142_n 0.0108589f $X=1.465 $Y=1.075 $X2=0 $Y2=0
cc_76 N_B_c_74_n N_A_30_517#_c_142_n 0.0223247f $X=1.4 $Y=2.26 $X2=0 $Y2=0
cc_77 N_B_M1003_g N_VPWR_c_196_n 0.0317375f $X=1.465 $Y=1.075 $X2=0.24 $Y2=0
cc_78 N_B_c_74_n N_VPWR_c_196_n 0.0656273f $X=1.4 $Y=2.26 $X2=0.24 $Y2=0
cc_79 N_B_M1003_g N_VPWR_c_199_n 6.36294e-19 $X=1.465 $Y=1.075 $X2=0 $Y2=0
cc_80 N_B_M1003_g N_VPWR_c_202_n 0.00598021f $X=1.465 $Y=1.075 $X2=0 $Y2=0
cc_81 N_B_M1003_g N_VGND_c_247_n 0.016332f $X=1.465 $Y=1.075 $X2=0 $Y2=0
cc_82 N_C_M1006_g N_A_30_517#_M1005_g 0.0220815f $X=2.245 $Y=2.795 $X2=0 $Y2=0
cc_83 C N_A_30_517#_M1001_g 5.5788e-19 $X=2.075 $Y=0.84 $X2=3.6 $Y2=0
cc_84 N_C_c_95_n N_A_30_517#_M1001_g 7.16196e-19 $X=2.09 $Y=1.56 $X2=3.6 $Y2=0
cc_85 N_C_c_96_n N_A_30_517#_M1001_g 0.00862659f $X=2.21 $Y=1.395 $X2=3.6 $Y2=0
cc_86 C N_A_30_517#_c_132_n 0.0486953f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_87 N_C_M1006_g N_A_30_517#_c_142_n 0.0290252f $X=2.245 $Y=2.795 $X2=0 $Y2=0
cc_88 N_C_M1006_g N_A_30_517#_c_133_n 0.0179837f $X=2.245 $Y=2.795 $X2=0 $Y2=0
cc_89 C N_A_30_517#_c_133_n 0.016986f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_90 N_C_c_95_n N_A_30_517#_c_133_n 0.0167117f $X=2.09 $Y=1.56 $X2=0 $Y2=0
cc_91 N_C_M1006_g N_A_30_517#_c_135_n 0.00141015f $X=2.245 $Y=2.795 $X2=0 $Y2=0
cc_92 C N_A_30_517#_c_135_n 0.0215307f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_93 N_C_c_95_n N_A_30_517#_c_135_n 0.00444457f $X=2.09 $Y=1.56 $X2=0 $Y2=0
cc_94 N_C_c_95_n N_A_30_517#_c_170_n 0.00115778f $X=2.09 $Y=1.56 $X2=0 $Y2=0
cc_95 C N_A_30_517#_c_136_n 0.00102611f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_96 N_C_c_95_n N_A_30_517#_c_136_n 0.0220815f $X=2.09 $Y=1.56 $X2=0 $Y2=0
cc_97 N_C_M1006_g N_VPWR_c_196_n 5.74502e-19 $X=2.245 $Y=2.795 $X2=0.24 $Y2=0
cc_98 N_C_M1006_g N_VPWR_c_199_n 0.0667798f $X=2.245 $Y=2.795 $X2=0 $Y2=0
cc_99 N_C_M1006_g N_VPWR_c_202_n 0.00598021f $X=2.245 $Y=2.795 $X2=0 $Y2=0
cc_100 C A_201_173# 0.00367414f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_101 C N_VGND_c_245_n 0.0247942f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_102 N_C_c_95_n N_VGND_c_245_n 0.00215536f $X=2.09 $Y=1.56 $X2=0 $Y2=0
cc_103 N_C_c_96_n N_VGND_c_245_n 0.00842317f $X=2.21 $Y=1.395 $X2=0 $Y2=0
cc_104 C N_VGND_c_247_n 0.0609311f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_105 N_C_c_96_n N_VGND_c_247_n 0.016332f $X=2.21 $Y=1.395 $X2=0 $Y2=0
cc_106 N_A_30_517#_c_140_n N_VPWR_c_196_n 0.0165118f $X=0.295 $Y=2.795 $X2=0.24
+ $Y2=0
cc_107 N_A_30_517#_c_132_n N_VPWR_c_196_n 0.001054f $X=1.77 $Y=1.91 $X2=0.24
+ $Y2=0
cc_108 N_A_30_517#_c_142_n N_VPWR_c_196_n 0.0123528f $X=1.855 $Y=2.795 $X2=0.24
+ $Y2=0
cc_109 N_A_30_517#_M1005_g N_VPWR_c_199_n 0.0702304f $X=3.14 $Y=2.965 $X2=0
+ $Y2=0
cc_110 N_A_30_517#_c_142_n N_VPWR_c_199_n 0.0647238f $X=1.855 $Y=2.795 $X2=0
+ $Y2=0
cc_111 N_A_30_517#_c_133_n N_VPWR_c_199_n 0.0548777f $X=2.91 $Y=1.91 $X2=0 $Y2=0
cc_112 N_A_30_517#_c_170_n N_VPWR_c_199_n 0.0182317f $X=3.075 $Y=1.83 $X2=0
+ $Y2=0
cc_113 N_A_30_517#_M1005_g N_VPWR_c_202_n 0.0130385f $X=3.14 $Y=2.965 $X2=0
+ $Y2=0
cc_114 N_A_30_517#_c_140_n N_VPWR_c_202_n 0.0113682f $X=0.295 $Y=2.795 $X2=0
+ $Y2=0
cc_115 N_A_30_517#_c_142_n N_VPWR_c_202_n 0.0112714f $X=1.855 $Y=2.795 $X2=0
+ $Y2=0
cc_116 N_A_30_517#_M1005_g X 0.00522528f $X=3.14 $Y=2.965 $X2=0.24 $Y2=0
cc_117 N_A_30_517#_c_136_n X 0.0010557f $X=3.075 $Y=1.83 $X2=0.24 $Y2=0
cc_118 N_A_30_517#_M1005_g N_X_c_226_n 0.00441217f $X=3.14 $Y=2.965 $X2=1.92
+ $Y2=0.058
cc_119 N_A_30_517#_M1001_g N_X_c_226_n 0.0207531f $X=3.175 $Y=0.91 $X2=1.92
+ $Y2=0.058
cc_120 N_A_30_517#_c_170_n N_X_c_226_n 0.0246163f $X=3.075 $Y=1.83 $X2=1.92
+ $Y2=0.058
cc_121 N_A_30_517#_c_136_n N_X_c_226_n 0.0344353f $X=3.075 $Y=1.83 $X2=1.92
+ $Y2=0.058
cc_122 N_A_30_517#_M1005_g X 0.0260387f $X=3.14 $Y=2.965 $X2=0 $Y2=0
cc_123 N_A_30_517#_M1001_g N_VGND_c_245_n 0.0568157f $X=3.175 $Y=0.91 $X2=0
+ $Y2=0
cc_124 N_A_30_517#_c_133_n N_VGND_c_245_n 0.0186107f $X=2.91 $Y=1.91 $X2=0 $Y2=0
cc_125 N_A_30_517#_c_170_n N_VGND_c_245_n 0.0150943f $X=3.075 $Y=1.83 $X2=0
+ $Y2=0
cc_126 N_A_30_517#_c_136_n N_VGND_c_245_n 0.001227f $X=3.075 $Y=1.83 $X2=0 $Y2=0
cc_127 N_A_30_517#_M1001_g N_VGND_c_247_n 0.0109073f $X=3.175 $Y=0.91 $X2=0
+ $Y2=0
cc_128 N_A_30_517#_c_131_n N_VGND_c_247_n 0.0163004f $X=0.34 $Y=1.075 $X2=0
+ $Y2=0
cc_129 N_VPWR_c_199_n X 0.0995832f $X=2.75 $Y=2.34 $X2=0 $Y2=0
cc_130 N_VPWR_c_202_n X 0.045435f $X=3.035 $Y=3.59 $X2=0 $Y2=0
cc_131 N_X_c_226_n N_VGND_c_245_n 0.0638037f $X=3.565 $Y=0.68 $X2=0 $Y2=0
cc_132 N_X_c_226_n N_VGND_c_247_n 0.0309744f $X=3.565 $Y=0.68 $X2=0 $Y2=0
