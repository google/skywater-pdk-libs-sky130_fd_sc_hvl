* File: sky130_fd_sc_hvl__buf_32.pex.spice
* Created: Wed Sep  2 09:04:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__BUF_32%VNB 5 7 17 25 27
r154 25 27 0.30797 $w=2.3e-07 $l=4.8e-07 $layer=MET1_cond $X=24.765 $Y=0
+ $X2=25.245 $Y2=0
r155 17 27 5.20662 $w=2.3e-07 $l=8.115e-06 $layer=MET1_cond $X=33.36 $Y=0
+ $X2=25.245 $Y2=0
r156 7 25 5.11038 $w=2.3e-07 $l=7.965e-06 $layer=MET1_cond $X=16.8 $Y=0
+ $X2=24.765 $Y2=0
r157 7 11 10.625 $w=2.3e-07 $l=1.656e-05 $layer=MET1_cond $X=16.8 $Y=0 $X2=0.24
+ $Y2=0
r158 5 17 0.265714 $w=1.7e-07 $l=5.95e-06 $layer=mcon $count=35 $X=33.36 $Y=0
+ $X2=33.36 $Y2=0
r159 5 11 0.265714 $w=1.7e-07 $l=5.95e-06 $layer=mcon $count=35 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_32%VPB 4 6 14 15 22 24
r256 22 24 0.30797 $w=2.3e-07 $l=4.8e-07 $layer=MET1_cond $X=24.765 $Y=4.07
+ $X2=25.245 $Y2=4.07
r257 15 24 5.20662 $w=2.3e-07 $l=8.115e-06 $layer=MET1_cond $X=33.36 $Y=4.07
+ $X2=25.245 $Y2=4.07
r258 14 15 0.265714 $w=1.7e-07 $l=5.95e-06 $layer=mcon $count=35 $X=33.36
+ $Y=4.07 $X2=33.36 $Y2=4.07
r259 9 14 2160.77 $w=1.68e-07 $l=3.312e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=33.36 $Y2=4.07
r260 9 10 0.265714 $w=1.7e-07 $l=5.95e-06 $layer=mcon $count=35 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r261 6 22 5.11038 $w=2.3e-07 $l=7.965e-06 $layer=MET1_cond $X=16.8 $Y=4.07
+ $X2=24.765 $Y2=4.07
r262 6 10 10.625 $w=2.3e-07 $l=1.656e-05 $layer=MET1_cond $X=16.8 $Y=4.07
+ $X2=0.24 $Y2=4.07
r263 4 14 5.2 $w=1.7e-07 $l=3.34025e-05 $layer=licon1_NTAP_notbjt $count=35 $X=0
+ $Y=3.985 $X2=33.36 $Y2=4.07
r264 4 9 5.2 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=35 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_32%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34
+ 36 38 41 43 45 48 50 52 55 57 59 62 64 66 69 71 72 73 74 75 76 77 96 101
c203 13 0 3.19988e-20 $X=1.445 $Y=2.965
r204 100 101 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=6.905 $Y=1.815
+ $X2=7.685 $Y2=1.815
r205 99 100 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=6.125 $Y=1.815
+ $X2=6.905 $Y2=1.815
r206 98 99 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=5.345 $Y=1.815
+ $X2=6.125 $Y2=1.815
r207 97 98 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=4.565 $Y=1.815
+ $X2=5.345 $Y2=1.815
r208 95 97 10.7006 $w=5e-07 $l=1e-07 $layer=POLY_cond $X=4.465 $Y=1.815
+ $X2=4.565 $Y2=1.815
r209 95 96 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6 $X=4.465
+ $Y=1.73 $X2=4.465 $Y2=1.73
r210 93 95 72.764 $w=5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.785 $Y=1.815
+ $X2=4.465 $Y2=1.815
r211 92 93 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.005 $Y=1.815
+ $X2=3.785 $Y2=1.815
r212 91 92 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.225 $Y=1.815
+ $X2=3.005 $Y2=1.815
r213 90 91 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.445 $Y=1.815
+ $X2=2.225 $Y2=1.815
r214 89 90 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.665 $Y=1.815
+ $X2=1.445 $Y2=1.815
r215 86 89 29.9617 $w=5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.385 $Y=1.815
+ $X2=0.665 $Y2=1.815
r216 86 87 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6 $X=0.385
+ $Y=1.73 $X2=0.385 $Y2=1.73
r217 77 96 42.4197 $w=2.33e-07 $l=8.65e-07 $layer=LI1_cond $X=3.6 $Y=1.697
+ $X2=4.465 $Y2=1.697
r218 76 77 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.697
+ $X2=3.6 $Y2=1.697
r219 75 76 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.697
+ $X2=3.12 $Y2=1.697
r220 74 75 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.697
+ $X2=2.64 $Y2=1.697
r221 73 74 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.697
+ $X2=2.16 $Y2=1.697
r222 72 73 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.697
+ $X2=1.68 $Y2=1.697
r223 71 72 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.697
+ $X2=1.2 $Y2=1.697
r224 71 87 16.4284 $w=2.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.72 $Y=1.697
+ $X2=0.385 $Y2=1.697
r225 67 101 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.685 $Y=2.065
+ $X2=7.685 $Y2=1.815
r226 67 69 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=7.685 $Y=2.065
+ $X2=7.685 $Y2=2.965
r227 64 101 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.685 $Y=1.565
+ $X2=7.685 $Y2=1.815
r228 64 66 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.685 $Y=1.565
+ $X2=7.685 $Y2=1.08
r229 60 100 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.905 $Y=2.065
+ $X2=6.905 $Y2=1.815
r230 60 62 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=6.905 $Y=2.065
+ $X2=6.905 $Y2=2.965
r231 57 100 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.905 $Y=1.565
+ $X2=6.905 $Y2=1.815
r232 57 59 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.905 $Y=1.565
+ $X2=6.905 $Y2=1.08
r233 53 99 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.125 $Y=2.065
+ $X2=6.125 $Y2=1.815
r234 53 55 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=6.125 $Y=2.065
+ $X2=6.125 $Y2=2.965
r235 50 99 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.125 $Y=1.565
+ $X2=6.125 $Y2=1.815
r236 50 52 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.125 $Y=1.565
+ $X2=6.125 $Y2=1.08
r237 46 98 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.345 $Y=2.065
+ $X2=5.345 $Y2=1.815
r238 46 48 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=5.345 $Y=2.065
+ $X2=5.345 $Y2=2.965
r239 43 98 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.345 $Y=1.565
+ $X2=5.345 $Y2=1.815
r240 43 45 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=5.345 $Y=1.565
+ $X2=5.345 $Y2=1.08
r241 39 97 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.565 $Y=2.065
+ $X2=4.565 $Y2=1.815
r242 39 41 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=4.565 $Y=2.065
+ $X2=4.565 $Y2=2.965
r243 36 97 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.565 $Y=1.565
+ $X2=4.565 $Y2=1.815
r244 36 38 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.565 $Y=1.565
+ $X2=4.565 $Y2=1.08
r245 32 93 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.785 $Y=2.065
+ $X2=3.785 $Y2=1.815
r246 32 34 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=3.785 $Y=2.065
+ $X2=3.785 $Y2=2.965
r247 29 93 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.785 $Y=1.565
+ $X2=3.785 $Y2=1.815
r248 29 31 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.785 $Y=1.565
+ $X2=3.785 $Y2=1.08
r249 25 92 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.005 $Y=2.065
+ $X2=3.005 $Y2=1.815
r250 25 27 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=3.005 $Y=2.065
+ $X2=3.005 $Y2=2.965
r251 22 92 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.005 $Y=1.565
+ $X2=3.005 $Y2=1.815
r252 22 24 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.005 $Y=1.565
+ $X2=3.005 $Y2=1.08
r253 18 91 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.225 $Y=2.065
+ $X2=2.225 $Y2=1.815
r254 18 20 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=2.225 $Y=2.065
+ $X2=2.225 $Y2=2.965
r255 15 91 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.225 $Y=1.565
+ $X2=2.225 $Y2=1.815
r256 15 17 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.225 $Y=1.565
+ $X2=2.225 $Y2=1.08
r257 11 90 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.445 $Y=2.065
+ $X2=1.445 $Y2=1.815
r258 11 13 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=1.445 $Y=2.065
+ $X2=1.445 $Y2=2.965
r259 8 90 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.445 $Y=1.565
+ $X2=1.445 $Y2=1.815
r260 8 10 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.445 $Y=1.565
+ $X2=1.445 $Y2=1.08
r261 4 89 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.665 $Y=2.065
+ $X2=0.665 $Y2=1.815
r262 4 6 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=0.665 $Y=2.065 $X2=0.665
+ $Y2=2.965
r263 1 89 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.665 $Y=1.565
+ $X2=0.665 $Y2=1.815
r264 1 3 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.665 $Y=1.565
+ $X2=0.665 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_32%A_183_141# 1 2 3 4 5 6 7 8 9 10 31 33 36 38
+ 40 43 45 47 50 52 54 57 59 61 64 66 68 71 73 75 78 80 82 85 87 89 92 94 96 99
+ 101 103 106 108 110 113 115 117 120 122 124 127 129 131 134 136 138 141 143
+ 145 148 150 152 155 157 159 162 164 166 169 171 173 176 178 180 183 185 187
+ 190 192 194 197 199 201 204 206 208 211 213 215 218 220 222 225 227 229 232
+ 234 236 239 241 243 246 248 250 253 257 261 265 266 267 268 271 275 279 281
+ 285 291 293 295 299 303 307 308 311 317 319 320 321 322 329 332 335 338 341
+ 344 347 350 353 356 359 362 365 368 371 373 374
r796 501 502 0.456075 $w=1.068e-06 $l=4e-08 $layer=LI1_cond $X=5.675 $Y=1.73
+ $X2=5.715 $Y2=1.73
r797 374 450 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=31.865
+ $Y=1.73 $X2=31.865 $Y2=1.73
r798 373 374 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=31.875 $Y=1.665
+ $X2=31.875 $Y2=1.665
r799 371 445 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=30.305
+ $Y=1.73 $X2=30.305 $Y2=1.73
r800 370 373 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=30.315 $Y=1.665
+ $X2=31.875 $Y2=1.665
r801 370 371 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=30.315 $Y=1.665
+ $X2=30.315 $Y2=1.665
r802 368 440 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=28.745
+ $Y=1.73 $X2=28.745 $Y2=1.73
r803 367 370 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=28.755 $Y=1.665
+ $X2=30.315 $Y2=1.665
r804 367 368 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=28.755 $Y=1.665
+ $X2=28.755 $Y2=1.665
r805 365 435 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=27.185
+ $Y=1.73 $X2=27.185 $Y2=1.73
r806 364 367 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=27.195 $Y=1.665
+ $X2=28.755 $Y2=1.665
r807 364 365 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=27.195 $Y=1.665
+ $X2=27.195 $Y2=1.665
r808 362 430 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=25.625
+ $Y=1.73 $X2=25.625 $Y2=1.73
r809 361 364 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=25.635 $Y=1.665
+ $X2=27.195 $Y2=1.665
r810 361 362 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=25.635 $Y=1.665
+ $X2=25.635 $Y2=1.665
r811 359 425 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=24.065
+ $Y=1.73 $X2=24.065 $Y2=1.73
r812 358 361 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=24.075 $Y=1.665
+ $X2=25.635 $Y2=1.665
r813 358 359 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=24.075 $Y=1.665
+ $X2=24.075 $Y2=1.665
r814 356 420 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=22.505
+ $Y=1.73 $X2=22.505 $Y2=1.73
r815 355 358 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=22.515 $Y=1.665
+ $X2=24.075 $Y2=1.665
r816 355 356 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=22.515 $Y=1.665
+ $X2=22.515 $Y2=1.665
r817 353 415 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=20.935
+ $Y=1.73 $X2=20.935 $Y2=1.73
r818 352 355 1.00732 $w=2.3e-07 $l=1.57e-06 $layer=MET1_cond $X=20.945 $Y=1.665
+ $X2=22.515 $Y2=1.665
r819 352 353 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.945 $Y=1.665
+ $X2=20.945 $Y2=1.665
r820 350 410 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=19.385
+ $Y=1.73 $X2=19.385 $Y2=1.73
r821 349 352 0.994487 $w=2.3e-07 $l=1.55e-06 $layer=MET1_cond $X=19.395 $Y=1.665
+ $X2=20.945 $Y2=1.665
r822 349 350 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=19.395 $Y=1.665
+ $X2=19.395 $Y2=1.665
r823 347 405 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=17.825
+ $Y=1.73 $X2=17.825 $Y2=1.73
r824 346 349 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=17.835 $Y=1.665
+ $X2=19.395 $Y2=1.665
r825 346 347 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.835 $Y=1.665
+ $X2=17.835 $Y2=1.665
r826 344 400 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=16.265
+ $Y=1.73 $X2=16.265 $Y2=1.73
r827 343 346 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=16.275 $Y=1.665
+ $X2=17.835 $Y2=1.665
r828 343 344 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.275 $Y=1.665
+ $X2=16.275 $Y2=1.665
r829 341 395 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.705
+ $Y=1.73 $X2=14.705 $Y2=1.73
r830 340 343 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=14.715 $Y=1.665
+ $X2=16.275 $Y2=1.665
r831 340 341 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.715 $Y=1.665
+ $X2=14.715 $Y2=1.665
r832 338 390 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.145
+ $Y=1.73 $X2=13.145 $Y2=1.73
r833 337 340 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=13.155 $Y=1.665
+ $X2=14.715 $Y2=1.665
r834 337 338 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.155 $Y=1.665
+ $X2=13.155 $Y2=1.665
r835 335 385 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.585
+ $Y=1.73 $X2=11.585 $Y2=1.73
r836 334 337 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=11.595 $Y=1.665
+ $X2=13.155 $Y2=1.665
r837 334 335 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.595 $Y=1.665
+ $X2=11.595 $Y2=1.665
r838 332 380 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.025
+ $Y=1.73 $X2=10.025 $Y2=1.73
r839 331 334 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=10.035 $Y=1.665
+ $X2=11.595 $Y2=1.665
r840 331 332 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.035 $Y=1.665
+ $X2=10.035 $Y2=1.665
r841 328 331 1.77724 $w=2.3e-07 $l=2.77e-06 $layer=MET1_cond $X=7.265 $Y=1.665
+ $X2=10.035 $Y2=1.665
r842 328 329 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.265
+ $Y=1.665 $X2=7.265 $Y2=1.665
r843 325 501 6.49907 $w=1.068e-06 $l=5.7e-07 $layer=LI1_cond $X=5.105 $Y=1.73
+ $X2=5.675 $Y2=1.73
r844 324 328 1.38587 $w=2.3e-07 $l=2.16e-06 $layer=MET1_cond $X=5.105 $Y=1.665
+ $X2=7.265 $Y2=1.665
r845 324 325 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.105
+ $Y=1.665 $X2=5.105 $Y2=1.665
r846 315 329 12.6925 $w=2.97e-07 $l=5.50768e-07 $layer=LI1_cond $X=7.267
+ $Y=1.195 $X2=7.235 $Y2=1.73
r847 315 317 14.1115 $w=2.43e-07 $l=3e-07 $layer=LI1_cond $X=7.267 $Y=1.195
+ $X2=7.267 $Y2=0.895
r848 311 313 41.1587 $w=3.48e-07 $l=1.25e-06 $layer=LI1_cond $X=7.235 $Y=2.34
+ $X2=7.235 $Y2=3.59
r849 309 329 12.6925 $w=2.97e-07 $l=5.35e-07 $layer=LI1_cond $X=7.235 $Y=2.265
+ $X2=7.235 $Y2=1.73
r850 309 311 2.46952 $w=3.48e-07 $l=7.5e-08 $layer=LI1_cond $X=7.235 $Y=2.265
+ $X2=7.235 $Y2=2.34
r851 308 502 2.22336 $w=1.068e-06 $l=1.95e-07 $layer=LI1_cond $X=5.91 $Y=1.73
+ $X2=5.715 $Y2=1.73
r852 307 329 2.56421 $w=1.07e-06 $l=1.75e-07 $layer=LI1_cond $X=7.06 $Y=1.73
+ $X2=7.235 $Y2=1.73
r853 307 308 13.1121 $w=1.068e-06 $l=1.15e-06 $layer=LI1_cond $X=7.06 $Y=1.73
+ $X2=5.91 $Y2=1.73
r854 303 305 46.4695 $w=3.08e-07 $l=1.25e-06 $layer=LI1_cond $X=5.675 $Y=2.34
+ $X2=5.675 $Y2=3.59
r855 301 501 8.1733 $w=3.1e-07 $l=5.35e-07 $layer=LI1_cond $X=5.675 $Y=2.265
+ $X2=5.675 $Y2=1.73
r856 301 303 2.78817 $w=3.08e-07 $l=7.5e-08 $layer=LI1_cond $X=5.675 $Y=2.265
+ $X2=5.675 $Y2=2.34
r857 297 502 6.72231 $w=3.9e-07 $l=5.35e-07 $layer=LI1_cond $X=5.715 $Y=1.195
+ $X2=5.715 $Y2=1.73
r858 297 299 8.86495 $w=3.88e-07 $l=3e-07 $layer=LI1_cond $X=5.715 $Y=1.195
+ $X2=5.715 $Y2=0.895
r859 296 321 6.19399 $w=2.8e-07 $l=1.75e-07 $layer=LI1_cond $X=4.29 $Y=2.125
+ $X2=4.115 $Y2=2.125
r860 295 325 7.57904 $w=5.35e-07 $l=5.25833e-07 $layer=LI1_cond $X=4.8 $Y=2.125
+ $X2=5.105 $Y2=1.73
r861 295 296 20.9909 $w=2.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.8 $Y=2.125
+ $X2=4.29 $Y2=2.125
r862 294 322 5.75112 $w=2.15e-07 $l=1.23e-07 $layer=LI1_cond $X=4.27 $Y=1.302
+ $X2=4.147 $Y2=1.302
r863 293 325 8.02838 $w=5.35e-07 $l=5.60111e-07 $layer=LI1_cond $X=4.8 $Y=1.302
+ $X2=5.105 $Y2=1.73
r864 293 294 28.4091 $w=2.13e-07 $l=5.3e-07 $layer=LI1_cond $X=4.8 $Y=1.302
+ $X2=4.27 $Y2=1.302
r865 289 322 0.876697 $w=2.45e-07 $l=1.07e-07 $layer=LI1_cond $X=4.147 $Y=1.195
+ $X2=4.147 $Y2=1.302
r866 289 291 14.1115 $w=2.43e-07 $l=3e-07 $layer=LI1_cond $X=4.147 $Y=1.195
+ $X2=4.147 $Y2=0.895
r867 285 287 41.1587 $w=3.48e-07 $l=1.25e-06 $layer=LI1_cond $X=4.115 $Y=2.34
+ $X2=4.115 $Y2=3.59
r868 283 321 0.552779 $w=3.5e-07 $l=1.4e-07 $layer=LI1_cond $X=4.115 $Y=2.265
+ $X2=4.115 $Y2=2.125
r869 283 285 2.46952 $w=3.48e-07 $l=7.5e-08 $layer=LI1_cond $X=4.115 $Y=2.265
+ $X2=4.115 $Y2=2.34
r870 282 319 8.20698 $w=2.15e-07 $l=1.95e-07 $layer=LI1_cond $X=2.79 $Y=1.302
+ $X2=2.595 $Y2=1.302
r871 281 322 5.75112 $w=2.15e-07 $l=1.22e-07 $layer=LI1_cond $X=4.025 $Y=1.302
+ $X2=4.147 $Y2=1.302
r872 281 282 66.1985 $w=2.13e-07 $l=1.235e-06 $layer=LI1_cond $X=4.025 $Y=1.302
+ $X2=2.79 $Y2=1.302
r873 280 320 5.6179 $w=2.8e-07 $l=1.55e-07 $layer=LI1_cond $X=2.71 $Y=2.125
+ $X2=2.555 $Y2=2.125
r874 279 321 6.19399 $w=2.8e-07 $l=1.75e-07 $layer=LI1_cond $X=3.94 $Y=2.125
+ $X2=4.115 $Y2=2.125
r875 279 280 50.6252 $w=2.78e-07 $l=1.23e-06 $layer=LI1_cond $X=3.94 $Y=2.125
+ $X2=2.71 $Y2=2.125
r876 275 277 46.4695 $w=3.08e-07 $l=1.25e-06 $layer=LI1_cond $X=2.555 $Y=2.34
+ $X2=2.555 $Y2=3.59
r877 273 320 0.978733 $w=3.1e-07 $l=1.4e-07 $layer=LI1_cond $X=2.555 $Y=2.265
+ $X2=2.555 $Y2=2.125
r878 273 275 2.78817 $w=3.08e-07 $l=7.5e-08 $layer=LI1_cond $X=2.555 $Y=2.265
+ $X2=2.555 $Y2=2.34
r879 269 319 0.684683 $w=3.9e-07 $l=1.07e-07 $layer=LI1_cond $X=2.595 $Y=1.195
+ $X2=2.595 $Y2=1.302
r880 269 271 8.86495 $w=3.88e-07 $l=3e-07 $layer=LI1_cond $X=2.595 $Y=1.195
+ $X2=2.595 $Y2=0.895
r881 267 319 8.20698 $w=2.15e-07 $l=1.95e-07 $layer=LI1_cond $X=2.4 $Y=1.302
+ $X2=2.595 $Y2=1.302
r882 267 268 65.9305 $w=2.13e-07 $l=1.23e-06 $layer=LI1_cond $X=2.4 $Y=1.302
+ $X2=1.17 $Y2=1.302
r883 265 320 5.6179 $w=2.8e-07 $l=1.55e-07 $layer=LI1_cond $X=2.4 $Y=2.125
+ $X2=2.555 $Y2=2.125
r884 265 266 51.0368 $w=2.78e-07 $l=1.24e-06 $layer=LI1_cond $X=2.4 $Y=2.125
+ $X2=1.16 $Y2=2.125
r885 261 263 46.4695 $w=3.08e-07 $l=1.25e-06 $layer=LI1_cond $X=1.005 $Y=2.34
+ $X2=1.005 $Y2=3.59
r886 259 266 6.83944 $w=2.8e-07 $l=2.13834e-07 $layer=LI1_cond $X=1.005 $Y=2.265
+ $X2=1.16 $Y2=2.125
r887 259 261 2.78817 $w=3.08e-07 $l=7.5e-08 $layer=LI1_cond $X=1.005 $Y=2.265
+ $X2=1.005 $Y2=2.34
r888 255 268 7.36541 $w=2.15e-07 $l=2.25233e-07 $layer=LI1_cond $X=0.992
+ $Y=1.195 $X2=1.17 $Y2=1.302
r889 255 257 8.92738 $w=3.53e-07 $l=2.75e-07 $layer=LI1_cond $X=0.992 $Y=1.195
+ $X2=0.992 $Y2=0.92
r890 248 253 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=32.885 $Y=2.005
+ $X2=32.885 $Y2=2.965
r891 248 250 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=32.885 $Y=1.565
+ $X2=32.885 $Y2=1.08
r892 241 248 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=32.105 $Y=1.785
+ $X2=32.885 $Y2=1.785
r893 241 450 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=32.105 $Y=1.785
+ $X2=31.865 $Y2=1.785
r894 241 246 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=32.105 $Y=2.005
+ $X2=32.105 $Y2=2.965
r895 241 243 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=32.105 $Y=1.565
+ $X2=32.105 $Y2=1.08
r896 234 450 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=31.325 $Y=1.785
+ $X2=31.865 $Y2=1.785
r897 234 239 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=31.325 $Y=2.005
+ $X2=31.325 $Y2=2.965
r898 234 236 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=31.325 $Y=1.565
+ $X2=31.325 $Y2=1.08
r899 227 234 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=30.545 $Y=1.785
+ $X2=31.325 $Y2=1.785
r900 227 445 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=30.545 $Y=1.785
+ $X2=30.305 $Y2=1.785
r901 227 232 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=30.545 $Y=2.005
+ $X2=30.545 $Y2=2.965
r902 227 229 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=30.545 $Y=1.565
+ $X2=30.545 $Y2=1.08
r903 220 445 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=29.765 $Y=1.785
+ $X2=30.305 $Y2=1.785
r904 220 225 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=29.765 $Y=2.005
+ $X2=29.765 $Y2=2.965
r905 220 222 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=29.765 $Y=1.565
+ $X2=29.765 $Y2=1.08
r906 213 220 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=28.985 $Y=1.785
+ $X2=29.765 $Y2=1.785
r907 213 440 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=28.985 $Y=1.785
+ $X2=28.745 $Y2=1.785
r908 213 218 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=28.985 $Y=2.005
+ $X2=28.985 $Y2=2.965
r909 213 215 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=28.985 $Y=1.565
+ $X2=28.985 $Y2=1.08
r910 206 440 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=28.205 $Y=1.785
+ $X2=28.745 $Y2=1.785
r911 206 211 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=28.205 $Y=2.005
+ $X2=28.205 $Y2=2.965
r912 206 208 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=28.205 $Y=1.565
+ $X2=28.205 $Y2=1.08
r913 199 206 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=27.425 $Y=1.785
+ $X2=28.205 $Y2=1.785
r914 199 435 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=27.425 $Y=1.785
+ $X2=27.185 $Y2=1.785
r915 199 204 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=27.425 $Y=2.005
+ $X2=27.425 $Y2=2.965
r916 199 201 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=27.425 $Y=1.565
+ $X2=27.425 $Y2=1.08
r917 192 435 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=26.645 $Y=1.785
+ $X2=27.185 $Y2=1.785
r918 192 197 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=26.645 $Y=2.005
+ $X2=26.645 $Y2=2.965
r919 192 194 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=26.645 $Y=1.565
+ $X2=26.645 $Y2=1.08
r920 185 192 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=25.865 $Y=1.785
+ $X2=26.645 $Y2=1.785
r921 185 430 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=25.865 $Y=1.785
+ $X2=25.625 $Y2=1.785
r922 185 190 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=25.865 $Y=2.005
+ $X2=25.865 $Y2=2.965
r923 185 187 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=25.865 $Y=1.565
+ $X2=25.865 $Y2=1.08
r924 178 430 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=25.085 $Y=1.785
+ $X2=25.625 $Y2=1.785
r925 178 183 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=25.085 $Y=2.005
+ $X2=25.085 $Y2=2.965
r926 178 180 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=25.085 $Y=1.565
+ $X2=25.085 $Y2=1.08
r927 171 178 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=24.305 $Y=1.785
+ $X2=25.085 $Y2=1.785
r928 171 425 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=24.305 $Y=1.785
+ $X2=24.065 $Y2=1.785
r929 171 176 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=24.305 $Y=2.005
+ $X2=24.305 $Y2=2.965
r930 171 173 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=24.305 $Y=1.565
+ $X2=24.305 $Y2=1.08
r931 164 425 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=23.525 $Y=1.785
+ $X2=24.065 $Y2=1.785
r932 164 169 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=23.525 $Y=2.005
+ $X2=23.525 $Y2=2.965
r933 164 166 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=23.525 $Y=1.565
+ $X2=23.525 $Y2=1.08
r934 157 164 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=22.745 $Y=1.785
+ $X2=23.525 $Y2=1.785
r935 157 420 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=22.745 $Y=1.785
+ $X2=22.505 $Y2=1.785
r936 157 162 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=22.745 $Y=2.005
+ $X2=22.745 $Y2=2.965
r937 157 159 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=22.745 $Y=1.565
+ $X2=22.745 $Y2=1.08
r938 150 420 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=21.965 $Y=1.785
+ $X2=22.505 $Y2=1.785
r939 150 155 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=21.965 $Y=2.005
+ $X2=21.965 $Y2=2.965
r940 150 152 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=21.965 $Y=1.565
+ $X2=21.965 $Y2=1.08
r941 143 150 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=21.185 $Y=1.785
+ $X2=21.965 $Y2=1.785
r942 143 415 31.5997 $w=4.4e-07 $l=2.5e-07 $layer=POLY_cond $X=21.185 $Y=1.785
+ $X2=20.935 $Y2=1.785
r943 143 148 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=21.185 $Y=2.005
+ $X2=21.185 $Y2=2.965
r944 143 145 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=21.185 $Y=1.565
+ $X2=21.185 $Y2=1.08
r945 136 415 66.9913 $w=4.4e-07 $l=5.3e-07 $layer=POLY_cond $X=20.405 $Y=1.785
+ $X2=20.935 $Y2=1.785
r946 136 141 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=20.405 $Y=2.005
+ $X2=20.405 $Y2=2.965
r947 136 138 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=20.405 $Y=1.565
+ $X2=20.405 $Y2=1.08
r948 129 136 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=19.625 $Y=1.785
+ $X2=20.405 $Y2=1.785
r949 129 410 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=19.625 $Y=1.785
+ $X2=19.385 $Y2=1.785
r950 129 134 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=19.625 $Y=2.005
+ $X2=19.625 $Y2=2.965
r951 129 131 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=19.625 $Y=1.565
+ $X2=19.625 $Y2=1.08
r952 122 410 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=18.845 $Y=1.785
+ $X2=19.385 $Y2=1.785
r953 122 127 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=18.845 $Y=2.005
+ $X2=18.845 $Y2=2.965
r954 122 124 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=18.845 $Y=1.565
+ $X2=18.845 $Y2=1.08
r955 115 122 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=18.065 $Y=1.785
+ $X2=18.845 $Y2=1.785
r956 115 405 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=18.065 $Y=1.785
+ $X2=17.825 $Y2=1.785
r957 115 120 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=18.065 $Y=2.005
+ $X2=18.065 $Y2=2.965
r958 115 117 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=18.065 $Y=1.565
+ $X2=18.065 $Y2=1.08
r959 108 405 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=17.285 $Y=1.785
+ $X2=17.825 $Y2=1.785
r960 108 113 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=17.285 $Y=2.005
+ $X2=17.285 $Y2=2.965
r961 108 110 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=17.285 $Y=1.565
+ $X2=17.285 $Y2=1.08
r962 101 108 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=16.505 $Y=1.785
+ $X2=17.285 $Y2=1.785
r963 101 400 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=16.505 $Y=1.785
+ $X2=16.265 $Y2=1.785
r964 101 106 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=16.505 $Y=2.005
+ $X2=16.505 $Y2=2.965
r965 101 103 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=16.505 $Y=1.565
+ $X2=16.505 $Y2=1.08
r966 94 400 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=15.725 $Y=1.785
+ $X2=16.265 $Y2=1.785
r967 94 99 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=15.725 $Y=2.005
+ $X2=15.725 $Y2=2.965
r968 94 96 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=15.725 $Y=1.565
+ $X2=15.725 $Y2=1.08
r969 87 94 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=14.945 $Y=1.785
+ $X2=15.725 $Y2=1.785
r970 87 395 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=14.945 $Y=1.785
+ $X2=14.705 $Y2=1.785
r971 87 92 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=14.945 $Y=2.005
+ $X2=14.945 $Y2=2.965
r972 87 89 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=14.945 $Y=1.565
+ $X2=14.945 $Y2=1.08
r973 80 395 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=14.165 $Y=1.785
+ $X2=14.705 $Y2=1.785
r974 80 85 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=14.165 $Y=2.005
+ $X2=14.165 $Y2=2.965
r975 80 82 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=14.165 $Y=1.565
+ $X2=14.165 $Y2=1.08
r976 73 80 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=13.385 $Y=1.785
+ $X2=14.165 $Y2=1.785
r977 73 390 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=13.385 $Y=1.785
+ $X2=13.145 $Y2=1.785
r978 73 78 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=13.385 $Y=2.005
+ $X2=13.385 $Y2=2.965
r979 73 75 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=13.385 $Y=1.565
+ $X2=13.385 $Y2=1.08
r980 66 390 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=12.605 $Y=1.785
+ $X2=13.145 $Y2=1.785
r981 66 71 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=12.605 $Y=2.005
+ $X2=12.605 $Y2=2.965
r982 66 68 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=12.605 $Y=1.565
+ $X2=12.605 $Y2=1.08
r983 59 66 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=11.825 $Y=1.785
+ $X2=12.605 $Y2=1.785
r984 59 385 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=11.825 $Y=1.785
+ $X2=11.585 $Y2=1.785
r985 59 64 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=11.825 $Y=2.005
+ $X2=11.825 $Y2=2.965
r986 59 61 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.825 $Y=1.565
+ $X2=11.825 $Y2=1.08
r987 52 385 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=11.045 $Y=1.785
+ $X2=11.585 $Y2=1.785
r988 52 57 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=11.045 $Y=2.005
+ $X2=11.045 $Y2=2.965
r989 52 54 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.045 $Y=1.565
+ $X2=11.045 $Y2=1.08
r990 45 52 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=10.265 $Y=1.785
+ $X2=11.045 $Y2=1.785
r991 45 380 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=10.265 $Y=1.785
+ $X2=10.025 $Y2=1.785
r992 45 50 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=10.265 $Y=2.005
+ $X2=10.265 $Y2=2.965
r993 45 47 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=10.265 $Y=1.565
+ $X2=10.265 $Y2=1.08
r994 38 380 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=9.485 $Y=1.785
+ $X2=10.025 $Y2=1.785
r995 38 43 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=9.485 $Y=2.005
+ $X2=9.485 $Y2=2.965
r996 38 40 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.485 $Y=1.565
+ $X2=9.485 $Y2=1.08
r997 31 38 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=8.705 $Y=1.785
+ $X2=9.485 $Y2=1.785
r998 31 36 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=8.705 $Y=2.005
+ $X2=8.705 $Y2=2.965
r999 31 33 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=8.705 $Y=1.565
+ $X2=8.705 $Y2=1.08
r1000 10 313 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=7.155
+ $Y=2.215 $X2=7.295 $Y2=3.59
r1001 10 311 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=7.155
+ $Y=2.215 $X2=7.295 $Y2=2.34
r1002 9 305 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=5.595
+ $Y=2.215 $X2=5.735 $Y2=3.59
r1003 9 303 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=5.595
+ $Y=2.215 $X2=5.735 $Y2=2.34
r1004 8 287 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=4.035
+ $Y=2.215 $X2=4.175 $Y2=3.59
r1005 8 285 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.035
+ $Y=2.215 $X2=4.175 $Y2=2.34
r1006 7 277 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.475
+ $Y=2.215 $X2=2.615 $Y2=3.59
r1007 7 275 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.475
+ $Y=2.215 $X2=2.615 $Y2=2.34
r1008 6 263 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=0.915
+ $Y=2.215 $X2=1.055 $Y2=3.59
r1009 6 261 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.915
+ $Y=2.215 $X2=1.055 $Y2=2.34
r1010 5 317 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=7.155
+ $Y=0.705 $X2=7.295 $Y2=0.895
r1011 4 299 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=5.595
+ $Y=0.705 $X2=5.735 $Y2=0.895
r1012 3 291 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=4.035
+ $Y=0.705 $X2=4.175 $Y2=0.895
r1013 2 271 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=2.475
+ $Y=0.705 $X2=2.615 $Y2=0.895
r1014 1 257 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=0.915
+ $Y=0.705 $X2=1.055 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_32%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 17 18 19 20 21 22 67 70 79 90 101 112 123 134 145 156 167 178 189 200 211 219
+ 230 241 252 263 274 285 296 300 336
c331 70 0 3.19988e-20 $X=0.275 $Y=2.36
r332 299 300 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=33.355 $Y=3.56
+ $X2=33.355 $Y2=3.56
r333 296 299 27.081 $w=5.28e-07 $l=1.2e-06 $layer=LI1_cond $X=33.175 $Y=2.36
+ $X2=33.175 $Y2=3.56
r334 291 300 0.491399 $w=3.7e-07 $l=1.28e-06 $layer=MET1_cond $X=32.075 $Y=3.63
+ $X2=33.355 $Y2=3.63
r335 289 291 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=31.355 $Y=3.63
+ $X2=32.075 $Y2=3.63
r336 288 293 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=31.715 $Y=3.56
+ $X2=31.715 $Y2=3.59
r337 288 291 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=32.075 $Y=3.56
+ $X2=32.075 $Y2=3.56
r338 288 289 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=31.355 $Y=3.56
+ $X2=31.355 $Y2=3.56
r339 285 288 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=31.715 $Y=2.34
+ $X2=31.715 $Y2=3.56
r340 280 289 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=30.515 $Y=3.63
+ $X2=31.355 $Y2=3.63
r341 278 280 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=29.795 $Y=3.63
+ $X2=30.515 $Y2=3.63
r342 277 282 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=30.155 $Y=3.56
+ $X2=30.155 $Y2=3.59
r343 277 280 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=30.515 $Y=3.56
+ $X2=30.515 $Y2=3.56
r344 277 278 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=29.795 $Y=3.56
+ $X2=29.795 $Y2=3.56
r345 274 277 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=30.155 $Y=2.34
+ $X2=30.155 $Y2=3.56
r346 269 278 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=28.955 $Y=3.63
+ $X2=29.795 $Y2=3.63
r347 267 269 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=28.235 $Y=3.63
+ $X2=28.955 $Y2=3.63
r348 266 271 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=28.595 $Y=3.56
+ $X2=28.595 $Y2=3.59
r349 266 269 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=28.955 $Y=3.56
+ $X2=28.955 $Y2=3.56
r350 266 267 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=28.235 $Y=3.56
+ $X2=28.235 $Y2=3.56
r351 263 266 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=28.595 $Y=2.34
+ $X2=28.595 $Y2=3.56
r352 258 267 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=27.395 $Y=3.63
+ $X2=28.235 $Y2=3.63
r353 256 258 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=26.675 $Y=3.63
+ $X2=27.395 $Y2=3.63
r354 255 260 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=27.035 $Y=3.56
+ $X2=27.035 $Y2=3.59
r355 255 258 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=27.395 $Y=3.56
+ $X2=27.395 $Y2=3.56
r356 255 256 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=26.675 $Y=3.56
+ $X2=26.675 $Y2=3.56
r357 252 255 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=27.035 $Y=2.34
+ $X2=27.035 $Y2=3.56
r358 247 256 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=25.835 $Y=3.63
+ $X2=26.675 $Y2=3.63
r359 245 247 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=25.115 $Y=3.63
+ $X2=25.835 $Y2=3.63
r360 245 336 0.134367 $w=3.7e-07 $l=3.5e-07 $layer=MET1_cond $X=25.115 $Y=3.63
+ $X2=24.765 $Y2=3.63
r361 244 249 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=25.475 $Y=3.56
+ $X2=25.475 $Y2=3.59
r362 244 247 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=25.835 $Y=3.56
+ $X2=25.835 $Y2=3.56
r363 244 245 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=25.115 $Y=3.56
+ $X2=25.115 $Y2=3.56
r364 241 244 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=25.475 $Y=2.34
+ $X2=25.475 $Y2=3.56
r365 236 336 0.188114 $w=3.7e-07 $l=4.9e-07 $layer=MET1_cond $X=24.275 $Y=3.63
+ $X2=24.765 $Y2=3.63
r366 234 236 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=23.555 $Y=3.63
+ $X2=24.275 $Y2=3.63
r367 233 238 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=23.915 $Y=3.56
+ $X2=23.915 $Y2=3.59
r368 233 236 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=24.275 $Y=3.56
+ $X2=24.275 $Y2=3.56
r369 233 234 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=23.555 $Y=3.56
+ $X2=23.555 $Y2=3.56
r370 230 233 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=23.915 $Y=2.34
+ $X2=23.915 $Y2=3.56
r371 225 234 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=22.715 $Y=3.63
+ $X2=23.555 $Y2=3.63
r372 223 225 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=21.995 $Y=3.63
+ $X2=22.715 $Y2=3.63
r373 222 227 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=22.355 $Y=3.56
+ $X2=22.355 $Y2=3.59
r374 222 225 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=22.715 $Y=3.56
+ $X2=22.715 $Y2=3.56
r375 222 223 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=21.995 $Y=3.56
+ $X2=21.995 $Y2=3.56
r376 219 222 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=22.355 $Y=2.34
+ $X2=22.355 $Y2=3.56
r377 215 223 0.429974 $w=3.7e-07 $l=1.12e-06 $layer=MET1_cond $X=20.875 $Y=3.63
+ $X2=21.995 $Y2=3.63
r378 214 215 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.875 $Y=3.56
+ $X2=20.875 $Y2=3.56
r379 211 214 27.081 $w=5.28e-07 $l=1.2e-06 $layer=LI1_cond $X=20.695 $Y=2.36
+ $X2=20.695 $Y2=3.56
r380 206 215 0.491399 $w=3.7e-07 $l=1.28e-06 $layer=MET1_cond $X=19.595 $Y=3.63
+ $X2=20.875 $Y2=3.63
r381 204 206 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=18.875 $Y=3.63
+ $X2=19.595 $Y2=3.63
r382 203 208 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=19.235 $Y=3.56
+ $X2=19.235 $Y2=3.59
r383 203 206 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=19.595 $Y=3.56
+ $X2=19.595 $Y2=3.56
r384 203 204 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=18.875 $Y=3.56
+ $X2=18.875 $Y2=3.56
r385 200 203 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=19.235 $Y=2.34
+ $X2=19.235 $Y2=3.56
r386 195 204 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=18.035 $Y=3.63
+ $X2=18.875 $Y2=3.63
r387 193 195 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=17.315 $Y=3.63
+ $X2=18.035 $Y2=3.63
r388 192 197 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=17.675 $Y=3.56
+ $X2=17.675 $Y2=3.59
r389 192 195 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=18.035 $Y=3.56
+ $X2=18.035 $Y2=3.56
r390 192 193 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.315 $Y=3.56
+ $X2=17.315 $Y2=3.56
r391 189 192 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=17.675 $Y=2.34
+ $X2=17.675 $Y2=3.56
r392 182 184 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=15.755 $Y=3.63
+ $X2=16.475 $Y2=3.63
r393 181 186 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=16.115 $Y=3.56
+ $X2=16.115 $Y2=3.59
r394 181 184 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.475 $Y=3.56
+ $X2=16.475 $Y2=3.56
r395 181 182 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.755 $Y=3.56
+ $X2=15.755 $Y2=3.56
r396 178 181 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=16.115 $Y=2.34
+ $X2=16.115 $Y2=3.56
r397 173 182 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=14.915 $Y=3.63
+ $X2=15.755 $Y2=3.63
r398 171 173 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=14.195 $Y=3.63
+ $X2=14.915 $Y2=3.63
r399 170 175 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=14.555 $Y=3.56
+ $X2=14.555 $Y2=3.59
r400 170 173 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.915 $Y=3.56
+ $X2=14.915 $Y2=3.56
r401 170 171 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.195 $Y=3.56
+ $X2=14.195 $Y2=3.56
r402 167 170 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=14.555 $Y=2.34
+ $X2=14.555 $Y2=3.56
r403 162 171 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=13.355 $Y=3.63
+ $X2=14.195 $Y2=3.63
r404 160 162 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=12.635 $Y=3.63
+ $X2=13.355 $Y2=3.63
r405 159 164 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=12.995 $Y=3.56
+ $X2=12.995 $Y2=3.59
r406 159 162 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.355 $Y=3.56
+ $X2=13.355 $Y2=3.56
r407 159 160 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.635 $Y=3.56
+ $X2=12.635 $Y2=3.56
r408 156 159 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=12.995 $Y=2.34
+ $X2=12.995 $Y2=3.56
r409 151 160 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=11.795 $Y=3.63
+ $X2=12.635 $Y2=3.63
r410 149 151 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=11.075 $Y=3.63
+ $X2=11.795 $Y2=3.63
r411 148 153 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=11.435 $Y=3.56
+ $X2=11.435 $Y2=3.59
r412 148 151 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.795 $Y=3.56
+ $X2=11.795 $Y2=3.56
r413 148 149 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.075 $Y=3.56
+ $X2=11.075 $Y2=3.56
r414 145 148 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=11.435 $Y=2.34
+ $X2=11.435 $Y2=3.56
r415 140 149 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=10.235 $Y=3.63
+ $X2=11.075 $Y2=3.63
r416 138 140 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=9.515 $Y=3.63
+ $X2=10.235 $Y2=3.63
r417 137 142 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=9.875 $Y=3.56
+ $X2=9.875 $Y2=3.59
r418 137 140 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.235 $Y=3.56
+ $X2=10.235 $Y2=3.56
r419 137 138 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.515 $Y=3.56
+ $X2=9.515 $Y2=3.56
r420 134 137 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=9.875 $Y=2.34
+ $X2=9.875 $Y2=3.56
r421 129 138 0.433813 $w=3.7e-07 $l=1.13e-06 $layer=MET1_cond $X=8.385 $Y=3.63
+ $X2=9.515 $Y2=3.63
r422 127 129 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.665 $Y=3.63
+ $X2=8.385 $Y2=3.63
r423 126 131 0.135556 $w=8.98e-07 $l=1e-08 $layer=LI1_cond $X=8.03 $Y=3.56
+ $X2=8.03 $Y2=3.57
r424 126 129 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.385 $Y=3.56
+ $X2=8.385 $Y2=3.56
r425 126 127 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.665 $Y=3.56
+ $X2=7.665 $Y2=3.56
r426 123 126 16.5378 $w=8.98e-07 $l=1.22e-06 $layer=LI1_cond $X=8.03 $Y=2.34
+ $X2=8.03 $Y2=3.56
r427 118 127 0.330159 $w=3.7e-07 $l=8.6e-07 $layer=MET1_cond $X=6.805 $Y=3.63
+ $X2=7.665 $Y2=3.63
r428 116 118 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=6.085 $Y=3.63
+ $X2=6.805 $Y2=3.63
r429 115 120 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=6.445 $Y=3.56
+ $X2=6.445 $Y2=3.57
r430 115 118 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.805 $Y=3.56
+ $X2=6.805 $Y2=3.56
r431 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.085 $Y=3.56
+ $X2=6.085 $Y2=3.56
r432 112 115 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=6.445 $Y=2.55
+ $X2=6.445 $Y2=3.56
r433 107 116 0.314802 $w=3.7e-07 $l=8.2e-07 $layer=MET1_cond $X=5.265 $Y=3.63
+ $X2=6.085 $Y2=3.63
r434 105 107 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=4.545 $Y=3.63
+ $X2=5.265 $Y2=3.63
r435 104 109 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=4.905 $Y=3.56
+ $X2=4.905 $Y2=3.57
r436 104 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.265 $Y=3.56
+ $X2=5.265 $Y2=3.56
r437 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.545 $Y=3.56
+ $X2=4.545 $Y2=3.56
r438 101 104 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=4.905 $Y=2.55
+ $X2=4.905 $Y2=3.56
r439 96 105 0.330159 $w=3.7e-07 $l=8.6e-07 $layer=MET1_cond $X=3.685 $Y=3.63
+ $X2=4.545 $Y2=3.63
r440 94 96 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.965 $Y=3.63
+ $X2=3.685 $Y2=3.63
r441 93 98 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=3.325 $Y=3.56
+ $X2=3.325 $Y2=3.57
r442 93 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.685 $Y=3.56
+ $X2=3.685 $Y2=3.56
r443 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.965 $Y=3.56
+ $X2=2.965 $Y2=3.56
r444 90 93 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=3.325 $Y=2.55
+ $X2=3.325 $Y2=3.56
r445 85 94 0.314802 $w=3.7e-07 $l=8.2e-07 $layer=MET1_cond $X=2.145 $Y=3.63
+ $X2=2.965 $Y2=3.63
r446 83 85 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.425 $Y=3.63
+ $X2=2.145 $Y2=3.63
r447 82 87 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=1.785 $Y=3.56
+ $X2=1.785 $Y2=3.57
r448 82 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.145 $Y=3.56
+ $X2=2.145 $Y2=3.56
r449 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.425 $Y=3.56
+ $X2=1.425 $Y2=3.56
r450 79 82 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=1.785 $Y=2.55
+ $X2=1.785 $Y2=3.56
r451 74 83 0.318641 $w=3.7e-07 $l=8.3e-07 $layer=MET1_cond $X=0.595 $Y=3.63
+ $X2=1.425 $Y2=3.63
r452 73 76 0.209838 $w=5.68e-07 $l=1e-08 $layer=LI1_cond $X=0.395 $Y=3.56
+ $X2=0.395 $Y2=3.57
r453 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.595 $Y=3.56
+ $X2=0.595 $Y2=3.56
r454 70 73 25.1806 $w=5.68e-07 $l=1.2e-06 $layer=LI1_cond $X=0.395 $Y=2.36
+ $X2=0.395 $Y2=3.56
r455 67 193 0.197711 $w=3.7e-07 $l=5.15e-07 $layer=MET1_cond $X=16.8 $Y=3.63
+ $X2=17.315 $Y2=3.63
r456 67 184 0.124769 $w=3.7e-07 $l=3.25e-07 $layer=MET1_cond $X=16.8 $Y=3.63
+ $X2=16.475 $Y2=3.63
r457 22 299 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=33.135
+ $Y=2.215 $X2=33.275 $Y2=3.57
r458 22 296 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=33.135
+ $Y=2.215 $X2=33.275 $Y2=2.36
r459 21 293 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=31.575
+ $Y=2.215 $X2=31.715 $Y2=3.59
r460 21 285 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=31.575
+ $Y=2.215 $X2=31.715 $Y2=2.34
r461 20 282 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=30.015
+ $Y=2.215 $X2=30.155 $Y2=3.59
r462 20 274 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=30.015
+ $Y=2.215 $X2=30.155 $Y2=2.34
r463 19 271 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=28.455
+ $Y=2.215 $X2=28.595 $Y2=3.59
r464 19 263 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=28.455
+ $Y=2.215 $X2=28.595 $Y2=2.34
r465 18 260 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=26.895
+ $Y=2.215 $X2=27.035 $Y2=3.59
r466 18 252 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=26.895
+ $Y=2.215 $X2=27.035 $Y2=2.34
r467 17 249 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=25.335
+ $Y=2.215 $X2=25.475 $Y2=3.59
r468 17 241 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=25.335
+ $Y=2.215 $X2=25.475 $Y2=2.34
r469 16 238 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=23.775
+ $Y=2.215 $X2=23.915 $Y2=3.59
r470 16 230 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=23.775
+ $Y=2.215 $X2=23.915 $Y2=2.34
r471 15 227 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=22.215
+ $Y=2.215 $X2=22.355 $Y2=3.59
r472 15 219 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=22.215
+ $Y=2.215 $X2=22.355 $Y2=2.34
r473 14 214 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=20.655
+ $Y=2.215 $X2=20.795 $Y2=3.57
r474 14 211 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=20.655
+ $Y=2.215 $X2=20.795 $Y2=2.36
r475 13 208 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=19.095
+ $Y=2.215 $X2=19.235 $Y2=3.59
r476 13 200 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=19.095
+ $Y=2.215 $X2=19.235 $Y2=2.34
r477 12 197 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=17.535
+ $Y=2.215 $X2=17.675 $Y2=3.59
r478 12 189 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=17.535
+ $Y=2.215 $X2=17.675 $Y2=2.34
r479 11 186 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=15.975
+ $Y=2.215 $X2=16.115 $Y2=3.59
r480 11 178 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=15.975
+ $Y=2.215 $X2=16.115 $Y2=2.34
r481 10 175 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=14.415
+ $Y=2.215 $X2=14.555 $Y2=3.59
r482 10 167 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=14.415
+ $Y=2.215 $X2=14.555 $Y2=2.34
r483 9 164 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=12.855
+ $Y=2.215 $X2=12.995 $Y2=3.59
r484 9 156 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=12.855
+ $Y=2.215 $X2=12.995 $Y2=2.34
r485 8 153 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=11.295
+ $Y=2.215 $X2=11.435 $Y2=3.59
r486 8 145 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=11.295
+ $Y=2.215 $X2=11.435 $Y2=2.34
r487 7 142 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=9.735
+ $Y=2.215 $X2=9.875 $Y2=3.59
r488 7 134 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=9.735
+ $Y=2.215 $X2=9.875 $Y2=2.34
r489 6 131 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=7.935
+ $Y=2.215 $X2=8.075 $Y2=3.57
r490 6 123 300 $w=1.7e-07 $l=4.38064e-07 $layer=licon1_PDIFF $count=2 $X=7.935
+ $Y=2.215 $X2=8.315 $Y2=2.34
r491 5 120 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=6.375
+ $Y=2.215 $X2=6.515 $Y2=3.57
r492 5 112 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=6.375
+ $Y=2.215 $X2=6.515 $Y2=2.55
r493 4 109 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=2.215 $X2=4.955 $Y2=3.57
r494 4 101 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=2.215 $X2=4.955 $Y2=2.55
r495 3 98 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=3.255
+ $Y=2.215 $X2=3.395 $Y2=3.57
r496 3 90 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=3.255
+ $Y=2.215 $X2=3.395 $Y2=2.55
r497 2 87 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=2.215 $X2=1.835 $Y2=3.57
r498 2 79 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=2.215 $X2=1.835 $Y2=2.55
r499 1 76 300 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.215 $X2=0.275 $Y2=3.57
r500 1 70 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.215 $X2=0.275 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_32%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17
+ 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 97 100 110 120 130 140 150 160
+ 170 180 190 200 210 220 230 240 250 255 270
r334 253 257 35.1355 $w=4.08e-07 $l=1.25e-06 $layer=LI1_cond $X=32.535 $Y=2.34
+ $X2=32.535 $Y2=3.59
r335 253 255 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=32.495 $Y=2.405
+ $X2=32.495 $Y2=2.405
r336 250 253 38.9301 $w=4.08e-07 $l=1.385e-06 $layer=LI1_cond $X=32.535 $Y=0.955
+ $X2=32.535 $Y2=2.34
r337 245 255 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=30.935 $Y=2.405
+ $X2=32.495 $Y2=2.405
r338 243 247 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=30.935 $Y=2.34
+ $X2=30.935 $Y2=3.59
r339 243 245 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=30.935 $Y=2.405
+ $X2=30.935 $Y2=2.405
r340 240 243 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=30.935 $Y=0.955
+ $X2=30.935 $Y2=2.34
r341 235 245 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=29.375 $Y=2.405
+ $X2=30.935 $Y2=2.405
r342 233 237 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=29.375 $Y=2.34
+ $X2=29.375 $Y2=3.59
r343 233 235 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=29.375 $Y=2.405
+ $X2=29.375 $Y2=2.405
r344 230 233 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=29.375 $Y=0.955
+ $X2=29.375 $Y2=2.34
r345 225 235 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=27.815 $Y=2.405
+ $X2=29.375 $Y2=2.405
r346 223 227 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=27.815 $Y=2.34
+ $X2=27.815 $Y2=3.59
r347 223 225 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=27.815 $Y=2.405
+ $X2=27.815 $Y2=2.405
r348 220 223 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=27.815 $Y=0.955
+ $X2=27.815 $Y2=2.34
r349 215 225 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=26.255 $Y=2.405
+ $X2=27.815 $Y2=2.405
r350 213 217 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=26.255 $Y=2.34
+ $X2=26.255 $Y2=3.59
r351 213 215 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=26.255 $Y=2.405
+ $X2=26.255 $Y2=2.405
r352 210 213 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=26.255 $Y=0.955
+ $X2=26.255 $Y2=2.34
r353 205 215 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=24.695 $Y=2.405
+ $X2=26.255 $Y2=2.405
r354 203 207 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=24.695 $Y=2.34
+ $X2=24.695 $Y2=3.59
r355 203 205 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.695 $Y=2.405
+ $X2=24.695 $Y2=2.405
r356 200 203 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=24.695 $Y=0.955
+ $X2=24.695 $Y2=2.34
r357 195 205 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=23.135 $Y=2.405
+ $X2=24.695 $Y2=2.405
r358 193 197 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=23.135 $Y=2.34
+ $X2=23.135 $Y2=3.59
r359 193 195 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=23.135 $Y=2.405
+ $X2=23.135 $Y2=2.405
r360 190 193 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=23.135 $Y=0.955
+ $X2=23.135 $Y2=2.34
r361 185 195 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=21.575 $Y=2.405
+ $X2=23.135 $Y2=2.405
r362 185 270 0.343258 $w=2.3e-07 $l=5.35e-07 $layer=MET1_cond $X=21.575 $Y=2.405
+ $X2=21.04 $Y2=2.405
r363 183 187 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=21.575 $Y=2.34
+ $X2=21.575 $Y2=3.59
r364 183 185 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.575 $Y=2.405
+ $X2=21.575 $Y2=2.405
r365 180 183 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=21.575 $Y=0.955
+ $X2=21.575 $Y2=2.34
r366 173 177 35.1355 $w=4.08e-07 $l=1.25e-06 $layer=LI1_cond $X=20.055 $Y=2.34
+ $X2=20.055 $Y2=3.59
r367 173 175 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.015 $Y=2.405
+ $X2=20.015 $Y2=2.405
r368 170 173 38.9301 $w=4.08e-07 $l=1.385e-06 $layer=LI1_cond $X=20.055 $Y=0.955
+ $X2=20.055 $Y2=2.34
r369 165 175 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=18.455 $Y=2.405
+ $X2=20.015 $Y2=2.405
r370 163 167 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=18.455 $Y=2.34
+ $X2=18.455 $Y2=3.59
r371 163 165 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.455 $Y=2.405
+ $X2=18.455 $Y2=2.405
r372 160 163 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=18.455 $Y=0.955
+ $X2=18.455 $Y2=2.34
r373 155 165 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=16.895 $Y=2.405
+ $X2=18.455 $Y2=2.405
r374 153 157 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=16.895 $Y=2.34
+ $X2=16.895 $Y2=3.59
r375 153 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.895 $Y=2.405
+ $X2=16.895 $Y2=2.405
r376 150 153 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=16.895 $Y=0.955
+ $X2=16.895 $Y2=2.34
r377 145 155 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=15.335 $Y=2.405
+ $X2=16.895 $Y2=2.405
r378 143 147 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=15.335 $Y=2.34
+ $X2=15.335 $Y2=3.59
r379 143 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.335 $Y=2.405
+ $X2=15.335 $Y2=2.405
r380 140 143 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=15.335 $Y=0.955
+ $X2=15.335 $Y2=2.34
r381 135 145 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=13.775 $Y=2.405
+ $X2=15.335 $Y2=2.405
r382 133 137 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=13.775 $Y=2.34
+ $X2=13.775 $Y2=3.59
r383 133 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.775 $Y=2.405
+ $X2=13.775 $Y2=2.405
r384 130 133 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=13.775 $Y=0.955
+ $X2=13.775 $Y2=2.34
r385 125 135 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=12.215 $Y=2.405
+ $X2=13.775 $Y2=2.405
r386 123 127 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=12.215 $Y=2.34
+ $X2=12.215 $Y2=3.59
r387 123 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.215 $Y=2.405
+ $X2=12.215 $Y2=2.405
r388 120 123 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=12.215 $Y=0.955
+ $X2=12.215 $Y2=2.34
r389 115 125 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=10.655 $Y=2.405
+ $X2=12.215 $Y2=2.405
r390 113 117 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=10.655 $Y=2.34
+ $X2=10.655 $Y2=3.59
r391 113 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.655 $Y=2.405
+ $X2=10.655 $Y2=2.405
r392 110 113 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=10.655 $Y=0.955
+ $X2=10.655 $Y2=2.34
r393 105 115 1.0009 $w=2.3e-07 $l=1.56e-06 $layer=MET1_cond $X=9.095 $Y=2.405
+ $X2=10.655 $Y2=2.405
r394 103 107 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=9.095 $Y=2.34
+ $X2=9.095 $Y2=3.59
r395 103 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.095 $Y=2.405
+ $X2=9.095 $Y2=2.405
r396 100 103 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=9.095 $Y=0.955
+ $X2=9.095 $Y2=2.34
r397 97 270 0.157193 $w=2.3e-07 $l=2.45e-07 $layer=MET1_cond $X=20.795 $Y=2.405
+ $X2=21.04 $Y2=2.405
r398 97 175 0.500451 $w=2.3e-07 $l=7.8e-07 $layer=MET1_cond $X=20.795 $Y=2.405
+ $X2=20.015 $Y2=2.405
r399 32 257 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=32.355
+ $Y=2.215 $X2=32.495 $Y2=3.59
r400 32 253 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=32.355
+ $Y=2.215 $X2=32.495 $Y2=2.34
r401 31 247 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=30.795
+ $Y=2.215 $X2=30.935 $Y2=3.59
r402 31 243 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=30.795
+ $Y=2.215 $X2=30.935 $Y2=2.34
r403 30 237 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=29.235
+ $Y=2.215 $X2=29.375 $Y2=3.59
r404 30 233 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=29.235
+ $Y=2.215 $X2=29.375 $Y2=2.34
r405 29 227 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=27.675
+ $Y=2.215 $X2=27.815 $Y2=3.59
r406 29 223 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=27.675
+ $Y=2.215 $X2=27.815 $Y2=2.34
r407 28 217 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=26.115
+ $Y=2.215 $X2=26.255 $Y2=3.59
r408 28 213 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=26.115
+ $Y=2.215 $X2=26.255 $Y2=2.34
r409 27 207 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=24.555
+ $Y=2.215 $X2=24.695 $Y2=3.59
r410 27 203 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=24.555
+ $Y=2.215 $X2=24.695 $Y2=2.34
r411 26 197 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=22.995
+ $Y=2.215 $X2=23.135 $Y2=3.59
r412 26 193 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=22.995
+ $Y=2.215 $X2=23.135 $Y2=2.34
r413 25 187 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=21.435
+ $Y=2.215 $X2=21.575 $Y2=3.59
r414 25 183 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=21.435
+ $Y=2.215 $X2=21.575 $Y2=2.34
r415 24 177 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=19.875
+ $Y=2.215 $X2=20.015 $Y2=3.59
r416 24 173 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=19.875
+ $Y=2.215 $X2=20.015 $Y2=2.34
r417 23 167 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=18.315
+ $Y=2.215 $X2=18.455 $Y2=3.59
r418 23 163 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=18.315
+ $Y=2.215 $X2=18.455 $Y2=2.34
r419 22 157 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=16.755
+ $Y=2.215 $X2=16.895 $Y2=3.59
r420 22 153 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=16.755
+ $Y=2.215 $X2=16.895 $Y2=2.34
r421 21 147 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=15.195
+ $Y=2.215 $X2=15.335 $Y2=3.59
r422 21 143 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=15.195
+ $Y=2.215 $X2=15.335 $Y2=2.34
r423 20 137 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=13.635
+ $Y=2.215 $X2=13.775 $Y2=3.59
r424 20 133 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=13.635
+ $Y=2.215 $X2=13.775 $Y2=2.34
r425 19 127 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=12.075
+ $Y=2.215 $X2=12.215 $Y2=3.59
r426 19 123 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=12.075
+ $Y=2.215 $X2=12.215 $Y2=2.34
r427 18 117 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=10.515
+ $Y=2.215 $X2=10.655 $Y2=3.59
r428 18 113 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=10.515
+ $Y=2.215 $X2=10.655 $Y2=2.34
r429 17 107 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=8.955
+ $Y=2.215 $X2=9.095 $Y2=3.59
r430 17 103 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=8.955
+ $Y=2.215 $X2=9.095 $Y2=2.34
r431 16 250 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=32.355
+ $Y=0.705 $X2=32.495 $Y2=0.955
r432 15 240 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=30.795
+ $Y=0.705 $X2=30.935 $Y2=0.955
r433 14 230 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=29.235
+ $Y=0.705 $X2=29.375 $Y2=0.955
r434 13 220 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=27.675
+ $Y=0.705 $X2=27.815 $Y2=0.955
r435 12 210 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=26.115
+ $Y=0.705 $X2=26.255 $Y2=0.955
r436 11 200 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=24.555
+ $Y=0.705 $X2=24.695 $Y2=0.955
r437 10 190 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=22.995
+ $Y=0.705 $X2=23.135 $Y2=0.955
r438 9 180 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=21.435
+ $Y=0.705 $X2=21.575 $Y2=0.955
r439 8 170 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=19.875
+ $Y=0.705 $X2=20.015 $Y2=0.955
r440 7 160 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=18.315
+ $Y=0.705 $X2=18.455 $Y2=0.955
r441 6 150 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=16.755
+ $Y=0.705 $X2=16.895 $Y2=0.955
r442 5 140 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=15.195
+ $Y=0.705 $X2=15.335 $Y2=0.955
r443 4 130 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=13.635
+ $Y=0.705 $X2=13.775 $Y2=0.955
r444 3 120 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=12.075
+ $Y=0.705 $X2=12.215 $Y2=0.955
r445 2 110 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=10.515
+ $Y=0.705 $X2=10.655 $Y2=0.955
r446 1 100 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=8.955
+ $Y=0.705 $X2=9.095 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_32%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 17 18 19 20 21 22 67 70 77 86 95 104 113 122 131 140 149 158 167 176 183 192
+ 201 210 219 228 237 246 247 253 292
r298 254 256 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.645 $Y=0.44
+ $X2=8.365 $Y2=0.44
r299 253 258 5.48465 $w=9.12e-07 $l=4.1e-07 $layer=LI1_cond $X=8.02 $Y=0.51
+ $X2=8.02 $Y2=0.92
r300 253 256 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.365 $Y=0.51
+ $X2=8.365 $Y2=0.51
r301 253 254 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.645 $Y=0.51
+ $X2=7.645 $Y2=0.51
r302 246 250 10.0425 $w=5.28e-07 $l=4.45e-07 $layer=LI1_cond $X=33.175 $Y=0.51
+ $X2=33.175 $Y2=0.955
r303 246 247 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=33.355 $Y=0.51
+ $X2=33.355 $Y2=0.51
r304 241 247 0.491399 $w=3.7e-07 $l=1.28e-06 $layer=MET1_cond $X=32.075 $Y=0.44
+ $X2=33.355 $Y2=0.44
r305 238 241 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=31.355 $Y=0.44
+ $X2=32.075 $Y2=0.44
r306 237 243 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=31.715 $Y=0.51
+ $X2=31.715 $Y2=0.92
r307 237 241 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=32.075 $Y=0.51
+ $X2=32.075 $Y2=0.51
r308 237 238 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=31.355 $Y=0.51
+ $X2=31.355 $Y2=0.51
r309 232 238 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=30.515 $Y=0.44
+ $X2=31.355 $Y2=0.44
r310 229 232 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=29.795 $Y=0.44
+ $X2=30.515 $Y2=0.44
r311 228 234 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=30.155 $Y=0.51
+ $X2=30.155 $Y2=0.92
r312 228 232 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=30.515 $Y=0.51
+ $X2=30.515 $Y2=0.51
r313 228 229 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=29.795 $Y=0.51
+ $X2=29.795 $Y2=0.51
r314 223 229 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=28.955 $Y=0.44
+ $X2=29.795 $Y2=0.44
r315 220 223 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=28.235 $Y=0.44
+ $X2=28.955 $Y2=0.44
r316 219 225 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=28.595 $Y=0.51
+ $X2=28.595 $Y2=0.92
r317 219 223 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=28.955 $Y=0.51
+ $X2=28.955 $Y2=0.51
r318 219 220 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=28.235 $Y=0.51
+ $X2=28.235 $Y2=0.51
r319 214 220 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=27.395 $Y=0.44
+ $X2=28.235 $Y2=0.44
r320 211 214 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=26.675 $Y=0.44
+ $X2=27.395 $Y2=0.44
r321 210 216 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=27.035 $Y=0.51
+ $X2=27.035 $Y2=0.92
r322 210 214 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=27.395 $Y=0.51
+ $X2=27.395 $Y2=0.51
r323 210 211 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=26.675 $Y=0.51
+ $X2=26.675 $Y2=0.51
r324 205 211 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=25.835 $Y=0.44
+ $X2=26.675 $Y2=0.44
r325 202 205 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=25.115 $Y=0.44
+ $X2=25.835 $Y2=0.44
r326 202 292 0.134367 $w=3.7e-07 $l=3.5e-07 $layer=MET1_cond $X=25.115 $Y=0.44
+ $X2=24.765 $Y2=0.44
r327 201 207 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=25.475 $Y=0.51
+ $X2=25.475 $Y2=0.92
r328 201 205 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=25.835 $Y=0.51
+ $X2=25.835 $Y2=0.51
r329 201 202 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=25.115 $Y=0.51
+ $X2=25.115 $Y2=0.51
r330 196 292 0.188114 $w=3.7e-07 $l=4.9e-07 $layer=MET1_cond $X=24.275 $Y=0.44
+ $X2=24.765 $Y2=0.44
r331 193 196 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=23.555 $Y=0.44
+ $X2=24.275 $Y2=0.44
r332 192 198 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=23.915 $Y=0.51
+ $X2=23.915 $Y2=0.92
r333 192 196 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=24.275 $Y=0.51
+ $X2=24.275 $Y2=0.51
r334 192 193 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=23.555 $Y=0.51
+ $X2=23.555 $Y2=0.51
r335 187 193 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=22.715 $Y=0.44
+ $X2=23.555 $Y2=0.44
r336 184 187 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=21.995 $Y=0.44
+ $X2=22.715 $Y2=0.44
r337 183 189 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=22.355 $Y=0.51
+ $X2=22.355 $Y2=0.92
r338 183 187 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=22.715 $Y=0.51
+ $X2=22.715 $Y2=0.51
r339 183 184 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=21.995 $Y=0.51
+ $X2=21.995 $Y2=0.51
r340 177 184 0.429974 $w=3.7e-07 $l=1.12e-06 $layer=MET1_cond $X=20.875 $Y=0.44
+ $X2=21.995 $Y2=0.44
r341 176 180 8.91417 $w=5.28e-07 $l=3.95e-07 $layer=LI1_cond $X=20.695 $Y=0.51
+ $X2=20.695 $Y2=0.905
r342 176 177 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.875 $Y=0.51
+ $X2=20.875 $Y2=0.51
r343 171 177 0.491399 $w=3.7e-07 $l=1.28e-06 $layer=MET1_cond $X=19.595 $Y=0.44
+ $X2=20.875 $Y2=0.44
r344 168 171 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=18.875 $Y=0.44
+ $X2=19.595 $Y2=0.44
r345 167 173 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=19.235 $Y=0.51
+ $X2=19.235 $Y2=0.92
r346 167 171 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=19.595 $Y=0.51
+ $X2=19.595 $Y2=0.51
r347 167 168 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=18.875 $Y=0.51
+ $X2=18.875 $Y2=0.51
r348 162 168 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=18.035 $Y=0.44
+ $X2=18.875 $Y2=0.44
r349 159 162 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=17.315 $Y=0.44
+ $X2=18.035 $Y2=0.44
r350 158 164 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=17.675 $Y=0.51
+ $X2=17.675 $Y2=0.92
r351 158 162 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=18.035 $Y=0.51
+ $X2=18.035 $Y2=0.51
r352 158 159 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.315 $Y=0.51
+ $X2=17.315 $Y2=0.51
r353 150 153 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=15.755 $Y=0.44
+ $X2=16.475 $Y2=0.44
r354 149 155 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=16.115 $Y=0.51
+ $X2=16.115 $Y2=0.92
r355 149 153 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.475 $Y=0.51
+ $X2=16.475 $Y2=0.51
r356 149 150 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.755 $Y=0.51
+ $X2=15.755 $Y2=0.51
r357 144 150 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=14.915 $Y=0.44
+ $X2=15.755 $Y2=0.44
r358 141 144 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=14.195 $Y=0.44
+ $X2=14.915 $Y2=0.44
r359 140 146 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=14.555 $Y=0.51
+ $X2=14.555 $Y2=0.92
r360 140 144 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.915 $Y=0.51
+ $X2=14.915 $Y2=0.51
r361 140 141 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.195 $Y=0.51
+ $X2=14.195 $Y2=0.51
r362 135 141 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=13.355 $Y=0.44
+ $X2=14.195 $Y2=0.44
r363 132 135 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=12.635 $Y=0.44
+ $X2=13.355 $Y2=0.44
r364 131 137 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=12.995 $Y=0.51
+ $X2=12.995 $Y2=0.92
r365 131 135 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.355 $Y=0.51
+ $X2=13.355 $Y2=0.51
r366 131 132 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.635 $Y=0.51
+ $X2=12.635 $Y2=0.51
r367 126 132 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=11.795 $Y=0.44
+ $X2=12.635 $Y2=0.44
r368 123 126 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=11.075 $Y=0.44
+ $X2=11.795 $Y2=0.44
r369 122 128 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=11.435 $Y=0.51
+ $X2=11.435 $Y2=0.92
r370 122 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.795 $Y=0.51
+ $X2=11.795 $Y2=0.51
r371 122 123 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.075 $Y=0.51
+ $X2=11.075 $Y2=0.51
r372 117 123 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=10.235 $Y=0.44
+ $X2=11.075 $Y2=0.44
r373 114 117 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=9.515 $Y=0.44
+ $X2=10.235 $Y2=0.44
r374 114 256 0.441491 $w=3.7e-07 $l=1.15e-06 $layer=MET1_cond $X=9.515 $Y=0.44
+ $X2=8.365 $Y2=0.44
r375 113 119 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=9.875 $Y=0.51
+ $X2=9.875 $Y2=0.92
r376 113 117 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.235 $Y=0.51
+ $X2=10.235 $Y2=0.51
r377 113 114 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.515 $Y=0.51
+ $X2=9.515 $Y2=0.51
r378 108 254 0.291768 $w=3.7e-07 $l=7.6e-07 $layer=MET1_cond $X=6.885 $Y=0.44
+ $X2=7.645 $Y2=0.44
r379 105 108 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=6.165 $Y=0.44
+ $X2=6.885 $Y2=0.44
r380 104 110 5.86145 $w=8.93e-07 $l=4.3e-07 $layer=LI1_cond $X=6.527 $Y=0.51
+ $X2=6.527 $Y2=0.94
r381 104 108 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.885 $Y=0.51
+ $X2=6.885 $Y2=0.51
r382 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.165 $Y=0.51
+ $X2=6.165 $Y2=0.51
r383 99 105 0.353193 $w=3.7e-07 $l=9.2e-07 $layer=MET1_cond $X=5.245 $Y=0.44
+ $X2=6.165 $Y2=0.44
r384 96 99 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=4.525 $Y=0.44
+ $X2=5.245 $Y2=0.44
r385 95 101 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=4.885 $Y=0.51
+ $X2=4.885 $Y2=0.92
r386 95 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.245 $Y=0.51
+ $X2=5.245 $Y2=0.51
r387 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.525 $Y=0.51
+ $X2=4.525 $Y2=0.51
r388 90 96 0.291768 $w=3.7e-07 $l=7.6e-07 $layer=MET1_cond $X=3.765 $Y=0.44
+ $X2=4.525 $Y2=0.44
r389 87 90 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.045 $Y=0.44
+ $X2=3.765 $Y2=0.44
r390 86 92 5.86145 $w=8.93e-07 $l=4.3e-07 $layer=LI1_cond $X=3.407 $Y=0.51
+ $X2=3.407 $Y2=0.94
r391 86 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.765 $Y=0.51
+ $X2=3.765 $Y2=0.51
r392 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.045 $Y=0.51
+ $X2=3.045 $Y2=0.51
r393 81 87 0.345515 $w=3.7e-07 $l=9e-07 $layer=MET1_cond $X=2.145 $Y=0.44
+ $X2=3.045 $Y2=0.44
r394 78 81 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.425 $Y=0.44
+ $X2=2.145 $Y2=0.44
r395 77 83 5.89438 $w=8.88e-07 $l=4.3e-07 $layer=LI1_cond $X=1.785 $Y=0.51
+ $X2=1.785 $Y2=0.94
r396 77 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.145 $Y=0.51
+ $X2=2.145 $Y2=0.51
r397 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.425 $Y=0.51
+ $X2=1.425 $Y2=0.51
r398 71 78 0.332078 $w=3.7e-07 $l=8.65e-07 $layer=MET1_cond $X=0.56 $Y=0.44
+ $X2=1.425 $Y2=0.44
r399 70 74 9.61334 $w=5.33e-07 $l=4.3e-07 $layer=LI1_cond $X=0.377 $Y=0.51
+ $X2=0.377 $Y2=0.94
r400 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.56 $Y=0.51
+ $X2=0.56 $Y2=0.51
r401 67 159 0.197711 $w=3.7e-07 $l=5.15e-07 $layer=MET1_cond $X=16.8 $Y=0.44
+ $X2=17.315 $Y2=0.44
r402 67 153 0.124769 $w=3.7e-07 $l=3.25e-07 $layer=MET1_cond $X=16.8 $Y=0.44
+ $X2=16.475 $Y2=0.44
r403 22 250 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=33.135
+ $Y=0.705 $X2=33.275 $Y2=0.955
r404 21 243 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=31.575
+ $Y=0.705 $X2=31.715 $Y2=0.92
r405 20 234 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=30.015
+ $Y=0.705 $X2=30.155 $Y2=0.92
r406 19 225 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=28.455
+ $Y=0.705 $X2=28.595 $Y2=0.92
r407 18 216 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=26.895
+ $Y=0.705 $X2=27.035 $Y2=0.92
r408 17 207 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=25.335
+ $Y=0.705 $X2=25.475 $Y2=0.92
r409 16 198 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=23.775
+ $Y=0.705 $X2=23.915 $Y2=0.92
r410 15 189 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=22.215
+ $Y=0.705 $X2=22.355 $Y2=0.92
r411 14 180 91 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=2 $X=20.655
+ $Y=0.705 $X2=20.795 $Y2=0.905
r412 13 173 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=19.095
+ $Y=0.705 $X2=19.235 $Y2=0.92
r413 12 164 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=17.535
+ $Y=0.705 $X2=17.675 $Y2=0.92
r414 11 155 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=15.975
+ $Y=0.705 $X2=16.115 $Y2=0.92
r415 10 146 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=14.415
+ $Y=0.705 $X2=14.555 $Y2=0.92
r416 9 137 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=12.855
+ $Y=0.705 $X2=12.995 $Y2=0.92
r417 8 128 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=11.295
+ $Y=0.705 $X2=11.435 $Y2=0.92
r418 7 119 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=9.735
+ $Y=0.705 $X2=9.875 $Y2=0.92
r419 6 258 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=7.935
+ $Y=0.705 $X2=8.075 $Y2=0.92
r420 5 110 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=6.375
+ $Y=0.705 $X2=6.515 $Y2=0.94
r421 4 101 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=4.815
+ $Y=0.705 $X2=4.955 $Y2=0.92
r422 3 92 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.255
+ $Y=0.705 $X2=3.395 $Y2=0.94
r423 2 83 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.705 $X2=1.835 $Y2=0.94
r424 1 74 91 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.705 $X2=0.275 $Y2=0.94
.ends

