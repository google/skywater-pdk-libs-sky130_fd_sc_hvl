* File: sky130_fd_sc_hvl__mux2_1.pex.spice
* Created: Fri Aug 28 09:37:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__MUX2_1%VNB 5 7 11 25
r37 7 25 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=0.057
+ $X2=2.64 $Y2=0.058
r38 7 11 0.00134943 $w=5.28e-06 $l=5.7e-08 $layer=MET1_cond $X=2.64 $Y=0.057
+ $X2=2.64 $Y2=0
r39 5 11 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r40 5 11 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX2_1%VPB 4 6 14 21
r34 10 21 0.00134943 $w=5.28e-06 $l=5.7e-08 $layer=MET1_cond $X=2.64 $Y=4.07
+ $X2=2.64 $Y2=4.013
r35 10 14 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=4.07
+ $X2=5.04 $Y2=4.07
r36 9 14 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=5.04
+ $Y2=4.07
r37 9 10 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r38 6 21 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=4.012
+ $X2=2.64 $Y2=4.013
r39 4 14 33.0909 $w=1.7e-07 $l=5.08232e-06 $layer=licon1_NTAP_notbjt $count=5
+ $X=0 $Y=3.985 $X2=5.04 $Y2=4.07
r40 4 9 33.0909 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=5
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX2_1%A_94_81# 1 2 7 10 11 13 14 16 17 23 27 29 35
+ 39
c77 27 0 1.62611e-19 $X=2.715 $Y=0.745
c78 13 0 3.21722e-20 $X=2.55 $Y=2.5
c79 11 0 3.90172e-20 $X=2.385 $Y=1.44
r80 29 32 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=2.5
+ $X2=2.715 $Y2=2.665
r81 24 27 6.72258 $w=4.18e-07 $l=2.45e-07 $layer=LI1_cond $X=2.47 $Y=0.705
+ $X2=2.715 $Y2=0.705
r82 21 39 148.203 $w=5e-07 $l=1.385e-06 $layer=POLY_cond $X=0.72 $Y=1.58
+ $X2=0.72 $Y2=2.965
r83 21 35 71.6939 $w=5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.72 $Y=1.58 $X2=0.72
+ $Y2=0.91
r84 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.785
+ $Y=1.58 $X2=0.785 $Y2=1.58
r85 17 20 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.785 $Y=1.44
+ $X2=0.785 $Y2=1.58
r86 15 24 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.47 $Y=0.915
+ $X2=2.47 $Y2=0.705
r87 15 16 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.47 $Y=0.915
+ $X2=2.47 $Y2=1.355
r88 13 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=2.5
+ $X2=2.715 $Y2=2.5
r89 13 14 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.55 $Y=2.5
+ $X2=2.115 $Y2=2.5
r90 12 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=1.44
+ $X2=2.03 $Y2=1.44
r91 11 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.385 $Y=1.44
+ $X2=2.47 $Y2=1.355
r92 11 12 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.385 $Y=1.44
+ $X2=2.115 $Y2=1.44
r93 10 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.03 $Y=2.415
+ $X2=2.115 $Y2=2.5
r94 9 23 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=1.525 $X2=2.03
+ $Y2=1.44
r95 9 10 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.03 $Y=1.525
+ $X2=2.03 $Y2=2.415
r96 8 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=1.44
+ $X2=0.785 $Y2=1.44
r97 7 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.945 $Y=1.44 $X2=2.03
+ $Y2=1.44
r98 7 8 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=1.945 $Y=1.44
+ $X2=0.95 $Y2=1.44
r99 2 32 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=2.455 $X2=2.715 $Y2=2.665
r100 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.575
+ $Y=0.535 $X2=2.715 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX2_1%S 3 6 7 9 10 11 13 14 18 22 25 31
c73 25 0 1.06818e-19 $X=4.595 $Y=0.745
c74 9 0 1.93882e-19 $X=3.145 $Y=3.095
r75 28 31 93.6302 $w=5e-07 $l=8.75e-07 $layer=POLY_cond $X=4.595 $Y=1.79
+ $X2=4.595 $Y2=2.665
r76 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.53
+ $Y=1.79 $X2=4.53 $Y2=1.79
r77 25 28 111.821 $w=5e-07 $l=1.045e-06 $layer=POLY_cond $X=4.595 $Y=0.745
+ $X2=4.595 $Y2=1.79
r78 14 29 9.10802 $w=3.08e-07 $l=2.45e-07 $layer=LI1_cond $X=4.52 $Y=2.035
+ $X2=4.52 $Y2=1.79
r79 13 29 4.64695 $w=3.08e-07 $l=1.25e-07 $layer=LI1_cond $X=4.52 $Y=1.665
+ $X2=4.52 $Y2=1.79
r80 12 14 3.71756 $w=3.08e-07 $l=1e-07 $layer=LI1_cond $X=4.52 $Y=2.135 $X2=4.52
+ $Y2=2.035
r81 10 12 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=4.365 $Y=2.22
+ $X2=4.52 $Y2=2.135
r82 10 11 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=4.365 $Y=2.22
+ $X2=3.23 $Y2=2.22
r83 8 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.145 $Y=2.305
+ $X2=3.23 $Y2=2.22
r84 8 9 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.145 $Y=2.305
+ $X2=3.145 $Y2=3.095
r85 6 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.06 $Y=3.18
+ $X2=3.145 $Y2=3.095
r86 6 7 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=3.06 $Y=3.18
+ $X2=1.765 $Y2=3.18
r87 4 22 93.6302 $w=5e-07 $l=8.75e-07 $layer=POLY_cond $X=1.615 $Y=1.79
+ $X2=1.615 $Y2=2.665
r88 4 18 111.821 $w=5e-07 $l=1.045e-06 $layer=POLY_cond $X=1.615 $Y=1.79
+ $X2=1.615 $Y2=0.745
r89 3 4 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.6 $Y=1.79
+ $X2=1.6 $Y2=1.79
r90 1 7 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.6 $Y=3.095
+ $X2=1.765 $Y2=3.18
r91 1 3 45.5739 $w=3.28e-07 $l=1.305e-06 $layer=LI1_cond $X=1.6 $Y=3.095 $X2=1.6
+ $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX2_1%A0 3 5 7 8 10 11 12 16 24
c61 16 0 2.00504e-19 $X=3.105 $Y=0.745
c62 12 0 1.06818e-19 $X=3.6 $Y=1.295
c63 8 0 1.93882e-19 $X=2.46 $Y=2.13
c64 7 0 5.77401e-20 $X=2.46 $Y=2.13
r65 16 19 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.105 $Y=0.745
+ $X2=3.105 $Y2=1.23
r66 11 12 18.7516 $w=2.93e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.242
+ $X2=3.6 $Y2=1.242
r67 11 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.23 $X2=3.17 $Y2=1.23
r68 10 11 8.39916 $w=2.93e-07 $l=2.15e-07 $layer=LI1_cond $X=2.905 $Y=1.242
+ $X2=3.12 $Y2=1.242
r69 8 24 21.1255 $w=5.7e-07 $l=2.15e-07 $layer=POLY_cond $X=2.36 $Y=2.13
+ $X2=2.36 $Y2=2.345
r70 7 8 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.46 $Y=2.13
+ $X2=2.46 $Y2=2.13
r71 5 7 13.6822 $w=3.21e-07 $l=4.58912e-07 $layer=LI1_cond $X=2.82 $Y=1.785
+ $X2=2.46 $Y2=2.01
r72 4 10 7.47753 $w=2.95e-07 $l=1.85699e-07 $layer=LI1_cond $X=2.82 $Y=1.39
+ $X2=2.905 $Y2=1.242
r73 4 5 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.82 $Y=1.39 $X2=2.82
+ $Y2=1.785
r74 3 24 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.325 $Y=2.665 $X2=2.325
+ $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX2_1%A1 1 3 5 9 12 15
c54 12 0 3.21722e-20 $X=3.17 $Y=1.79
c55 5 0 8.21802e-20 $X=2.855 $Y=1.68
r56 12 15 93.6302 $w=5e-07 $l=8.75e-07 $layer=POLY_cond $X=3.105 $Y=1.79
+ $X2=3.105 $Y2=2.665
r57 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.79 $X2=3.17 $Y2=1.79
r58 9 13 12.8714 $w=3.83e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=1.762 $X2=3.17
+ $Y2=1.762
r59 8 12 3.74521 $w=5e-07 $l=3.5e-08 $layer=POLY_cond $X=3.105 $Y=1.755
+ $X2=3.105 $Y2=1.79
r60 6 7 32.9344 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.615 $Y=1.68
+ $X2=2.345 $Y2=1.68
r61 5 8 38.6381 $w=1.5e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.855 $Y=1.68
+ $X2=3.105 $Y2=1.755
r62 5 6 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.855 $Y=1.68
+ $X2=2.615 $Y2=1.68
r63 1 7 54.2318 $w=5.31e-07 $l=6.04917e-07 $layer=POLY_cond $X=2.325 $Y=1.085
+ $X2=2.345 $Y2=1.68
r64 1 3 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.325 $Y=1.085 $X2=2.325
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX2_1%A_713_81# 1 2 9 11 13 17 21 25 28 30
c46 28 0 2.43667e-19 $X=3.95 $Y=1.27
c47 11 0 5.77401e-20 $X=3.815 $Y=2.325
c48 9 0 1.62611e-19 $X=3.815 $Y=0.745
r49 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.95
+ $Y=1.27 $X2=3.95 $Y2=1.27
r50 23 30 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=1.275
+ $X2=5.025 $Y2=1.19
r51 23 25 64.0758 $w=2.48e-07 $l=1.39e-06 $layer=LI1_cond $X=5.025 $Y=1.275
+ $X2=5.025 $Y2=2.665
r52 19 30 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=1.105
+ $X2=5.025 $Y2=1.19
r53 19 21 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=5.025 $Y=1.105
+ $X2=5.025 $Y2=0.745
r54 18 28 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.115 $Y=1.19
+ $X2=3.99 $Y2=1.19
r55 17 30 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.9 $Y=1.19
+ $X2=5.025 $Y2=1.19
r56 17 18 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=4.9 $Y=1.19
+ $X2=4.115 $Y2=1.19
r57 11 29 92.6485 $w=5.52e-07 $l=1.07236e-06 $layer=POLY_cond $X=3.815 $Y=2.325
+ $X2=3.85 $Y2=1.27
r58 11 13 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.815 $Y=2.325
+ $X2=3.815 $Y2=2.665
r59 7 29 16.6811 $w=5.52e-07 $l=2.01742e-07 $layer=POLY_cond $X=3.815 $Y=1.085
+ $X2=3.85 $Y2=1.27
r60 7 9 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.815 $Y=1.085 $X2=3.815
+ $Y2=0.745
r61 2 25 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.845
+ $Y=2.455 $X2=4.985 $Y2=2.665
r62 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.535 $X2=4.985 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX2_1%X 1 2 7 8 9 10 11 12 13 24 48
r14 32 48 2.33603 $w=3.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.31 $Y=2.11
+ $X2=0.31 $Y2=2.035
r15 13 43 13.8605 $w=3.68e-07 $l=4.45e-07 $layer=LI1_cond $X=0.31 $Y=3.145
+ $X2=0.31 $Y2=3.59
r16 12 13 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.31 $Y=2.775
+ $X2=0.31 $Y2=3.145
r17 11 12 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.31 $Y=2.405
+ $X2=0.31 $Y2=2.775
r18 11 35 2.02456 $w=3.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.31 $Y=2.405
+ $X2=0.31 $Y2=2.34
r19 10 48 0.155736 $w=3.68e-07 $l=5e-09 $layer=LI1_cond $X=0.31 $Y=2.03 $X2=0.31
+ $Y2=2.035
r20 10 46 3.84076 $w=3.68e-07 $l=1.05e-07 $layer=LI1_cond $X=0.31 $Y=2.03
+ $X2=0.31 $Y2=1.925
r21 10 35 7.0081 $w=3.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.31 $Y=2.115
+ $X2=0.31 $Y2=2.34
r22 10 32 0.155736 $w=3.68e-07 $l=5e-09 $layer=LI1_cond $X=0.31 $Y=2.115
+ $X2=0.31 $Y2=2.11
r23 9 46 10.3322 $w=2.88e-07 $l=2.6e-07 $layer=LI1_cond $X=0.27 $Y=1.665
+ $X2=0.27 $Y2=1.925
r24 8 9 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.665
r25 7 8 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=0.925 $X2=0.27
+ $Y2=1.295
r26 7 24 10.5309 $w=2.88e-07 $l=2.65e-07 $layer=LI1_cond $X=0.27 $Y=0.925
+ $X2=0.27 $Y2=0.66
r27 2 43 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.185
+ $Y=2.215 $X2=0.33 $Y2=3.59
r28 2 35 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.185
+ $Y=2.215 $X2=0.33 $Y2=2.34
r29 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.185
+ $Y=0.535 $X2=0.33 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX2_1%VPWR 1 2 7 10 18 24
r32 22 24 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=3.525 $Y=3.63
+ $X2=4.605 $Y2=3.63
r33 21 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.605 $Y=3.59
+ $X2=4.605 $Y2=3.59
r34 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.525 $Y=3.59
+ $X2=3.525 $Y2=3.59
r35 18 21 8.6145 $w=1.308e-06 $l=9.25e-07 $layer=LI1_cond $X=4.065 $Y=2.665
+ $X2=4.065 $Y2=3.59
r36 13 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.145 $Y=3.59
+ $X2=1.145 $Y2=3.59
r37 10 13 25.7776 $w=5.78e-07 $l=1.25e-06 $layer=LI1_cond $X=0.965 $Y=2.34
+ $X2=0.965 $Y2=3.59
r38 7 22 0.339756 $w=3.7e-07 $l=8.85e-07 $layer=MET1_cond $X=2.64 $Y=3.63
+ $X2=3.525 $Y2=3.63
r39 7 15 0.573939 $w=3.7e-07 $l=1.495e-06 $layer=MET1_cond $X=2.64 $Y=3.63
+ $X2=1.145 $Y2=3.63
r40 2 18 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.065
+ $Y=2.455 $X2=4.205 $Y2=2.665
r41 1 13 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=0.97
+ $Y=2.215 $X2=1.11 $Y2=3.59
r42 1 10 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.97
+ $Y=2.215 $X2=1.11 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX2_1%VGND 1 2 7 10 25 26
r43 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.61 $Y=0.48
+ $X2=4.61 $Y2=0.48
r44 23 25 8.80749 $w=5.48e-07 $l=4.05e-07 $layer=LI1_cond $X=4.205 $Y=0.64
+ $X2=4.61 $Y2=0.64
r45 20 26 0.552824 $w=3.7e-07 $l=1.44e-06 $layer=MET1_cond $X=3.17 $Y=0.44
+ $X2=4.61 $Y2=0.44
r46 19 23 22.508 $w=5.48e-07 $l=1.035e-06 $layer=LI1_cond $X=3.17 $Y=0.64
+ $X2=4.205 $Y2=0.64
r47 19 20 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.17 $Y=0.48
+ $X2=3.17 $Y2=0.48
r48 11 14 0.552824 $w=3.7e-07 $l=1.44e-06 $layer=MET1_cond $X=0.68 $Y=0.44
+ $X2=2.12 $Y2=0.44
r49 10 16 1.36398 $w=1.608e-06 $l=1.8e-07 $layer=LI1_cond $X=1.4 $Y=0.48 $X2=1.4
+ $Y2=0.66
r50 10 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.12 $Y=0.48
+ $X2=2.12 $Y2=0.48
r51 10 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.68 $Y=0.48
+ $X2=0.68 $Y2=0.48
r52 7 20 0.20347 $w=3.7e-07 $l=5.3e-07 $layer=MET1_cond $X=2.64 $Y=0.44 $X2=3.17
+ $Y2=0.44
r53 7 14 0.199631 $w=3.7e-07 $l=5.2e-07 $layer=MET1_cond $X=2.64 $Y=0.44
+ $X2=2.12 $Y2=0.44
r54 2 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.065
+ $Y=0.535 $X2=4.205 $Y2=0.745
r55 1 16 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.97
+ $Y=0.535 $X2=1.11 $Y2=0.66
.ends

