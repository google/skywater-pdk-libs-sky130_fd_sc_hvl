* File: sky130_fd_sc_hvl__inv_16.spice
* Created: Wed Sep  2 09:06:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__inv_16.pex.spice"
.subckt sky130_fd_sc_hvl__inv_16  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1002_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000 SB=250012
+ A=0.375 P=2.5 MULT=1
MM1003 N_Y_M1002_d N_A_M1003_g N_VGND_M1003_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250001 SB=250011
+ A=0.375 P=2.5 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VGND_M1003_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250002 SB=250010
+ A=0.375 P=2.5 MULT=1
MM1006 N_Y_M1005_d N_A_M1006_g N_VGND_M1006_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250002 SB=250009
+ A=0.375 P=2.5 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_VGND_M1006_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250003 SB=250009
+ A=0.375 P=2.5 MULT=1
MM1012 N_Y_M1007_d N_A_M1012_g N_VGND_M1012_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250004 SB=250008
+ A=0.375 P=2.5 MULT=1
MM1013 N_Y_M1013_d N_A_M1013_g N_VGND_M1012_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250005 SB=250007
+ A=0.375 P=2.5 MULT=1
MM1016 N_Y_M1013_d N_A_M1016_g N_VGND_M1016_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250005 SB=250006
+ A=0.375 P=2.5 MULT=1
MM1018 N_Y_M1018_d N_A_M1018_g N_VGND_M1016_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250006 SB=250005
+ A=0.375 P=2.5 MULT=1
MM1020 N_Y_M1018_d N_A_M1020_g N_VGND_M1020_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250007 SB=250005
+ A=0.375 P=2.5 MULT=1
MM1021 N_Y_M1021_d N_A_M1021_g N_VGND_M1020_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250008 SB=250004
+ A=0.375 P=2.5 MULT=1
MM1023 N_Y_M1021_d N_A_M1023_g N_VGND_M1023_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250009 SB=250003
+ A=0.375 P=2.5 MULT=1
MM1025 N_Y_M1025_d N_A_M1025_g N_VGND_M1023_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250009 SB=250002
+ A=0.375 P=2.5 MULT=1
MM1028 N_Y_M1025_d N_A_M1028_g N_VGND_M1028_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250010 SB=250002
+ A=0.375 P=2.5 MULT=1
MM1030 N_Y_M1030_d N_A_M1030_g N_VGND_M1028_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250011 SB=250001
+ A=0.375 P=2.5 MULT=1
MM1031 N_Y_M1030_d N_A_M1031_g N_VGND_M1031_s N_VNB_M1002_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.2025 PD=1.03 PS=2.04 NRD=0 NRS=0 M=1 R=1.5 SA=250012 SB=250000
+ A=0.375 P=2.5 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250000 SB=250012
+ A=0.75 P=4 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1000_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001 SB=250011 A=0.75
+ P=4 MULT=1
MM1004 N_VPWR_M1001_d N_A_M1004_g N_Y_M1004_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002 SB=250010 A=0.75
+ P=4 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g N_Y_M1004_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002 SB=250009 A=0.75
+ P=4 MULT=1
MM1009 N_VPWR_M1008_d N_A_M1009_g N_Y_M1009_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250003 SB=250009 A=0.75
+ P=4 MULT=1
MM1010 N_VPWR_M1010_d N_A_M1010_g N_Y_M1009_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250004 SB=250008 A=0.75
+ P=4 MULT=1
MM1011 N_VPWR_M1010_d N_A_M1011_g N_Y_M1011_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250005 SB=250007 A=0.75
+ P=4 MULT=1
MM1014 N_VPWR_M1014_d N_A_M1014_g N_Y_M1011_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250005 SB=250006 A=0.75
+ P=4 MULT=1
MM1015 N_VPWR_M1014_d N_A_M1015_g N_Y_M1015_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250006 SB=250005 A=0.75
+ P=4 MULT=1
MM1017 N_VPWR_M1017_d N_A_M1017_g N_Y_M1015_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250007 SB=250005 A=0.75
+ P=4 MULT=1
MM1019 N_VPWR_M1017_d N_A_M1019_g N_Y_M1019_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250008 SB=250004 A=0.75
+ P=4 MULT=1
MM1022 N_VPWR_M1022_d N_A_M1022_g N_Y_M1019_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250009 SB=250003 A=0.75
+ P=4 MULT=1
MM1024 N_VPWR_M1022_d N_A_M1024_g N_Y_M1024_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250009 SB=250002 A=0.75
+ P=4 MULT=1
MM1026 N_VPWR_M1026_d N_A_M1026_g N_Y_M1024_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250010 SB=250002 A=0.75
+ P=4 MULT=1
MM1027 N_VPWR_M1026_d N_A_M1027_g N_Y_M1027_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250011 SB=250001 A=0.75
+ P=4 MULT=1
MM1029 N_VPWR_M1029_d N_A_M1029_g N_Y_M1027_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250012 SB=250000
+ A=0.75 P=4 MULT=1
DX32_noxref N_VNB_M1002_b N_VPB_M1000_b NWDIODE A=36.66 P=33.4
*
.include "sky130_fd_sc_hvl__inv_16.pxi.spice"
*
.ends
*
*
