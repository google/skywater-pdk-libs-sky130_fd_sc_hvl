* File: sky130_fd_sc_hvl__buf_4.spice
* Created: Wed Sep  2 09:04:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__buf_4.pex.spice"
.subckt sky130_fd_sc_hvl__buf_4  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_149_81#_M1000_g N_X_M1000_s N_VNB_M1000_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.105 PD=2.07 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250003 A=0.375 P=2.5 MULT=1
MM1002 N_VGND_M1002_d N_A_149_81#_M1002_g N_X_M1000_s N_VNB_M1000_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250001
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1003 N_VGND_M1002_d N_A_149_81#_M1003_g N_X_M1003_s N_VNB_M1000_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250002
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1005 N_VGND_M1005_d N_A_149_81#_M1005_g N_X_M1003_s N_VNB_M1000_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250002
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1007 N_A_149_81#_M1007_d N_A_M1007_g N_VGND_M1005_d N_VNB_M1000_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.105 PD=2.07 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250003
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_A_149_81#_M1004_g N_X_M1004_s N_VPB_M1004_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.21 PD=3.57 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250003 A=0.75 P=4 MULT=1
MM1006 N_VPWR_M1006_d N_A_149_81#_M1006_g N_X_M1004_s N_VPB_M1004_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001 SB=250002
+ A=0.75 P=4 MULT=1
MM1008 N_VPWR_M1006_d N_A_149_81#_M1008_g N_X_M1008_s N_VPB_M1004_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002 SB=250002
+ A=0.75 P=4 MULT=1
MM1009 N_VPWR_M1009_d N_A_149_81#_M1009_g N_X_M1008_s N_VPB_M1004_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002 SB=250001
+ A=0.75 P=4 MULT=1
MM1001 N_A_149_81#_M1001_d N_A_M1001_g N_VPWR_M1009_d N_VPB_M1004_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.21 PD=3.57 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250003
+ SB=250000 A=0.75 P=4 MULT=1
DX10_noxref N_VNB_M1000_b N_VPB_M1004_b NWDIODE A=14.196 P=16.12
*
.include "sky130_fd_sc_hvl__buf_4.pxi.spice"
*
.ends
*
*
