* File: sky130_fd_sc_hvl__mux4_1.pex.spice
* Created: Fri Aug 28 09:37:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__MUX4_1%VNB 5 7 11 25
c92 5 0 2.5389e-19 $X=-0.33 $Y=-0.265
r93 7 25 1.0016e-05 $w=1.248e-05 $l=1e-09 $layer=MET1_cond $X=6.24 $Y=0.057
+ $X2=6.24 $Y2=0.058
r94 7 11 0.000570913 $w=1.248e-05 $l=5.7e-08 $layer=MET1_cond $X=6.24 $Y=0.057
+ $X2=6.24 $Y2=0
r95 5 11 0.715385 $w=1.7e-07 $l=2.21e-06 $layer=mcon $count=13 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r96 5 11 0.715385 $w=1.7e-07 $l=2.21e-06 $layer=mcon $count=13 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%VPB 4 6 14 21
r124 10 21 0.000570913 $w=1.248e-05 $l=5.7e-08 $layer=MET1_cond $X=6.24 $Y=4.07
+ $X2=6.24 $Y2=4.013
r125 10 14 0.715385 $w=1.7e-07 $l=2.21e-06 $layer=mcon $count=13 $X=12.24
+ $Y=4.07 $X2=12.24 $Y2=4.07
r126 9 14 782.888 $w=1.68e-07 $l=1.2e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=12.24 $Y2=4.07
r127 9 10 0.715385 $w=1.7e-07 $l=2.21e-06 $layer=mcon $count=13 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r128 6 21 1.0016e-05 $w=1.248e-05 $l=1e-09 $layer=MET1_cond $X=6.24 $Y=4.012
+ $X2=6.24 $Y2=4.013
r129 4 14 14 $w=1.7e-07 $l=1.22824e-05 $layer=licon1_NTAP_notbjt $count=13 $X=0
+ $Y=3.985 $X2=12.24 $Y2=4.07
r130 4 9 14 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=13 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%S0 1 3 7 9 12 16 23 25 26 27 28 30 31 32 35
+ 37 39 46 48 49 50 55 59 65 67 68
c173 65 0 1.01701e-19 $X=5.31 $Y=1.265
c174 35 0 1.95782e-19 $X=2.87 $Y=1.53
c175 30 0 1.97986e-19 $X=2.77 $Y=2.8
c176 27 0 6.16607e-20 $X=2.89 $Y=3.72
c177 25 0 1.87716e-19 $X=2.03 $Y=2.5
c178 12 0 1.23038e-19 $X=6.015 $Y=3.345
r179 65 67 18.3095 $w=5.7e-07 $l=1.85e-07 $layer=POLY_cond $X=5.41 $Y=1.265
+ $X2=5.41 $Y2=1.08
r180 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.31
+ $Y=1.265 $X2=5.31 $Y2=1.265
r181 50 68 2.85366 $w=4.95e-07 $l=1.62e-07 $layer=LI1_cond $X=5.172 $Y=1.607
+ $X2=5.172 $Y2=1.445
r182 49 68 3.62448 $w=4.93e-07 $l=1.5e-07 $layer=LI1_cond $X=5.172 $Y=1.295
+ $X2=5.172 $Y2=1.445
r183 49 66 0.724896 $w=4.93e-07 $l=3e-08 $layer=LI1_cond $X=5.172 $Y=1.295
+ $X2=5.172 $Y2=1.265
r184 48 66 8.21549 $w=4.93e-07 $l=3.4e-07 $layer=LI1_cond $X=5.172 $Y=0.925
+ $X2=5.172 $Y2=1.265
r185 44 46 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.77 $Y=2.885
+ $X2=2.975 $Y2=2.885
r186 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.07
+ $Y=2.47 $X2=2.07 $Y2=2.47
r187 40 59 95.7703 $w=5e-07 $l=8.95e-07 $layer=POLY_cond $X=0.665 $Y=2.45
+ $X2=0.665 $Y2=3.345
r188 40 55 182.445 $w=5e-07 $l=1.705e-06 $layer=POLY_cond $X=0.665 $Y=2.45
+ $X2=0.665 $Y2=0.745
r189 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.73
+ $Y=2.45 $X2=0.73 $Y2=2.45
r190 36 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=2.97
+ $X2=2.975 $Y2=2.885
r191 36 37 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.975 $Y=2.97
+ $X2=2.975 $Y2=3.635
r192 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.53 $X2=2.87 $Y2=1.53
r193 32 34 0.531897 $w=3.23e-07 $l=1.5e-08 $layer=LI1_cond $X=2.855 $Y=1.607
+ $X2=2.87 $Y2=1.607
r194 31 50 4.35095 $w=3.25e-07 $l=2.47e-07 $layer=LI1_cond $X=4.925 $Y=1.607
+ $X2=5.172 $Y2=1.607
r195 31 34 72.8699 $w=3.23e-07 $l=2.055e-06 $layer=LI1_cond $X=4.925 $Y=1.607
+ $X2=2.87 $Y2=1.607
r196 30 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.77 $Y=2.8
+ $X2=2.77 $Y2=2.885
r197 29 32 7.72402 $w=3.25e-07 $l=2.01057e-07 $layer=LI1_cond $X=2.77 $Y=1.77
+ $X2=2.855 $Y2=1.607
r198 29 30 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.77 $Y=1.77
+ $X2=2.77 $Y2=2.8
r199 27 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.89 $Y=3.72
+ $X2=2.975 $Y2=3.635
r200 27 28 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.89 $Y=3.72
+ $X2=2.155 $Y2=3.72
r201 26 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.03 $Y=3.635
+ $X2=2.155 $Y2=3.72
r202 25 42 2.96623 $w=2.5e-07 $l=9.8e-08 $layer=LI1_cond $X=2.03 $Y=2.5 $X2=2.03
+ $Y2=2.402
r203 25 26 52.3209 $w=2.48e-07 $l=1.135e-06 $layer=LI1_cond $X=2.03 $Y=2.5
+ $X2=2.03 $Y2=3.635
r204 24 39 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.415
+ $X2=0.73 $Y2=2.415
r205 23 42 4.17693 $w=1.7e-07 $l=1.31339e-07 $layer=LI1_cond $X=1.905 $Y=2.415
+ $X2=2.03 $Y2=2.402
r206 23 24 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.905 $Y=2.415
+ $X2=0.895 $Y2=2.415
r207 18 35 49.6017 $w=4.8e-07 $l=4.45e-07 $layer=POLY_cond $X=2.945 $Y=1.085
+ $X2=2.945 $Y2=1.53
r208 16 18 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.935 $Y=0.745
+ $X2=2.935 $Y2=1.085
r209 10 20 6.82538 $w=5e-07 $l=4.25e-07 $layer=POLY_cond $X=6.015 $Y=2.795
+ $X2=6.015 $Y2=2.37
r210 10 12 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.015 $Y=2.795
+ $X2=6.015 $Y2=3.345
r211 9 20 49.2584 $w=5.92e-07 $l=7.89398e-07 $layer=POLY_cond $X=5.41 $Y=1.945
+ $X2=6.015 $Y2=2.37
r212 8 65 9.38648 $w=5.7e-07 $l=1e-07 $layer=POLY_cond $X=5.41 $Y=1.365 $X2=5.41
+ $Y2=1.265
r213 8 9 54.4416 $w=5.7e-07 $l=5.8e-07 $layer=POLY_cond $X=5.41 $Y=1.365
+ $X2=5.41 $Y2=1.945
r214 7 67 32.294 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.375 $Y=0.745
+ $X2=5.375 $Y2=1.08
r215 1 43 36.4082 $w=5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.155 $Y=2.83
+ $X2=2.155 $Y2=2.47
r216 1 3 55.108 $w=5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.155 $Y=2.83 $X2=2.155
+ $Y2=3.345
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%A2 2 5 9 11 12 13 17
c39 2 0 1.87716e-19 $X=1.43 $Y=2.74
r40 17 19 18.909 $w=5.3e-07 $l=1.85e-07 $layer=POLY_cond $X=1.43 $Y=1.665
+ $X2=1.43 $Y2=1.48
r41 12 13 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.3 $Y=1.665 $X2=1.3
+ $Y2=2.035
r42 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.35
+ $Y=1.665 $X2=1.35 $Y2=1.665
r43 9 11 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.445 $Y=3.345 $X2=1.445
+ $Y2=3.005
r44 5 19 78.6493 $w=5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.445 $Y=0.745
+ $X2=1.445 $Y2=1.48
r45 2 11 26.9849 $w=5.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.43 $Y=2.74
+ $X2=1.43 $Y2=3.005
r46 1 17 8.07592 $w=5.3e-07 $l=8e-08 $layer=POLY_cond $X=1.43 $Y=1.745 $X2=1.43
+ $Y2=1.665
r47 1 2 100.444 $w=5.3e-07 $l=9.95e-07 $layer=POLY_cond $X=1.43 $Y=1.745
+ $X2=1.43 $Y2=2.74
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%A_30_107# 1 2 9 13 18 22 26 31 35 36 38 42
+ 45 47 48 51 53 56 62 67
c142 67 0 1.10319e-19 $X=2.935 $Y=2.097
c143 51 0 1.48072e-19 $X=3.12 $Y=2.115
c144 38 0 1.53558e-19 $X=5.91 $Y=2.035
c145 35 0 1.23038e-19 $X=5.17 $Y=2.47
c146 22 0 4.77099e-20 $X=1.905 $Y=1.26
r147 54 67 60.25 $w=6.24e-07 $l=1.01546e-06 $layer=POLY_cond $X=2.155 $Y=1.555
+ $X2=2.935 $Y2=2.097
r148 52 67 14.2901 $w=6.24e-07 $l=1.85e-07 $layer=POLY_cond $X=3.12 $Y=2.097
+ $X2=2.935 $Y2=2.097
r149 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.12
+ $Y=2.115 $X2=3.12 $Y2=2.115
r150 47 48 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.275 $Y=3.345
+ $X2=0.275 $Y2=3.115
r151 43 62 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.155 $Y=1.23
+ $X2=6.155 $Y2=0.745
r152 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.075
+ $Y=1.23 $X2=6.075 $Y2=1.23
r153 40 42 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=6.075 $Y=1.95
+ $X2=6.075 $Y2=1.23
r154 39 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=2.035
+ $X2=5.17 $Y2=2.035
r155 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.91 $Y=2.035
+ $X2=6.075 $Y2=1.95
r156 38 39 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=5.91 $Y=2.035
+ $X2=5.335 $Y2=2.035
r157 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.17
+ $Y=2.47 $X2=5.17 $Y2=2.47
r158 33 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=2.12
+ $X2=5.17 $Y2=2.035
r159 33 35 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=5.17 $Y=2.12
+ $X2=5.17 $Y2=2.47
r160 32 51 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.285 $Y=2.035
+ $X2=3.16 $Y2=2.035
r161 31 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.005 $Y=2.035
+ $X2=5.17 $Y2=2.035
r162 31 32 112.214 $w=1.68e-07 $l=1.72e-06 $layer=LI1_cond $X=5.005 $Y=2.035
+ $X2=3.285 $Y2=2.035
r163 27 54 2.67515 $w=5e-07 $l=2.5e-08 $layer=POLY_cond $X=2.155 $Y=1.53
+ $X2=2.155 $Y2=1.555
r164 27 56 83.9996 $w=5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.155 $Y=1.53
+ $X2=2.155 $Y2=0.745
r165 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.07
+ $Y=1.53 $X2=2.07 $Y2=1.53
r166 24 26 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=2.03 $Y=1.345
+ $X2=2.03 $Y2=1.53
r167 23 45 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.44 $Y=1.26
+ $X2=0.275 $Y2=1.26
r168 22 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.905 $Y=1.26
+ $X2=2.03 $Y2=1.345
r169 22 23 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=1.905 $Y=1.26
+ $X2=0.44 $Y2=1.26
r170 20 45 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.195 $Y=1.345
+ $X2=0.275 $Y2=1.26
r171 20 48 115.476 $w=1.68e-07 $l=1.77e-06 $layer=LI1_cond $X=0.195 $Y=1.345
+ $X2=0.195 $Y2=3.115
r172 16 45 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.275 $Y=1.175
+ $X2=0.275 $Y2=1.26
r173 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.275 $Y=1.175
+ $X2=0.275 $Y2=0.745
r174 14 36 88.205 $w=3.5e-07 $l=5.35e-07 $layer=POLY_cond $X=5.16 $Y=3.005
+ $X2=5.16 $Y2=2.47
r175 13 14 41.2577 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.235 $Y=3.345
+ $X2=5.235 $Y2=3.005
r176 7 67 8.04834 $w=5e-07 $l=5.43e-07 $layer=POLY_cond $X=2.935 $Y=2.64
+ $X2=2.935 $Y2=2.097
r177 7 9 75.4392 $w=5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.935 $Y=2.64
+ $X2=2.935 $Y2=3.345
r178 2 47 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=3.135 $X2=0.275 $Y2=3.345
r179 1 18 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.535 $X2=0.275 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%A3 3 7 12 13 14 18 20
c48 18 0 1.97986e-19 $X=3.68 $Y=2.435
c49 12 0 5.704e-20 $X=3.71 $Y=1.585
c50 7 0 6.16607e-20 $X=3.745 $Y=3.345
c51 3 0 4.7602e-20 $X=3.645 $Y=0.745
r52 18 21 57.7743 $w=5.3e-07 $l=5.7e-07 $layer=POLY_cond $X=3.76 $Y=2.435
+ $X2=3.76 $Y2=3.005
r53 18 20 18.909 $w=5.3e-07 $l=1.85e-07 $layer=POLY_cond $X=3.76 $Y=2.435
+ $X2=3.76 $Y2=2.25
r54 13 14 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.665 $Y=2.405
+ $X2=3.665 $Y2=2.775
r55 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.68
+ $Y=2.435 $X2=3.68 $Y2=2.435
r56 12 20 71.1589 $w=5e-07 $l=6.65e-07 $layer=POLY_cond $X=3.775 $Y=1.585
+ $X2=3.775 $Y2=2.25
r57 11 12 42.4627 $w=6.3e-07 $l=5e-07 $layer=POLY_cond $X=3.71 $Y=1.085 $X2=3.71
+ $Y2=1.585
r58 7 21 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.745 $Y=3.345 $X2=3.745
+ $Y2=3.005
r59 3 11 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.645 $Y=0.745 $X2=3.645
+ $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%A1 3 7 8 9 10 15 18
r41 15 18 93.6302 $w=5e-07 $l=8.75e-07 $layer=POLY_cond $X=4.525 $Y=2.47
+ $X2=4.525 $Y2=3.345
r42 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.565 $Y=2.775
+ $X2=4.565 $Y2=3.145
r43 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.565 $Y=2.405
+ $X2=4.565 $Y2=2.775
r44 8 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.565
+ $Y=2.47 $X2=4.565 $Y2=2.47
r45 7 15 94.7002 $w=5e-07 $l=8.85e-07 $layer=POLY_cond $X=4.525 $Y=1.585
+ $X2=4.525 $Y2=2.47
r46 6 7 41.7992 $w=6.4e-07 $l=5e-07 $layer=POLY_cond $X=4.595 $Y=1.085 $X2=4.595
+ $Y2=1.585
r47 3 6 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.665 $Y=0.745 $X2=4.665
+ $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%A0 3 7 11 12 14 15 16 21
c44 12 0 1.23747e-19 $X=6.88 $Y=1.35
c45 11 0 1.53558e-19 $X=6.81 $Y=2.475
r46 15 16 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=6.935 $Y=1.95
+ $X2=6.935 $Y2=2.405
r47 15 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.935
+ $Y=1.95 $X2=6.935 $Y2=1.95
r48 14 15 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=6.935 $Y=1.665
+ $X2=6.935 $Y2=1.95
r49 12 21 60.5694 $w=5.3e-07 $l=6e-07 $layer=POLY_cond $X=6.88 $Y=1.35 $X2=6.88
+ $Y2=1.95
r50 12 13 26.9849 $w=5.3e-07 $l=2.65e-07 $layer=POLY_cond $X=6.88 $Y=1.35
+ $X2=6.88 $Y2=1.085
r51 10 21 2.52372 $w=5.3e-07 $l=2.5e-08 $layer=POLY_cond $X=6.88 $Y=1.975
+ $X2=6.88 $Y2=1.95
r52 10 11 50.7079 $w=5.3e-07 $l=5e-07 $layer=POLY_cond $X=6.81 $Y=1.975 $X2=6.81
+ $Y2=2.475
r53 7 13 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.865 $Y=0.745 $X2=6.865
+ $Y2=1.085
r54 3 11 93.0951 $w=5e-07 $l=8.7e-07 $layer=POLY_cond $X=6.725 $Y=3.345
+ $X2=6.725 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%S1 3 5 7 9 11 13 16 18 19 20 23 27 29 30 31
+ 32 37
c87 5 0 9.36113e-20 $X=9.435 $Y=1.295
r88 37 40 54.2411 $w=5.3e-07 $l=5.35e-07 $layer=POLY_cond $X=8.08 $Y=2.41
+ $X2=8.08 $Y2=2.945
r89 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.03
+ $Y=2.41 $X2=8.03 $Y2=2.41
r90 32 38 10.2596 $w=4.08e-07 $l=3.65e-07 $layer=LI1_cond $X=8.015 $Y=2.775
+ $X2=8.015 $Y2=2.41
r91 31 38 0.140542 $w=4.08e-07 $l=5e-09 $layer=LI1_cond $X=8.015 $Y=2.405
+ $X2=8.015 $Y2=2.41
r92 30 31 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=8.015 $Y=2.035
+ $X2=8.015 $Y2=2.405
r93 28 32 3.09192 $w=4.08e-07 $l=1.1e-07 $layer=LI1_cond $X=8.015 $Y=2.885
+ $X2=8.015 $Y2=2.775
r94 27 29 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=9.205 $Y=2.885
+ $X2=9.205 $Y2=1.985
r95 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.285
+ $Y=1.48 $X2=9.285 $Y2=1.48
r96 21 29 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=9.245 $Y=1.86
+ $X2=9.245 $Y2=1.985
r97 21 23 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=9.245 $Y=1.86
+ $X2=9.245 $Y2=1.48
r98 20 28 39.3849 $w=6.2e-08 $l=2.43824e-07 $layer=LI1_cond $X=8.22 $Y=2.97
+ $X2=8.015 $Y2=2.885
r99 19 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.12 $Y=2.97
+ $X2=9.205 $Y2=2.885
r100 19 20 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=9.12 $Y=2.97 $X2=8.22
+ $Y2=2.97
r101 14 18 20.4101 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=10.825 $Y=1.985
+ $X2=10.825 $Y2=1.735
r102 14 16 47.0826 $w=5e-07 $l=4.4e-07 $layer=POLY_cond $X=10.825 $Y=1.985
+ $X2=10.825 $Y2=2.425
r103 11 18 20.4101 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=10.825 $Y=1.485
+ $X2=10.825 $Y2=1.735
r104 11 13 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.825 $Y=1.485
+ $X2=10.825 $Y2=1.165
r105 10 24 13.111 $w=5e-07 $l=3.24731e-07 $layer=POLY_cond $X=9.685 $Y=1.735
+ $X2=9.4 $Y2=1.65
r106 9 18 5.30422 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=10.575 $Y=1.735
+ $X2=10.825 $Y2=1.735
r107 9 10 95.2352 $w=5e-07 $l=8.9e-07 $layer=POLY_cond $X=10.575 $Y=1.735
+ $X2=9.685 $Y2=1.735
r108 5 24 13.8197 $w=5e-07 $l=3.72089e-07 $layer=POLY_cond $X=9.435 $Y=1.295
+ $X2=9.4 $Y2=1.65
r109 5 7 54.573 $w=5e-07 $l=5.1e-07 $layer=POLY_cond $X=9.435 $Y=1.295 $X2=9.435
+ $Y2=0.785
r110 3 40 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=8.095 $Y=3.285
+ $X2=8.095 $Y2=2.945
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%A_1681_89# 1 2 8 11 14 18 21 25 27
c68 21 0 9.36113e-20 $X=10.435 $Y=1.165
r69 27 29 7.94589 $w=4.99e-07 $l=4.22788e-07 $layer=LI1_cond $X=10.21 $Y=2.425
+ $X2=9.985 $Y2=2.75
r70 25 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.985
+ $Y=2.75 $X2=9.985 $Y2=2.75
r71 24 27 0.366733 $w=4.99e-07 $l=1.5e-08 $layer=LI1_cond $X=10.21 $Y=2.41
+ $X2=10.21 $Y2=2.425
r72 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.985
+ $Y=2.41 $X2=9.985 $Y2=2.41
r73 19 24 10.2476 $w=4.99e-07 $l=3.76298e-07 $layer=LI1_cond $X=10.395 $Y=2.115
+ $X2=10.21 $Y2=2.41
r74 19 21 43.7928 $w=2.48e-07 $l=9.5e-07 $layer=LI1_cond $X=10.395 $Y=2.115
+ $X2=10.395 $Y2=1.165
r75 17 25 61.4149 $w=7.2e-07 $l=8.6e-07 $layer=POLY_cond $X=9.125 $Y=2.585
+ $X2=9.985 $Y2=2.585
r76 17 18 2.9237 $w=7.2e-07 $l=2.5e-07 $layer=POLY_cond $X=9.125 $Y=2.585
+ $X2=8.875 $Y2=2.585
r77 14 16 46.6574 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=8.655 $Y=0.785
+ $X2=8.655 $Y2=1.125
r78 9 18 32.8342 $w=3.9e-07 $l=3.6e-07 $layer=POLY_cond $X=8.875 $Y=2.945
+ $X2=8.875 $Y2=2.585
r79 9 11 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=8.875 $Y=2.945 $X2=8.875
+ $Y2=3.285
r80 8 18 32.8342 $w=3.9e-07 $l=4.11339e-07 $layer=POLY_cond $X=8.765 $Y=2.225
+ $X2=8.875 $Y2=2.585
r81 8 16 235.663 $w=2.8e-07 $l=1.1e-06 $layer=POLY_cond $X=8.765 $Y=2.225
+ $X2=8.765 $Y2=1.125
r82 2 27 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=10.31
+ $Y=2.215 $X2=10.435 $Y2=2.425
r83 1 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=10.29
+ $Y=0.955 $X2=10.435 $Y2=1.165
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%A_1669_615# 1 2 9 11 12 15 17 18 20 22 25 28
+ 30 34
c72 15 0 1.48312e-19 $X=9.045 $Y=0.7
r73 26 34 128.942 $w=5e-07 $l=1.205e-06 $layer=POLY_cond $X=11.815 $Y=1.76
+ $X2=11.815 $Y2=2.965
r74 26 30 81.3245 $w=5e-07 $l=7.6e-07 $layer=POLY_cond $X=11.815 $Y=1.76
+ $X2=11.815 $Y2=1
r75 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.75
+ $Y=1.76 $X2=11.75 $Y2=1.76
r76 23 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.87 $Y=1.76
+ $X2=10.785 $Y2=1.76
r77 23 25 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=10.87 $Y=1.76
+ $X2=11.75 $Y2=1.76
r78 21 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.785 $Y=1.925
+ $X2=10.785 $Y2=1.76
r79 21 22 111.561 $w=1.68e-07 $l=1.71e-06 $layer=LI1_cond $X=10.785 $Y=1.925
+ $X2=10.785 $Y2=3.635
r80 20 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.785 $Y=1.595
+ $X2=10.785 $Y2=1.76
r81 19 20 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=10.785 $Y=0.435
+ $X2=10.785 $Y2=1.595
r82 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.7 $Y=0.35
+ $X2=10.785 $Y2=0.435
r83 17 18 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=10.7 $Y=0.35
+ $X2=9.21 $Y2=0.35
r84 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.045 $Y=0.435
+ $X2=9.21 $Y2=0.35
r85 13 15 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=9.045 $Y=0.435
+ $X2=9.045 $Y2=0.7
r86 11 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.7 $Y=3.72
+ $X2=10.785 $Y2=3.635
r87 11 12 133.743 $w=1.68e-07 $l=2.05e-06 $layer=LI1_cond $X=10.7 $Y=3.72
+ $X2=8.65 $Y2=3.72
r88 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.485 $Y=3.635
+ $X2=8.65 $Y2=3.72
r89 7 9 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=8.485 $Y=3.635
+ $X2=8.485 $Y2=3.345
r90 2 9 600 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=8.345
+ $Y=3.075 $X2=8.485 $Y2=3.345
r91 1 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=8.905
+ $Y=0.575 $X2=9.045 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%VPWR 1 2 3 4 13 16 32 41 45 54
r95 51 54 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=11.135 $Y=3.63
+ $X2=11.855 $Y2=3.63
r96 50 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.855 $Y=3.59
+ $X2=11.855 $Y2=3.59
r97 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.135 $Y=3.59
+ $X2=11.135 $Y2=3.59
r98 48 50 11.4461 $w=8.88e-07 $l=8.35e-07 $layer=LI1_cond $X=11.495 $Y=2.755
+ $X2=11.495 $Y2=3.59
r99 45 48 5.68876 $w=8.88e-07 $l=4.15e-07 $layer=LI1_cond $X=11.495 $Y=2.34
+ $X2=11.495 $Y2=2.755
r100 42 51 1.5241 $w=3.7e-07 $l=3.97e-06 $layer=MET1_cond $X=7.165 $Y=3.63
+ $X2=11.135 $Y2=3.63
r101 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.165 $Y=3.59
+ $X2=7.165 $Y2=3.59
r102 39 41 0.980392 $w=6.08e-07 $l=5e-08 $layer=LI1_cond $X=7.115 $Y=3.4
+ $X2=7.165 $Y2=3.4
r103 36 42 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=6.445 $Y=3.63
+ $X2=7.165 $Y2=3.63
r104 35 39 13.1373 $w=6.08e-07 $l=6.7e-07 $layer=LI1_cond $X=6.445 $Y=3.4
+ $X2=7.115 $Y2=3.4
r105 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.445 $Y=3.59
+ $X2=6.445 $Y2=3.59
r106 29 32 0.588235 $w=6.08e-07 $l=3e-08 $layer=LI1_cond $X=4.105 $Y=3.4
+ $X2=4.135 $Y2=3.4
r107 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.105 $Y=3.59
+ $X2=4.105 $Y2=3.59
r108 26 30 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.385 $Y=3.63
+ $X2=4.105 $Y2=3.63
r109 25 29 14.1176 $w=6.08e-07 $l=7.2e-07 $layer=LI1_cond $X=3.385 $Y=3.4
+ $X2=4.105 $Y2=3.4
r110 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.385 $Y=3.59
+ $X2=3.385 $Y2=3.59
r111 22 26 0.740937 $w=3.7e-07 $l=1.93e-06 $layer=MET1_cond $X=1.455 $Y=3.63
+ $X2=3.385 $Y2=3.63
r112 20 22 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.735 $Y=3.63
+ $X2=1.455 $Y2=3.63
r113 19 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.455 $Y=3.59
+ $X2=1.455 $Y2=3.59
r114 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.735 $Y=3.59
+ $X2=0.735 $Y2=3.59
r115 16 19 3.14632 $w=9.48e-07 $l=2.45e-07 $layer=LI1_cond $X=1.095 $Y=3.345
+ $X2=1.095 $Y2=3.59
r116 13 36 0.0787006 $w=3.7e-07 $l=2.05e-07 $layer=MET1_cond $X=6.24 $Y=3.63
+ $X2=6.445 $Y2=3.63
r117 13 30 0.819638 $w=3.7e-07 $l=2.135e-06 $layer=MET1_cond $X=6.24 $Y=3.63
+ $X2=4.105 $Y2=3.63
r118 4 50 400 $w=1.7e-07 $l=1.49708e-06 $layer=licon1_PDIFF $count=1 $X=11.075
+ $Y=2.215 $X2=11.33 $Y2=3.59
r119 4 48 400 $w=1.7e-07 $l=6.5521e-07 $layer=licon1_PDIFF $count=1 $X=11.075
+ $Y=2.215 $X2=11.33 $Y2=2.755
r120 4 45 600 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=1 $X=11.075
+ $Y=2.215 $X2=11.33 $Y2=2.34
r121 3 39 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.975
+ $Y=3.135 $X2=7.115 $Y2=3.345
r122 2 32 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.995
+ $Y=3.135 $X2=4.135 $Y2=3.345
r123 1 16 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.915
+ $Y=3.135 $X2=1.055 $Y2=3.345
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%A_481_107# 1 2 3 4 15 18 19 22 23 24 26 27
+ 28 30 31 32 34 35 36 37 38 39 43 46
c155 34 0 1.05578e-19 $X=8.615 $Y=0.965
c156 24 0 4.7602e-20 $X=4.55 $Y=0.35
c157 22 0 5.704e-20 $X=4.465 $Y=1.095
c158 19 0 2.1202e-19 $X=4.38 $Y=1.18
r159 40 43 5.14483 $w=2.78e-07 $l=1.25e-07 $layer=LI1_cond $X=2.42 $Y=3.315
+ $X2=2.545 $Y2=3.315
r160 38 46 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=9.635 $Y=3.115
+ $X2=9.635 $Y2=3.285
r161 37 38 129.176 $w=1.68e-07 $l=1.98e-06 $layer=LI1_cond $X=9.635 $Y=1.135
+ $X2=9.635 $Y2=3.115
r162 35 37 6.58872 $w=3.88e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.55 $Y=1.05
+ $X2=9.635 $Y2=1.135
r163 35 49 8.33247 $w=3.88e-07 $l=3.58504e-07 $layer=LI1_cond $X=9.55 $Y=1.05
+ $X2=9.77 $Y2=0.785
r164 35 36 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=9.55 $Y=1.05
+ $X2=8.7 $Y2=1.05
r165 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.615 $Y=0.965
+ $X2=8.7 $Y2=1.05
r166 33 34 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.615 $Y=0.435
+ $X2=8.615 $Y2=0.965
r167 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.53 $Y=0.35
+ $X2=8.615 $Y2=0.435
r168 31 32 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.53 $Y=0.35 $X2=8
+ $Y2=0.35
r169 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.915 $Y=0.435
+ $X2=8 $Y2=0.35
r170 29 30 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=7.915 $Y=0.435
+ $X2=7.915 $Y2=1.175
r171 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.83 $Y=1.26
+ $X2=7.915 $Y2=1.175
r172 27 28 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=7.83 $Y=1.26
+ $X2=6.94 $Y2=1.26
r173 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.855 $Y=1.175
+ $X2=6.94 $Y2=1.26
r174 25 26 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.855 $Y=0.435
+ $X2=6.855 $Y2=1.175
r175 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.77 $Y=0.35
+ $X2=6.855 $Y2=0.435
r176 23 24 144.834 $w=1.68e-07 $l=2.22e-06 $layer=LI1_cond $X=6.77 $Y=0.35
+ $X2=4.55 $Y2=0.35
r177 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.465 $Y=0.435
+ $X2=4.55 $Y2=0.35
r178 21 22 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.465 $Y=0.435
+ $X2=4.465 $Y2=1.095
r179 20 39 3.08518 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=2.71 $Y=1.18
+ $X2=2.522 $Y2=1.18
r180 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.38 $Y=1.18
+ $X2=4.465 $Y2=1.095
r181 19 20 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=4.38 $Y=1.18
+ $X2=2.71 $Y2=1.18
r182 18 40 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.42 $Y=3.175
+ $X2=2.42 $Y2=3.315
r183 17 39 3.43356 $w=2.72e-07 $l=1.38109e-07 $layer=LI1_cond $X=2.42 $Y=1.265
+ $X2=2.522 $Y2=1.18
r184 17 18 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=2.42 $Y=1.265
+ $X2=2.42 $Y2=3.175
r185 13 39 3.43356 $w=2.72e-07 $l=8.5e-08 $layer=LI1_cond $X=2.522 $Y=1.095
+ $X2=2.522 $Y2=1.18
r186 13 15 10.7561 $w=3.73e-07 $l=3.5e-07 $layer=LI1_cond $X=2.522 $Y=1.095
+ $X2=2.522 $Y2=0.745
r187 4 46 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=9.125
+ $Y=3.075 $X2=9.635 $Y2=3.285
r188 3 43 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=3.135 $X2=2.545 $Y2=3.315
r189 2 49 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.685
+ $Y=0.575 $X2=9.825 $Y2=0.785
r190 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.405
+ $Y=0.535 $X2=2.545 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%A_1097_627# 1 2 3 4 13 15 17 23 24 26 27 30
+ 32 33 34 37 39 40 41 45
r109 42 45 4.39026 $w=4.18e-07 $l=1.6e-07 $layer=LI1_cond $X=7.545 $Y=3.325
+ $X2=7.705 $Y2=3.325
r110 35 37 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=8.265 $Y=1.57
+ $X2=8.265 $Y2=0.825
r111 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.18 $Y=1.655
+ $X2=8.265 $Y2=1.57
r112 33 34 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=8.18 $Y=1.655
+ $X2=7.63 $Y2=1.655
r113 32 42 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=7.545 $Y=3.115
+ $X2=7.545 $Y2=3.325
r114 31 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.545 $Y=2.915
+ $X2=7.545 $Y2=2.83
r115 31 32 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.545 $Y=2.915
+ $X2=7.545 $Y2=3.115
r116 30 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.545 $Y=2.745
+ $X2=7.545 $Y2=2.83
r117 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.545 $Y=1.74
+ $X2=7.63 $Y2=1.655
r118 29 30 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=7.545 $Y=1.74
+ $X2=7.545 $Y2=2.745
r119 28 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.59 $Y=2.83
+ $X2=6.505 $Y2=2.83
r120 27 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.46 $Y=2.83
+ $X2=7.545 $Y2=2.83
r121 27 28 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=7.46 $Y=2.83
+ $X2=6.59 $Y2=2.83
r122 26 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=2.745
+ $X2=6.505 $Y2=2.83
r123 25 26 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=6.505 $Y=0.915
+ $X2=6.505 $Y2=2.745
r124 23 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=2.83
+ $X2=6.505 $Y2=2.83
r125 23 24 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=6.42 $Y=2.83
+ $X2=5.79 $Y2=2.83
r126 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.705 $Y=2.915
+ $X2=5.79 $Y2=2.83
r127 21 39 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.705 $Y=2.915
+ $X2=5.705 $Y2=3.095
r128 17 25 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=6.42 $Y=0.765
+ $X2=6.505 $Y2=0.915
r129 17 19 25.1617 $w=2.98e-07 $l=6.55e-07 $layer=LI1_cond $X=6.42 $Y=0.765
+ $X2=5.765 $Y2=0.765
r130 13 39 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.625 $Y=3.26
+ $X2=5.625 $Y2=3.095
r131 13 15 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.625 $Y=3.26
+ $X2=5.625 $Y2=3.345
r132 4 45 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=7.56
+ $Y=3.075 $X2=7.705 $Y2=3.285
r133 3 15 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.485
+ $Y=3.135 $X2=5.625 $Y2=3.345
r134 2 37 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=8.12
+ $Y=0.575 $X2=8.265 $Y2=0.825
r135 1 19 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=5.625
+ $Y=0.535 $X2=5.765 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%X 1 2 7 8 9 10 11 12 13 22
r13 13 40 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=12.245 $Y=3.145
+ $X2=12.245 $Y2=3.57
r14 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=12.245 $Y=2.775
+ $X2=12.245 $Y2=3.145
r15 11 12 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=12.245 $Y=2.36
+ $X2=12.245 $Y2=2.775
r16 10 11 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=12.245 $Y=2.035
+ $X2=12.245 $Y2=2.36
r17 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=12.245 $Y=1.665
+ $X2=12.245 $Y2=2.035
r18 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=12.245 $Y=1.295
+ $X2=12.245 $Y2=1.665
r19 7 8 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=12.245 $Y=0.925
+ $X2=12.245 $Y2=1.295
r20 7 22 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=12.245 $Y=0.925
+ $X2=12.245 $Y2=0.77
r21 2 40 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=12.065
+ $Y=2.215 $X2=12.205 $Y2=3.57
r22 2 11 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=12.065
+ $Y=2.215 $X2=12.205 $Y2=2.36
r23 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.065
+ $Y=0.625 $X2=12.205 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HVL__MUX4_1%VGND 1 2 3 4 13 16 31 35 42 46
c81 46 0 1.23747e-19 $X=11.855 $Y=0.48
r82 48 50 6.85393 $w=8.88e-07 $l=5e-07 $layer=LI1_cond $X=11.495 $Y=0.75
+ $X2=11.495 $Y2=1.25
r83 43 46 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=11.135 $Y=0.44
+ $X2=11.855 $Y2=0.44
r84 42 48 3.70112 $w=8.88e-07 $l=2.7e-07 $layer=LI1_cond $X=11.495 $Y=0.48
+ $X2=11.495 $Y2=0.75
r85 42 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.855 $Y=0.48
+ $X2=11.855 $Y2=0.48
r86 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.135 $Y=0.48
+ $X2=11.135 $Y2=0.48
r87 36 43 1.37054 $w=3.7e-07 $l=3.57e-06 $layer=MET1_cond $X=7.565 $Y=0.44
+ $X2=11.135 $Y2=0.44
r88 35 39 5.98039 $w=5.28e-07 $l=2.65e-07 $layer=LI1_cond $X=7.385 $Y=0.48
+ $X2=7.385 $Y2=0.745
r89 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.565 $Y=0.48
+ $X2=7.565 $Y2=0.48
r90 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.085 $Y=0.48
+ $X2=4.085 $Y2=0.48
r91 29 31 1.08734 $w=5.48e-07 $l=5e-08 $layer=LI1_cond $X=4.035 $Y=0.64
+ $X2=4.085 $Y2=0.64
r92 26 32 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.365 $Y=0.44
+ $X2=4.085 $Y2=0.44
r93 25 29 14.5704 $w=5.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.365 $Y=0.64
+ $X2=4.035 $Y2=0.64
r94 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.365 $Y=0.48
+ $X2=3.365 $Y2=0.48
r95 20 26 0.733259 $w=3.7e-07 $l=1.91e-06 $layer=MET1_cond $X=1.455 $Y=0.44
+ $X2=3.365 $Y2=0.44
r96 17 20 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.735 $Y=0.44
+ $X2=1.455 $Y2=0.44
r97 16 22 3.40316 $w=9.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.095 $Y=0.48
+ $X2=1.095 $Y2=0.745
r98 16 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.455 $Y=0.48
+ $X2=1.455 $Y2=0.48
r99 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.735 $Y=0.48
+ $X2=0.735 $Y2=0.48
r100 13 36 0.508675 $w=3.7e-07 $l=1.325e-06 $layer=MET1_cond $X=6.24 $Y=0.44
+ $X2=7.565 $Y2=0.44
r101 13 32 0.827316 $w=3.7e-07 $l=2.155e-06 $layer=MET1_cond $X=6.24 $Y=0.44
+ $X2=4.085 $Y2=0.44
r102 4 50 182 $w=1.7e-07 $l=4.75132e-07 $layer=licon1_NDIFF $count=1 $X=11.075
+ $Y=0.955 $X2=11.425 $Y2=1.25
r103 4 48 182 $w=1.7e-07 $l=4.40738e-07 $layer=licon1_NDIFF $count=1 $X=11.075
+ $Y=0.955 $X2=11.425 $Y2=0.75
r104 3 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.115
+ $Y=0.535 $X2=7.255 $Y2=0.745
r105 2 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.895
+ $Y=0.535 $X2=4.035 $Y2=0.745
r106 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.915
+ $Y=0.535 $X2=1.055 $Y2=0.745
.ends

