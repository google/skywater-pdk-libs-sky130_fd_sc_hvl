* File: sky130_fd_sc_hvl__lsbufhv2hv_hl_1.pex.spice
* Created: Wed Sep  2 09:07:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%VNB 9 11 12 17 43
r24 12 29 0.00083912 $w=8.64e-06 $l=5.8e-08 $layer=MET1_cond $X=4.32 $Y=8.082
+ $X2=4.32 $Y2=8.14
r25 11 43 1.44676e-05 $w=8.64e-06 $l=1e-09 $layer=MET1_cond $X=4.32 $Y=0.057
+ $X2=4.32 $Y2=0.058
r26 11 17 0.000824653 $w=8.64e-06 $l=5.7e-08 $layer=MET1_cond $X=4.32 $Y=0.057
+ $X2=4.32 $Y2=0
r27 9 29 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=8.4 $Y=8.14
+ $X2=8.4 $Y2=8.14
r28 9 29 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=0.24 $Y=8.14
+ $X2=0.24 $Y2=8.14
r29 9 17 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r30 9 17 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%VPB 7 8 11 14 20 21
c21 21 0 2.74381e-19 $X=8.4 $Y=4.07
r22 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=4.07 $X2=8.4
+ $Y2=4.07
r23 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r24 11 21 2.61775 $w=2.3e-07 $l=4.08e-06 $layer=MET1_cond $X=4.32 $Y=4.07
+ $X2=8.4 $Y2=4.07
r25 11 15 2.61775 $w=2.3e-07 $l=4.08e-06 $layer=MET1_cond $X=4.32 $Y=4.07
+ $X2=0.24 $Y2=4.07
r26 8 20 91 $w=1.7e-07 $l=6.86185e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=7.755 $Y=3.985 $X2=8.4 $Y2=4.07
r27 7 14 182 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=1 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%LOWHVPWR 1 7 11 13 16 19
c33 1 0 1.29121e-19 $X=3.915 $Y=2.525
r34 22 25 14.2758 $w=6.18e-07 $l=7.4e-07 $layer=LI1_cond $X=3.875 $Y=3.16
+ $X2=3.875 $Y2=3.9
r35 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.075 $Y=3.16
+ $X2=4.075 $Y2=3.16
r36 19 22 9.83871 $w=6.18e-07 $l=5.1e-07 $layer=LI1_cond $X=3.875 $Y=2.65
+ $X2=3.875 $Y2=3.16
r37 16 23 0.122109 $w=2.85e-07 $l=2.45e-07 $layer=MET1_cond $X=4.32 $Y=3.162
+ $X2=4.075 $Y2=3.162
r38 13 25 7.04143 $w=6.18e-07 $l=3.65e-07 $layer=LI1_cond $X=3.875 $Y=4.265
+ $X2=3.875 $Y2=3.9
r39 13 15 3.33324 $w=6.2e-07 $l=3.78622e-07 $layer=LI1_cond $X=3.875 $Y=4.265
+ $X2=3.657 $Y2=4.55
r40 9 15 3.49891 $w=5.7e-07 $l=5.28e-07 $layer=LI1_cond $X=4.185 $Y=4.55
+ $X2=3.657 $Y2=4.55
r41 9 11 14.7936 $w=5.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.185 $Y=4.55
+ $X2=4.89 $Y2=4.55
r42 7 15 36.4 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=5
+ $X=3.13 $Y=4.295 $X2=3.335 $Y2=4.38
r43 7 11 36.4 $w=1.7e-07 $l=1.802e-06 $layer=licon1_NTAP_notbjt $count=5 $X=3.13
+ $Y=4.295 $X2=4.89 $Y2=4.38
r44 1 25 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=3.915
+ $Y=2.525 $X2=4.055 $Y2=3.9
r45 1 19 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=3.915
+ $Y=2.525 $X2=4.055 $Y2=2.65
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%A_662_81# 1 2 9 12 16 20 24 27 28
+ 29 31
c42 12 0 1.42604e-19 $X=3.665 $Y=3.275
r43 28 32 31.3954 $w=6.05e-07 $l=3.35e-07 $layer=POLY_cond $X=3.612 $Y=1.56
+ $X2=3.612 $Y2=1.895
r44 28 31 16.3616 $w=6.05e-07 $l=1.65e-07 $layer=POLY_cond $X=3.612 $Y=1.56
+ $X2=3.612 $Y2=1.395
r45 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.73
+ $Y=1.56 $X2=3.73 $Y2=1.56
r46 22 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=1.605
+ $X2=4.99 $Y2=1.52
r47 22 24 48.1721 $w=2.48e-07 $l=1.045e-06 $layer=LI1_cond $X=4.99 $Y=1.605
+ $X2=4.99 $Y2=2.65
r48 18 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=1.435
+ $X2=4.99 $Y2=1.52
r49 18 20 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=4.99 $Y=1.435
+ $X2=4.99 $Y2=0.745
r50 17 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=1.52
+ $X2=3.73 $Y2=1.52
r51 16 29 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.865 $Y=1.52
+ $X2=4.99 $Y2=1.52
r52 16 17 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=4.865 $Y=1.52
+ $X2=3.895 $Y2=1.52
r53 12 32 147.668 $w=5e-07 $l=1.38e-06 $layer=POLY_cond $X=3.665 $Y=3.275
+ $X2=3.665 $Y2=1.895
r54 9 31 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.56 $Y=0.91 $X2=3.56
+ $Y2=1.395
r55 2 24 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.81
+ $Y=2.525 $X2=4.95 $Y2=2.65
r56 1 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.81
+ $Y=0.535 $X2=4.95 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%A 1 2 3 8 12 14
c20 12 0 1.42604e-19 $X=4.52 $Y=1.86
r21 11 14 111.286 $w=5e-07 $l=1.04e-06 $layer=POLY_cond $X=4.56 $Y=1.86 $X2=4.56
+ $Y2=2.9
r22 11 12 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.52
+ $Y=1.86 $X2=4.52 $Y2=1.86
r23 8 11 119.312 $w=5e-07 $l=1.115e-06 $layer=POLY_cond $X=4.56 $Y=0.745
+ $X2=4.56 $Y2=1.86
r24 2 3 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=2.405 $X2=4.52
+ $Y2=2.775
r25 1 2 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=2.035 $X2=4.52
+ $Y2=2.405
r26 1 12 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=4.52 $Y=2.035
+ $X2=4.52 $Y2=1.86
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%X 1 2 7 8 9 10 11 12 13 22
c17 2 0 1.45261e-19 $X=3.13 $Y=2.525
r18 13 41 21.7524 $w=3.98e-07 $l=7.55e-07 $layer=LI1_cond $X=3.195 $Y=3.145
+ $X2=3.195 $Y2=3.9
r19 12 13 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.195 $Y=2.775
+ $X2=3.195 $Y2=3.145
r20 12 35 3.60138 $w=3.98e-07 $l=1.25e-07 $layer=LI1_cond $X=3.195 $Y=2.775
+ $X2=3.195 $Y2=2.65
r21 11 35 7.05871 $w=3.98e-07 $l=2.45e-07 $layer=LI1_cond $X=3.195 $Y=2.405
+ $X2=3.195 $Y2=2.65
r22 10 11 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.195 $Y=2.035
+ $X2=3.195 $Y2=2.405
r23 9 10 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.195 $Y=1.665
+ $X2=3.195 $Y2=2.035
r24 8 9 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.195 $Y=1.295
+ $X2=3.195 $Y2=1.665
r25 7 8 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.195 $Y=0.925
+ $X2=3.195 $Y2=1.295
r26 7 22 7.05871 $w=3.98e-07 $l=2.45e-07 $layer=LI1_cond $X=3.195 $Y=0.925
+ $X2=3.195 $Y2=0.68
r27 2 41 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.525 $X2=3.275 $Y2=3.9
r28 2 35 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.525 $X2=3.275 $Y2=2.65
r29 1 22 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=3.045
+ $Y=0.535 $X2=3.17 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_HL_1%VGND 1 4 5 9
r18 15 17 5.32947 $w=9.48e-07 $l=4.15e-07 $layer=LI1_cond $X=4.04 $Y=0.745
+ $X2=4.04 $Y2=1.16
r19 9 15 3.40316 $w=9.48e-07 $l=2.65e-07 $layer=LI1_cond $X=4.04 $Y=0.48
+ $X2=4.04 $Y2=0.745
r20 9 10 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.68 $Y=0.48
+ $X2=3.68 $Y2=0.48
r21 4 10 0.245699 $w=3.7e-07 $l=6.4e-07 $layer=MET1_cond $X=4.32 $Y=0.44
+ $X2=3.68 $Y2=0.44
r22 4 9 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.4 $Y=0.48 $X2=4.4
+ $Y2=0.48
r23 1 17 182 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_NDIFF $count=1 $X=3.81
+ $Y=0.535 $X2=3.95 $Y2=1.16
r24 1 15 182 $w=1.7e-07 $l=4.5299e-07 $layer=licon1_NDIFF $count=1 $X=3.81
+ $Y=0.535 $X2=4.17 $Y2=0.745
.ends

