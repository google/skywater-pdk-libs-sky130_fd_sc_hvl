* NGSPICE file created from sky130_fd_sc_hvl__a21o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_83_283# B1 VGND VNB nhv w=750000u l=500000u
+  ad=2.1e+11p pd=2.06e+06u as=8.5875e+11p ps=5.29e+06u
M1001 VGND a_83_283# X VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=2.1375e+11p ps=2.07e+06u
M1002 VPWR a_83_283# X VPB phv w=1.5e+06u l=500000u
+  ad=8.475e+11p pd=7.13e+06u as=3.975e+11p ps=3.53e+06u
M1003 VPWR A1 a_469_443# VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=8.175e+11p ps=7.09e+06u
M1004 a_469_443# B1 a_83_283# VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=4.275e+11p ps=3.57e+06u
M1005 a_469_443# A2 VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_631_107# A1 a_83_283# VNB nhv w=750000u l=500000u
+  ad=1.575e+11p pd=1.92e+06u as=0p ps=0u
M1007 VGND A2 a_631_107# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends

