* File: sky130_fd_sc_hvl__o22a_1.spice
* Created: Fri Aug 28 09:38:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__o22a_1.pex.spice"
.subckt sky130_fd_sc_hvl__o22a_1  VNB VPB A1 B1 B2 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* B2	B2
* B1	B1
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_87_81#_M1003_g N_X_M1003_s N_VNB_M1003_b NHV L=0.5
+ W=0.75 AD=0.125625 AS=0.21375 PD=1.085 PS=2.07 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250003 A=0.375 P=2.5 MULT=1
MM1007 N_A_354_107#_M1007_d N_A1_M1007_g N_VGND_M1003_d N_VNB_M1003_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.125625 PD=1.03 PS=1.085 NRD=0 NRS=8.3562 M=1 R=1.5
+ SA=250001 SB=250002 A=0.375 P=2.5 MULT=1
MM1002 N_A_87_81#_M1002_d N_B1_M1002_g N_A_354_107#_M1007_d N_VNB_M1003_b NHV
+ L=0.5 W=0.75 AD=0.121875 AS=0.105 PD=1.075 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250002 SB=250002 A=0.375 P=2.5 MULT=1
MM1004 N_A_354_107#_M1004_d N_B2_M1004_g N_A_87_81#_M1002_d N_VNB_M1003_b NHV
+ L=0.5 W=0.75 AD=0.105 AS=0.121875 PD=1.03 PS=1.075 NRD=0 NRS=6.8286 M=1 R=1.5
+ SA=250002 SB=250001 A=0.375 P=2.5 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_354_107#_M1004_d N_VNB_M1003_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.105 PD=2.07 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250003
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1008 N_VPWR_M1008_d N_A_87_81#_M1008_g N_X_M1008_s N_VPB_M1008_b PHV L=0.5
+ W=1.5 AD=0.9225 AS=0.4275 PD=2.73 PS=3.57 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250004 A=0.75 P=4 MULT=1
MM1009 A_533_443# N_B1_M1009_g N_VPWR_M1008_d N_VPB_M1008_b PHV L=0.5 W=1.5
+ AD=0.1575 AS=0.9225 PD=1.71 PS=2.73 NRD=6.3603 NRS=120.96 M=1 R=3 SA=250002
+ SB=250002 A=0.75 P=4 MULT=1
MM1000 N_A_87_81#_M1000_d N_B2_M1000_g A_533_443# N_VPB_M1008_b PHV L=0.5 W=1.5
+ AD=0.21 AS=0.1575 PD=1.78 PS=1.71 NRD=0 NRS=6.3603 M=1 R=3 SA=250002 SB=250002
+ A=0.75 P=4 MULT=1
MM1005 A_831_443# N_A2_M1005_g N_A_87_81#_M1000_d N_VPB_M1008_b PHV L=0.5 W=1.5
+ AD=0.1575 AS=0.21 PD=1.71 PS=1.78 NRD=6.3603 NRS=0 M=1 R=3 SA=250003 SB=250001
+ A=0.75 P=4 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g A_831_443# N_VPB_M1008_b PHV L=0.5 W=1.5
+ AD=0.3975 AS=0.1575 PD=3.53 PS=1.71 NRD=0 NRS=6.3603 M=1 R=3 SA=250004
+ SB=250000 A=0.75 P=4 MULT=1
DX10_noxref N_VNB_M1003_b N_VPB_M1008_b NWDIODE A=15.444 P=17.08
*
.include "sky130_fd_sc_hvl__o22a_1.pxi.spice"
*
.ends
*
*
