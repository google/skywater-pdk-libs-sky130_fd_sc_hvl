* File: sky130_fd_sc_hvl__sdlclkp_1.pex.spice
* Created: Wed Sep  2 09:10:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%VNB 5 7 17 24
c88 5 0 6.67964e-20 $X=-0.33 $Y=-0.265
r89 11 24 3.0797 $w=2.3e-07 $l=4.8e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=5.04
+ $Y2=0
r90 7 17 3.38767 $w=2.3e-07 $l=5.28e-06 $layer=MET1_cond $X=5.52 $Y=0 $X2=10.8
+ $Y2=0
r91 7 24 0.30797 $w=2.3e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r92 5 17 0.808696 $w=1.7e-07 $l=1.955e-06 $layer=mcon $count=11 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r93 5 11 0.808696 $w=1.7e-07 $l=1.955e-06 $layer=mcon $count=11 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%VPB 4 6 14 15 21
r97 14 15 0.808696 $w=1.7e-07 $l=1.955e-06 $layer=mcon $count=11 $X=10.8 $Y=4.07
+ $X2=10.8 $Y2=4.07
r98 10 21 3.0797 $w=2.3e-07 $l=4.8e-06 $layer=MET1_cond $X=0.24 $Y=4.07 $X2=5.04
+ $Y2=4.07
r99 9 14 688.941 $w=1.68e-07 $l=1.056e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=10.8 $Y2=4.07
r100 9 10 0.808696 $w=1.7e-07 $l=1.955e-06 $layer=mcon $count=11 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r101 6 15 3.38767 $w=2.3e-07 $l=5.28e-06 $layer=MET1_cond $X=5.52 $Y=4.07
+ $X2=10.8 $Y2=4.07
r102 6 21 0.30797 $w=2.3e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=4.07
+ $X2=5.04 $Y2=4.07
r103 4 14 15.8261 $w=1.7e-07 $l=1.08424e-05 $layer=licon1_NTAP_notbjt $count=11
+ $X=0 $Y=3.985 $X2=10.8 $Y2=4.07
r104 4 9 15.8261 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=11
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%SCE 1 2 6 12
r18 9 12 111.286 $w=5e-07 $l=1.04e-06 $layer=POLY_cond $X=0.845 $Y=1.62
+ $X2=0.845 $Y2=2.66
r19 6 9 65.8086 $w=5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.845 $Y=1.005
+ $X2=0.845 $Y2=1.62
r20 1 2 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.76 $Y=1.62 $X2=0.76
+ $Y2=2.035
r21 1 9 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.76 $Y=1.62
+ $X2=0.76 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%GATE 1 2 6 12
r22 9 12 111.286 $w=5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.625 $Y=1.62
+ $X2=1.625 $Y2=2.66
r23 6 9 65.8086 $w=5e-07 $l=6.15e-07 $layer=POLY_cond $X=1.625 $Y=1.005
+ $X2=1.625 $Y2=1.62
r24 1 2 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.64 $Y=1.62 $X2=1.64
+ $Y2=2.035
r25 1 9 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.64 $Y=1.62
+ $X2=1.64 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%A_423_71# 1 2 9 12 14 17 19 22 25 28 32
+ 37 38 40 41 43 44 45 47 51 55
c113 19 0 4.52609e-21 $X=3.6 $Y=0.45
c114 12 0 1.75473e-19 $X=5.845 $Y=2.495
r115 41 57 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.8 $Y=3.13
+ $X2=5.8 $Y2=2.965
r116 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.97
+ $Y=3.13 $X2=5.97 $Y2=3.13
r117 38 40 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=5.03 $Y=3.11
+ $X2=5.97 $Y2=3.11
r118 35 38 6.81649 $w=2.1e-07 $l=1.48492e-07 $layer=LI1_cond $X=4.925 $Y=3.005
+ $X2=5.03 $Y2=3.11
r119 35 37 30.368 $w=2.08e-07 $l=5.75e-07 $layer=LI1_cond $X=4.925 $Y=3.005
+ $X2=4.925 $Y2=2.43
r120 34 45 3.98977 $w=2.3e-07 $l=9.44722e-08 $layer=LI1_cond $X=4.925 $Y=1.295
+ $X2=4.905 $Y2=1.21
r121 34 37 59.9437 $w=2.08e-07 $l=1.135e-06 $layer=LI1_cond $X=4.925 $Y=1.295
+ $X2=4.925 $Y2=2.43
r122 30 45 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=1.125
+ $X2=4.905 $Y2=1.21
r123 30 32 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.905 $Y=1.125
+ $X2=4.905 $Y2=0.87
r124 29 44 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.93 $Y=1.21
+ $X2=3.765 $Y2=1.21
r125 28 45 2.45049 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.78 $Y=1.21
+ $X2=4.905 $Y2=1.21
r126 28 29 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=4.78 $Y=1.21
+ $X2=3.93 $Y2=1.21
r127 26 51 128.407 $w=5e-07 $l=1.2e-06 $layer=POLY_cond $X=3.735 $Y=1.46
+ $X2=3.735 $Y2=2.66
r128 26 47 63.1335 $w=5e-07 $l=5.9e-07 $layer=POLY_cond $X=3.735 $Y=1.46
+ $X2=3.735 $Y2=0.87
r129 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.765
+ $Y=1.46 $X2=3.765 $Y2=1.46
r130 23 44 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=1.295
+ $X2=3.765 $Y2=1.21
r131 23 25 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=1.295
+ $X2=3.765 $Y2=1.46
r132 22 44 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.685 $Y=1.125
+ $X2=3.765 $Y2=1.21
r133 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.685 $Y=0.535
+ $X2=3.685 $Y2=1.125
r134 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.6 $Y=0.45
+ $X2=3.685 $Y2=0.535
r135 19 43 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.6 $Y=0.45
+ $X2=2.825 $Y2=0.45
r136 17 55 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.45 $Y=0.52
+ $X2=2.45 $Y2=0.685
r137 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.62
+ $Y=0.52 $X2=2.62 $Y2=0.52
r138 14 43 7.98337 $w=3.03e-07 $l=1.52e-07 $layer=LI1_cond $X=2.673 $Y=0.517
+ $X2=2.825 $Y2=0.517
r139 14 16 2.00261 $w=3.03e-07 $l=5.3e-08 $layer=LI1_cond $X=2.673 $Y=0.517
+ $X2=2.62 $Y2=0.517
r140 12 57 50.2928 $w=5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.845 $Y=2.495
+ $X2=5.845 $Y2=2.965
r141 9 55 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.405 $Y=1.005
+ $X2=2.405 $Y2=0.685
r142 2 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.765
+ $Y=2.285 $X2=4.905 $Y2=2.43
r143 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.765
+ $Y=0.66 $X2=4.905 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%A_431_431# 1 2 9 13 15 18 21 25 26 29 30
+ 31 34 35 37 39 42 44 45 48
c121 45 0 2.11044e-19 $X=6.1 $Y=1.78
c122 37 0 1.1081e-19 $X=6.39 $Y=3.385
c123 13 0 2.1354e-20 $X=5.845 $Y=1.005
r124 46 48 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.18 $Y=2.51
+ $X2=6.39 $Y2=2.51
r125 45 54 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.93 $Y=1.78
+ $X2=5.93 $Y2=1.615
r126 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.1
+ $Y=1.78 $X2=6.1 $Y2=1.78
r127 39 41 10.2694 $w=2.48e-07 $l=2.1e-07 $layer=LI1_cond $X=3.305 $Y=0.87
+ $X2=3.305 $Y2=1.08
r128 36 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=2.595
+ $X2=6.39 $Y2=2.51
r129 36 37 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.39 $Y=2.595
+ $X2=6.39 $Y2=3.385
r130 35 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.18 $Y=2.425
+ $X2=6.18 $Y2=2.51
r131 34 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.18 $Y=1.945
+ $X2=6.18 $Y2=1.78
r132 34 35 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6.18 $Y=1.945
+ $X2=6.18 $Y2=2.425
r133 30 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.305 $Y=3.47
+ $X2=6.39 $Y2=3.385
r134 30 31 107.973 $w=1.68e-07 $l=1.655e-06 $layer=LI1_cond $X=6.305 $Y=3.47
+ $X2=4.65 $Y2=3.47
r135 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.565 $Y=3.385
+ $X2=4.65 $Y2=3.47
r136 28 29 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.565 $Y=2.315
+ $X2=4.565 $Y2=3.385
r137 27 42 2.06925 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.455 $Y=2.23
+ $X2=3.345 $Y2=2.23
r138 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.48 $Y=2.23
+ $X2=4.565 $Y2=2.315
r139 26 27 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=4.48 $Y=2.23
+ $X2=3.455 $Y2=2.23
r140 23 25 41.6451 $w=2.18e-07 $l=7.95e-07 $layer=LI1_cond $X=3.345 $Y=3.225
+ $X2=3.345 $Y2=2.43
r141 22 42 4.36305 $w=2.07e-07 $l=8.5e-08 $layer=LI1_cond $X=3.345 $Y=2.315
+ $X2=3.345 $Y2=2.23
r142 22 25 6.02413 $w=2.18e-07 $l=1.15e-07 $layer=LI1_cond $X=3.345 $Y=2.315
+ $X2=3.345 $Y2=2.43
r143 21 42 4.36305 $w=2.07e-07 $l=9.12688e-08 $layer=LI1_cond $X=3.332 $Y=2.145
+ $X2=3.345 $Y2=2.23
r144 21 41 60.5734 $w=1.93e-07 $l=1.065e-06 $layer=LI1_cond $X=3.332 $Y=2.145
+ $X2=3.332 $Y2=1.08
r145 18 51 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.49 $Y=3.36
+ $X2=2.49 $Y2=3.195
r146 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.66
+ $Y=3.36 $X2=2.66 $Y2=3.36
r147 15 23 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=3.235 $Y=3.335
+ $X2=3.345 $Y2=3.225
r148 15 17 30.1207 $w=2.18e-07 $l=5.75e-07 $layer=LI1_cond $X=3.235 $Y=3.335
+ $X2=2.66 $Y2=3.335
r149 13 54 65.2736 $w=5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.845 $Y=1.005
+ $X2=5.845 $Y2=1.615
r150 9 51 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.405 $Y=2.66
+ $X2=2.405 $Y2=3.195
r151 2 25 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=3.22
+ $Y=2.285 $X2=3.345 $Y2=2.43
r152 1 39 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.66 $X2=3.345 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%A_1261_133# 1 2 9 14 19 20 22 23 26 30 32
+ 34 37 44 48
c78 23 0 1.53715e-19 $X=6.805 $Y=1.98
c79 9 0 1.06584e-19 $X=6.555 $Y=1.005
r80 38 48 111.286 $w=5e-07 $l=1.04e-06 $layer=POLY_cond $X=8.665 $Y=1.55
+ $X2=8.665 $Y2=2.59
r81 38 44 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=8.665 $Y=1.55
+ $X2=8.665 $Y2=1.065
r82 37 40 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=8.58 $Y=1.55
+ $X2=8.58 $Y2=1.72
r83 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.58
+ $Y=1.55 $X2=8.58 $Y2=1.55
r84 34 35 11.0976 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.755 $Y=1.72
+ $X2=7.755 $Y2=1.98
r85 33 34 2.2115 $w=2.1e-07 $l=1.35e-07 $layer=LI1_cond $X=7.89 $Y=1.72
+ $X2=7.755 $Y2=1.72
r86 32 40 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=8.415 $Y=1.72
+ $X2=8.58 $Y2=1.72
r87 32 33 27.7273 $w=2.08e-07 $l=5.25e-07 $layer=LI1_cond $X=8.415 $Y=1.72
+ $X2=7.89 $Y2=1.72
r88 28 35 4.48172 $w=2.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.755 $Y=2.085
+ $X2=7.755 $Y2=1.98
r89 28 30 17.5001 $w=2.68e-07 $l=4.1e-07 $layer=LI1_cond $X=7.755 $Y=2.085
+ $X2=7.755 $Y2=2.495
r90 24 34 4.48172 $w=2.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.755 $Y=1.615
+ $X2=7.755 $Y2=1.72
r91 24 26 26.0367 $w=2.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.755 $Y=1.615
+ $X2=7.755 $Y2=1.005
r92 22 35 2.2115 $w=2.1e-07 $l=1.35e-07 $layer=LI1_cond $X=7.62 $Y=1.98
+ $X2=7.755 $Y2=1.98
r93 22 23 43.0433 $w=2.08e-07 $l=8.15e-07 $layer=LI1_cond $X=7.62 $Y=1.98
+ $X2=6.805 $Y2=1.98
r94 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.64
+ $Y=1.62 $X2=6.64 $Y2=1.62
r95 17 23 7.26367 $w=2.1e-07 $l=2.11069e-07 $layer=LI1_cond $X=6.64 $Y=1.875
+ $X2=6.805 $Y2=1.98
r96 17 19 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.64 $Y=1.875
+ $X2=6.64 $Y2=1.62
r97 15 20 93.5508 $w=3.3e-07 $l=5.35e-07 $layer=POLY_cond $X=6.64 $Y=2.155
+ $X2=6.64 $Y2=1.62
r98 14 15 42.5715 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.555 $Y=2.495
+ $X2=6.555 $Y2=2.155
r99 11 20 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=6.64 $Y=1.345
+ $X2=6.64 $Y2=1.62
r100 9 11 42.5715 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.555 $Y=1.005
+ $X2=6.555 $Y2=1.345
r101 2 30 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.585
+ $Y=2.285 $X2=7.725 $Y2=2.495
r102 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.585
+ $Y=0.795 $X2=7.725 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%A_495_311# 1 2 3 4 14 15 16 17 18 19 22
+ 26 31 34 41 48 50 52 53 56 64 69 71 74
c141 71 0 1.1081e-19 $X=7.335 $Y=1.005
c142 52 0 1.24125e-19 $X=5.455 $Y=2.495
c143 48 0 2.1354e-20 $X=5.477 $Y=0.395
c144 34 0 1.06584e-19 $X=7.085 $Y=1.28
r145 69 71 34.2419 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.335 $Y=0.685
+ $X2=7.335 $Y2=1.005
r146 65 69 52.6077 $w=3.39e-07 $l=3.7e-07 $layer=POLY_cond $X=7.705 $Y=0.495
+ $X2=7.335 $Y2=0.495
r147 64 65 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.705
+ $Y=0.52 $X2=7.705 $Y2=0.52
r148 61 64 12.4391 $w=3.13e-07 $l=3.4e-07 $layer=LI1_cond $X=7.365 $Y=0.512
+ $X2=7.705 $Y2=0.512
r149 59 74 107.541 $w=5e-07 $l=1.005e-06 $layer=POLY_cond $X=7.335 $Y=1.49
+ $X2=7.335 $Y2=2.495
r150 59 71 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.335 $Y=1.49
+ $X2=7.335 $Y2=1.005
r151 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.25
+ $Y=1.49 $X2=7.25 $Y2=1.49
r152 52 53 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=5.477 $Y=2.495
+ $X2=5.477 $Y2=2.33
r153 45 48 10.5778 $w=2.78e-07 $l=2.57e-07 $layer=LI1_cond $X=5.22 $Y=0.395
+ $X2=5.477 $Y2=0.395
r154 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.22
+ $Y=0.41 $X2=5.22 $Y2=0.41
r155 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.98
+ $Y=1.72 $X2=2.98 $Y2=1.72
r156 38 41 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.795 $Y=1.72
+ $X2=2.98 $Y2=1.72
r157 36 61 4.34843 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=7.365 $Y=0.67
+ $X2=7.365 $Y2=0.512
r158 36 56 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=7.365 $Y=0.67
+ $X2=7.365 $Y2=1.195
r159 35 50 2.40986 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.62 $Y=1.28
+ $X2=5.477 $Y2=1.28
r160 34 58 6.63049 $w=3.63e-07 $l=2.1e-07 $layer=LI1_cond $X=7.267 $Y=1.28
+ $X2=7.267 $Y2=1.49
r161 34 56 5.9984 $w=3.63e-07 $l=8.5e-08 $layer=LI1_cond $X=7.267 $Y=1.28
+ $X2=7.267 $Y2=1.195
r162 34 35 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=7.085 $Y=1.28
+ $X2=5.62 $Y2=1.28
r163 32 50 4.02809 $w=2.27e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.42 $Y=1.365
+ $X2=5.477 $Y2=1.28
r164 32 53 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=5.42 $Y=1.365
+ $X2=5.42 $Y2=2.33
r165 29 50 4.02809 $w=2.27e-07 $l=8.5e-08 $layer=LI1_cond $X=5.477 $Y=1.195
+ $X2=5.477 $Y2=1.28
r166 29 31 7.68295 $w=2.83e-07 $l=1.9e-07 $layer=LI1_cond $X=5.477 $Y=1.195
+ $X2=5.477 $Y2=1.005
r167 28 48 0.630043 $w=2.85e-07 $l=1.4e-07 $layer=LI1_cond $X=5.477 $Y=0.535
+ $X2=5.477 $Y2=0.395
r168 28 31 19.0052 $w=2.83e-07 $l=4.7e-07 $layer=LI1_cond $X=5.477 $Y=0.535
+ $X2=5.477 $Y2=1.005
r169 24 38 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=1.885
+ $X2=2.795 $Y2=1.72
r170 24 26 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=2.795 $Y=1.885
+ $X2=2.795 $Y2=2.43
r171 20 38 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=1.555
+ $X2=2.795 $Y2=1.72
r172 20 22 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=2.795 $Y=1.555
+ $X2=2.795 $Y2=1.005
r173 19 42 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.995 $Y=1.72
+ $X2=2.98 $Y2=1.72
r174 18 46 38.9663 $w=3.64e-07 $l=1.68953e-07 $layer=POLY_cond $X=5.385 $Y=0.38
+ $X2=5.22 $Y2=0.372
r175 17 69 50.756 $w=3.39e-07 $l=3.02076e-07 $layer=POLY_cond $X=7.085 $Y=0.38
+ $X2=7.335 $Y2=0.495
r176 17 18 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=7.085 $Y=0.38
+ $X2=5.385 $Y2=0.38
r177 15 46 38.9663 $w=3.64e-07 $l=2.19499e-07 $layer=POLY_cond $X=5.055 $Y=0.245
+ $X2=5.22 $Y2=0.372
r178 15 16 979.383 $w=1.5e-07 $l=1.91e-06 $layer=POLY_cond $X=5.055 $Y=0.245
+ $X2=3.145 $Y2=0.245
r179 14 19 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.07 $Y=1.555
+ $X2=2.995 $Y2=1.72
r180 13 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.07 $Y=0.32
+ $X2=3.145 $Y2=0.245
r181 13 14 633.266 $w=1.5e-07 $l=1.235e-06 $layer=POLY_cond $X=3.07 $Y=0.32
+ $X2=3.07 $Y2=1.555
r182 4 52 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=5.33
+ $Y=2.285 $X2=5.455 $Y2=2.495
r183 3 26 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.655
+ $Y=2.285 $X2=2.795 $Y2=2.43
r184 2 31 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.33
+ $Y=0.795 $X2=5.455 $Y2=1.005
r185 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.655
+ $Y=0.795 $X2=2.795 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%CLK 1 3 4 7 8 9 10 13 14 20 25 26 27 30
+ 34 37 44 48
c102 37 0 4.52609e-21 $X=4.515 $Y=0.87
c103 10 0 1.82094e-19 $X=9.195 $Y=3.38
c104 1 0 8.39567e-20 $X=4.515 $Y=2.21
r105 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.485
+ $Y=1.55 $X2=4.485 $Y2=1.55
r106 37 40 72.764 $w=5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.515 $Y=0.87
+ $X2=4.515 $Y2=1.55
r107 34 41 1.75894 $w=5.08e-07 $l=7.5e-08 $layer=LI1_cond $X=4.56 $Y=1.72
+ $X2=4.485 $Y2=1.72
r108 31 48 74.9041 $w=5e-07 $l=7e-07 $layer=POLY_cond $X=9.445 $Y=1.89 $X2=9.445
+ $Y2=2.59
r109 31 44 88.2799 $w=5e-07 $l=8.25e-07 $layer=POLY_cond $X=9.445 $Y=1.89
+ $X2=9.445 $Y2=1.065
r110 30 33 5.41921 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=9.475 $Y=1.89
+ $X2=9.475 $Y2=2.025
r111 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.475
+ $Y=1.89 $X2=9.475 $Y2=1.89
r112 27 33 50.7075 $w=2.48e-07 $l=1.1e-06 $layer=LI1_cond $X=9.435 $Y=3.125
+ $X2=9.435 $Y2=2.025
r113 25 27 6.36223 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=9.377 $Y=3.29
+ $X2=9.377 $Y2=3.125
r114 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.36
+ $Y=3.29 $X2=9.36 $Y2=3.29
r115 21 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.36 $Y=3.305
+ $X2=9.36 $Y2=3.29
r116 20 26 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=9.36 $Y=3.095
+ $X2=9.36 $Y2=3.29
r117 18 48 27.2865 $w=5e-07 $l=2.55e-07 $layer=POLY_cond $X=9.445 $Y=2.845
+ $X2=9.445 $Y2=2.59
r118 18 20 32.941 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=9.445 $Y=2.845
+ $X2=9.445 $Y2=3.095
r119 14 16 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=6.42 $Y=3.38 $X2=6.42
+ $Y2=3.58
r120 12 40 54.573 $w=5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.515 $Y=2.06
+ $X2=4.515 $Y2=1.55
r121 12 13 6.88608 $w=5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.515 $Y=2.06
+ $X2=4.515 $Y2=2.135
r122 11 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.495 $Y=3.38
+ $X2=6.42 $Y2=3.38
r123 10 21 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=9.195 $Y=3.38
+ $X2=9.36 $Y2=3.305
r124 10 11 1384.47 $w=1.5e-07 $l=2.7e-06 $layer=POLY_cond $X=9.195 $Y=3.38
+ $X2=6.495 $Y2=3.38
r125 8 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.345 $Y=3.58
+ $X2=6.42 $Y2=3.58
r126 8 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=6.345 $Y=3.58
+ $X2=5.255 $Y2=3.58
r127 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.18 $Y=3.505
+ $X2=5.255 $Y2=3.58
r128 6 7 664.032 $w=1.5e-07 $l=1.295e-06 $layer=POLY_cond $X=5.18 $Y=2.21
+ $X2=5.18 $Y2=3.505
r129 5 13 23.237 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.765 $Y=2.135
+ $X2=4.515 $Y2=2.135
r130 4 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.105 $Y=2.135
+ $X2=5.18 $Y2=2.21
r131 4 5 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.105 $Y=2.135
+ $X2=4.765 $Y2=2.135
r132 1 13 6.88608 $w=5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.515 $Y=2.21
+ $X2=4.515 $Y2=2.135
r133 1 3 43.38 $w=5e-07 $l=4.5e-07 $layer=POLY_cond $X=4.515 $Y=2.21 $X2=4.515
+ $Y2=2.66
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%A_1630_171# 1 2 9 12 14 19 22 26 28 29 30
+ 33
r59 29 34 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.24 $Y=1.56
+ $X2=10.24 $Y2=1.725
r60 29 33 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.24 $Y=1.56
+ $X2=10.24 $Y2=1.395
r61 28 30 19.9963 $w=3.38e-07 $l=5.05e-07 $layer=LI1_cond $X=10.41 $Y=1.555
+ $X2=9.905 $Y2=1.555
r62 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.41
+ $Y=1.56 $X2=10.41 $Y2=1.56
r63 25 26 2.36881 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=9.14 $Y=1.47
+ $X2=9.027 $Y2=1.47
r64 25 30 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=9.14 $Y=1.47
+ $X2=9.905 $Y2=1.47
r65 20 26 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=9.027 $Y=1.555
+ $X2=9.027 $Y2=1.47
r66 20 22 41.2318 $w=2.23e-07 $l=8.05e-07 $layer=LI1_cond $X=9.027 $Y=1.555
+ $X2=9.027 $Y2=2.36
r67 19 26 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=9.027 $Y=1.385
+ $X2=9.027 $Y2=1.47
r68 18 19 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=9.027 $Y=1.215
+ $X2=9.027 $Y2=1.385
r69 14 18 7.1387 $w=3.3e-07 $l=2.13787e-07 $layer=LI1_cond $X=8.915 $Y=1.05
+ $X2=9.027 $Y2=1.215
r70 14 16 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=8.915 $Y=1.05
+ $X2=8.275 $Y2=1.05
r71 12 34 132.687 $w=5e-07 $l=1.24e-06 $layer=POLY_cond $X=10.285 $Y=2.965
+ $X2=10.285 $Y2=1.725
r72 9 33 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=10.285 $Y=0.91
+ $X2=10.285 $Y2=1.395
r73 2 22 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.915
+ $Y=2.215 $X2=9.055 $Y2=2.36
r74 1 16 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=8.15
+ $Y=0.855 $X2=8.275 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%VPWR 1 2 3 4 5 16 18 22 24 26 28 32 36 41
+ 43 44 45 47 70 74 75 81 83 84 93
c116 83 0 1.82094e-19 $X=10.32 $Y=3.56
c117 75 0 8.39567e-20 $X=4.125 $Y=3.63
c118 26 0 1.75473e-19 $X=6.945 $Y=2.495
r119 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.56
+ $X2=10.32 $Y2=3.56
r120 80 83 13.2375 $w=3.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.895 $Y=3.63
+ $X2=10.32 $Y2=3.63
r121 80 81 7.556 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.895 $Y=3.63
+ $X2=9.73 $Y2=3.63
r122 78 79 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.76 $Y=3.56
+ $X2=6.76 $Y2=3.56
r123 73 93 0.353193 $w=3.7e-07 $l=9.2e-07 $layer=MET1_cond $X=4.12 $Y=3.63
+ $X2=5.04 $Y2=3.63
r124 72 75 0.155736 $w=3.68e-07 $l=5e-09 $layer=LI1_cond $X=4.12 $Y=3.63
+ $X2=4.125 $Y2=3.63
r125 72 74 17.8345 $w=3.68e-07 $l=4.95e-07 $layer=LI1_cond $X=4.12 $Y=3.63
+ $X2=3.625 $Y2=3.63
r126 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.12 $Y=3.56
+ $X2=4.12 $Y2=3.56
r127 68 70 4.9085 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=1.905 $Y=3.63
+ $X2=1.985 $Y2=3.63
r128 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.905 $Y=3.7
+ $X2=1.905 $Y2=3.7
r129 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.465 $Y=3.56
+ $X2=0.465 $Y2=3.56
r130 63 84 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=9.6 $Y=3.63
+ $X2=10.32 $Y2=3.63
r131 62 81 7.20909 $w=1.98e-07 $l=1.3e-07 $layer=LI1_cond $X=9.6 $Y=3.715
+ $X2=9.73 $Y2=3.715
r132 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.6 $Y=3.7 $X2=9.6
+ $Y2=3.7
r133 59 63 0.399262 $w=3.7e-07 $l=1.04e-06 $layer=MET1_cond $X=8.56 $Y=3.63
+ $X2=9.6 $Y2=3.63
r134 59 79 0.69103 $w=3.7e-07 $l=1.8e-06 $layer=MET1_cond $X=8.56 $Y=3.63
+ $X2=6.76 $Y2=3.63
r135 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.56 $Y=3.56
+ $X2=8.56 $Y2=3.56
r136 56 73 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.4 $Y=3.63
+ $X2=4.12 $Y2=3.63
r137 56 69 0.573939 $w=3.7e-07 $l=1.495e-06 $layer=MET1_cond $X=3.4 $Y=3.63
+ $X2=1.905 $Y2=3.63
r138 55 74 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=3.4 $Y=3.715
+ $X2=3.625 $Y2=3.715
r139 55 70 78.4682 $w=1.98e-07 $l=1.415e-06 $layer=LI1_cond $X=3.4 $Y=3.715
+ $X2=1.985 $Y2=3.715
r140 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.4 $Y=3.7
+ $X2=3.4 $Y2=3.7
r141 51 69 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=1.545 $Y=3.63
+ $X2=1.905 $Y2=3.63
r142 51 66 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=1.545 $Y=3.63
+ $X2=0.465 $Y2=3.63
r143 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.545 $Y=3.56
+ $X2=1.545 $Y2=3.56
r144 48 65 3.22716 $w=3.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=3.63
+ $X2=0.455 $Y2=3.63
r145 48 50 28.8111 $w=3.68e-07 $l=9.25e-07 $layer=LI1_cond $X=0.62 $Y=3.63
+ $X2=1.545 $Y2=3.63
r146 47 68 3.27045 $w=3.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.8 $Y=3.63
+ $X2=1.905 $Y2=3.63
r147 47 50 7.94251 $w=3.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.8 $Y=3.63
+ $X2=1.545 $Y2=3.63
r148 45 79 0.476043 $w=3.7e-07 $l=1.24e-06 $layer=MET1_cond $X=5.52 $Y=3.63
+ $X2=6.76 $Y2=3.63
r149 45 93 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.63
+ $X2=5.04 $Y2=3.63
r150 44 62 31.8864 $w=1.98e-07 $l=5.75e-07 $layer=LI1_cond $X=9.025 $Y=3.715
+ $X2=9.6 $Y2=3.715
r151 43 58 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.84 $Y=3.63
+ $X2=8.56 $Y2=3.63
r152 43 44 8.17894 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.84 $Y=3.63
+ $X2=9.025 $Y2=3.63
r153 40 58 3.73765 $w=3.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.44 $Y=3.63
+ $X2=8.56 $Y2=3.63
r154 40 41 4.69202 $w=3.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.44 $Y=3.63
+ $X2=8.275 $Y2=3.63
r155 36 39 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=9.895 $Y=2.36
+ $X2=9.895 $Y2=3.23
r156 34 80 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=9.895 $Y=3.445
+ $X2=9.895 $Y2=3.63
r157 34 39 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=9.895 $Y=3.445
+ $X2=9.895 $Y2=3.23
r158 30 41 1.75761 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=8.275 $Y=3.445
+ $X2=8.275 $Y2=3.63
r159 30 32 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=8.275 $Y=3.445
+ $X2=8.275 $Y2=2.36
r160 29 78 3.28189 $w=3.7e-07 $l=2.33e-07 $layer=LI1_cond $X=7.11 $Y=3.63
+ $X2=6.877 $Y2=3.63
r161 28 41 4.69202 $w=3.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.11 $Y=3.63
+ $X2=8.275 $Y2=3.63
r162 28 29 31.1471 $w=3.68e-07 $l=1e-06 $layer=LI1_cond $X=8.11 $Y=3.63 $X2=7.11
+ $Y2=3.63
r163 24 78 3.56359 $w=3.3e-07 $l=2.16345e-07 $layer=LI1_cond $X=6.945 $Y=3.445
+ $X2=6.877 $Y2=3.63
r164 24 26 33.1764 $w=3.28e-07 $l=9.5e-07 $layer=LI1_cond $X=6.945 $Y=3.445
+ $X2=6.945 $Y2=2.495
r165 20 75 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=4.125 $Y=3.445
+ $X2=4.125 $Y2=3.63
r166 20 22 30.5572 $w=3.28e-07 $l=8.75e-07 $layer=LI1_cond $X=4.125 $Y=3.445
+ $X2=4.125 $Y2=2.57
r167 16 65 3.61833 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=0.455 $Y=3.445
+ $X2=0.455 $Y2=3.63
r168 16 18 35.4464 $w=3.28e-07 $l=1.015e-06 $layer=LI1_cond $X=0.455 $Y=3.445
+ $X2=0.455 $Y2=2.43
r169 5 39 300 $w=1.7e-07 $l=1.11051e-06 $layer=licon1_PDIFF $count=2 $X=9.695
+ $Y=2.215 $X2=9.895 $Y2=3.23
r170 5 36 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=9.695
+ $Y=2.215 $X2=9.895 $Y2=2.36
r171 4 32 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=8.15
+ $Y=2.215 $X2=8.275 $Y2=2.36
r172 3 26 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.805
+ $Y=2.285 $X2=6.945 $Y2=2.495
r173 2 22 300 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=2 $X=3.985
+ $Y=2.285 $X2=4.125 $Y2=2.57
r174 1 18 300 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=2 $X=0.29
+ $Y=2.285 $X2=0.455 $Y2=2.43
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%A_58_159# 1 2 3 12 14 15 18 24 26 27
r37 26 27 7.32568 $w=2.93e-07 $l=1.35e-07 $layer=LI1_cond $X=1.997 $Y=2.43
+ $X2=1.997 $Y2=2.295
r38 22 24 3.95216 $w=2.32e-07 $l=1.12161e-07 $layer=LI1_cond $X=2.06 $Y=1.365
+ $X2=1.997 $Y2=1.28
r39 22 27 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.06 $Y=1.365
+ $X2=2.06 $Y2=2.295
r40 16 24 3.95216 $w=2.32e-07 $l=8.5e-08 $layer=LI1_cond $X=1.997 $Y=1.195
+ $X2=1.997 $Y2=1.28
r41 16 18 7.42251 $w=2.93e-07 $l=1.9e-07 $layer=LI1_cond $X=1.997 $Y=1.195
+ $X2=1.997 $Y2=1.005
r42 14 24 2.49072 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=1.85 $Y=1.28
+ $X2=1.997 $Y2=1.28
r43 14 15 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=1.85 $Y=1.28
+ $X2=0.62 $Y2=1.28
r44 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.455 $Y=1.195
+ $X2=0.62 $Y2=1.28
r45 10 12 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.455 $Y=1.195
+ $X2=0.455 $Y2=1.005
r46 3 26 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.875
+ $Y=2.285 $X2=2.015 $Y2=2.43
r47 2 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.875
+ $Y=0.795 $X2=2.015 $Y2=1.005
r48 1 12 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.29
+ $Y=0.795 $X2=0.455 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%GCLK 1 2 9 11 12 13 22 38
r21 29 31 38.2043 $w=3.63e-07 $l=1.21e-06 $layer=LI1_cond $X=10.772 $Y=2.36
+ $X2=10.772 $Y2=3.57
r22 26 38 1.3261 $w=3.63e-07 $l=4.2e-08 $layer=LI1_cond $X=10.772 $Y=2.077
+ $X2=10.772 $Y2=2.035
r23 22 34 3.41465 $w=2.68e-07 $l=8e-08 $layer=LI1_cond $X=10.82 $Y=1.295
+ $X2=10.82 $Y2=1.215
r24 13 38 0.694623 $w=3.63e-07 $l=2.2e-08 $layer=LI1_cond $X=10.772 $Y=2.013
+ $X2=10.772 $Y2=2.035
r25 13 36 4.52998 $w=3.63e-07 $l=1.18e-07 $layer=LI1_cond $X=10.772 $Y=2.013
+ $X2=10.772 $Y2=1.895
r26 13 29 8.27233 $w=3.63e-07 $l=2.62e-07 $layer=LI1_cond $X=10.772 $Y=2.098
+ $X2=10.772 $Y2=2.36
r27 13 26 0.663049 $w=3.63e-07 $l=2.1e-08 $layer=LI1_cond $X=10.772 $Y=2.098
+ $X2=10.772 $Y2=2.077
r28 12 36 9.81711 $w=2.68e-07 $l=2.3e-07 $layer=LI1_cond $X=10.82 $Y=1.665
+ $X2=10.82 $Y2=1.895
r29 11 34 0.898996 $w=3.63e-07 $l=3e-09 $layer=LI1_cond $X=10.772 $Y=1.212
+ $X2=10.772 $Y2=1.215
r30 11 12 15.7074 $w=2.68e-07 $l=3.68e-07 $layer=LI1_cond $X=10.82 $Y=1.297
+ $X2=10.82 $Y2=1.665
r31 11 22 0.0853661 $w=2.68e-07 $l=2e-09 $layer=LI1_cond $X=10.82 $Y=1.297
+ $X2=10.82 $Y2=1.295
r32 7 11 5.65171 $w=3.63e-07 $l=1.79e-07 $layer=LI1_cond $X=10.772 $Y=1.033
+ $X2=10.772 $Y2=1.212
r33 7 9 11.1455 $w=3.63e-07 $l=3.53e-07 $layer=LI1_cond $X=10.772 $Y=1.033
+ $X2=10.772 $Y2=0.68
r34 2 31 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=10.535
+ $Y=2.215 $X2=10.675 $Y2=3.57
r35 2 29 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=10.535
+ $Y=2.215 $X2=10.675 $Y2=2.36
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.535
+ $Y=0.535 $X2=10.675 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLCLKP_1%VGND 1 2 3 4 15 17 19 23 28 29 30 37 40
+ 45 53 63 64 72
r107 63 64 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=10.305 $Y=0.51
+ $X2=10.305 $Y2=0.51
r108 61 63 12.7703 $w=3.68e-07 $l=4.1e-07 $layer=LI1_cond $X=9.895 $Y=0.44
+ $X2=10.305 $Y2=0.44
r109 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.995 $Y=0.51
+ $X2=6.995 $Y2=0.51
r110 57 72 0.107494 $w=3.7e-07 $l=2.8e-07 $layer=MET1_cond $X=4.76 $Y=0.44
+ $X2=5.04 $Y2=0.44
r111 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.76 $Y=0.44
+ $X2=4.76 $Y2=0.44
r112 54 57 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=4.4 $Y=0.44
+ $X2=4.76 $Y2=0.44
r113 53 56 9.42489 $w=4.66e-07 $l=4.34741e-07 $layer=LI1_cond $X=4.4 $Y=0.605
+ $X2=4.76 $Y2=0.44
r114 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.4 $Y=0.51
+ $X2=4.4 $Y2=0.51
r115 51 53 7.19957 $w=4.66e-07 $l=2.75e-07 $layer=LI1_cond $X=4.125 $Y=0.605
+ $X2=4.4 $Y2=0.605
r116 48 64 0.829236 $w=3.7e-07 $l=2.16e-06 $layer=MET1_cond $X=8.145 $Y=0.44
+ $X2=10.305 $Y2=0.44
r117 48 60 0.441491 $w=3.7e-07 $l=1.15e-06 $layer=MET1_cond $X=8.145 $Y=0.44
+ $X2=6.995 $Y2=0.44
r118 47 48 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.145 $Y=0.44
+ $X2=8.145 $Y2=0.44
r119 45 61 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.73 $Y=0.44
+ $X2=9.895 $Y2=0.44
r120 45 47 49.3682 $w=3.68e-07 $l=1.585e-06 $layer=LI1_cond $X=9.73 $Y=0.44
+ $X2=8.145 $Y2=0.44
r121 43 60 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=5.915 $Y=0.44
+ $X2=6.995 $Y2=0.44
r122 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.915 $Y=0.44
+ $X2=5.915 $Y2=0.44
r123 40 59 3.22716 $w=3.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.78 $Y=0.44
+ $X2=6.945 $Y2=0.44
r124 40 42 26.9422 $w=3.68e-07 $l=8.65e-07 $layer=LI1_cond $X=6.78 $Y=0.44
+ $X2=5.915 $Y2=0.44
r125 38 54 1.07685 $w=3.7e-07 $l=2.805e-06 $layer=MET1_cond $X=1.595 $Y=0.44
+ $X2=4.4 $Y2=0.44
r126 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.595 $Y=0.51
+ $X2=1.595 $Y2=0.51
r127 34 38 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.875 $Y=0.44
+ $X2=1.595 $Y2=0.44
r128 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.875 $Y=0.51
+ $X2=0.875 $Y2=0.51
r129 30 43 0.151643 $w=3.7e-07 $l=3.95e-07 $layer=MET1_cond $X=5.52 $Y=0.44
+ $X2=5.915 $Y2=0.44
r130 30 72 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0.44
+ $X2=5.04 $Y2=0.44
r131 28 33 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=1.07 $Y=0.495
+ $X2=0.875 $Y2=0.495
r132 28 29 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=0.495
+ $X2=1.235 $Y2=0.495
r133 27 37 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=1.4 $Y=0.495
+ $X2=1.595 $Y2=0.495
r134 27 29 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=0.495
+ $X2=1.235 $Y2=0.495
r135 23 25 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=9.895 $Y=0.68
+ $X2=9.895 $Y2=1.09
r136 21 61 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=9.895 $Y=0.625
+ $X2=9.895 $Y2=0.44
r137 21 23 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=9.895 $Y=0.625
+ $X2=9.895 $Y2=0.68
r138 17 59 3.61833 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=6.945 $Y=0.625
+ $X2=6.945 $Y2=0.44
r139 17 19 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=6.945 $Y=0.625
+ $X2=6.945 $Y2=0.94
r140 13 29 0.499868 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=1.235 $Y=0.625
+ $X2=1.235 $Y2=0.495
r141 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.235 $Y=0.625
+ $X2=1.235 $Y2=0.92
r142 4 25 182 $w=1.7e-07 $l=3.19726e-07 $layer=licon1_NDIFF $count=1 $X=9.695
+ $Y=0.855 $X2=9.895 $Y2=1.09
r143 4 23 182 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_NDIFF $count=1 $X=9.695
+ $Y=0.855 $X2=9.895 $Y2=0.68
r144 3 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.805
+ $Y=0.795 $X2=6.945 $Y2=0.94
r145 2 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.985
+ $Y=0.66 $X2=4.125 $Y2=0.87
r146 1 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.795 $X2=1.235 $Y2=0.92
.ends

