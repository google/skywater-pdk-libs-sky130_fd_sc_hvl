# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__buf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.775000 2.775000 2.120000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.630000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.550000 1.390000 1.720000 ;
        RECT 0.125000 1.720000 1.370000 1.780000 ;
        RECT 1.200000 1.780000 1.370000 3.755000 ;
        RECT 1.220000 0.495000 1.390000 1.550000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.360000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.360000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.985000 3.360000 4.155000 ;
      RECT 0.090000  0.365000 1.040000 1.325000 ;
      RECT 0.090000  2.175000 1.020000 3.755000 ;
      RECT 1.550000  2.300000 2.800000 3.755000 ;
      RECT 1.570000  0.365000 2.820000 1.245000 ;
      RECT 1.570000  1.425000 3.250000 1.595000 ;
      RECT 1.570000  1.595000 1.865000 1.755000 ;
      RECT 2.980000  1.595000 3.250000 3.005000 ;
      RECT 3.000000  0.825000 3.250000 1.425000 ;
    LAYER mcon ;
      RECT 0.110000  3.505000 0.280000 3.675000 ;
      RECT 0.120000  0.395000 0.290000 0.565000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.470000  3.505000 0.640000 3.675000 ;
      RECT 0.480000  0.395000 0.650000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.830000  3.505000 1.000000 3.675000 ;
      RECT 0.840000  0.395000 1.010000 0.565000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.550000  3.505000 1.720000 3.675000 ;
      RECT 1.570000  0.395000 1.740000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.910000  3.505000 2.080000 3.675000 ;
      RECT 1.930000  0.395000 2.100000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.270000  3.505000 2.440000 3.675000 ;
      RECT 2.290000  0.395000 2.460000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.630000  3.505000 2.800000 3.675000 ;
      RECT 2.650000  0.395000 2.820000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
  END
END sky130_fd_sc_hvl__buf_2
END LIBRARY
