* File: sky130_fd_sc_hvl__buf_8.pex.spice
* Created: Fri Aug 28 09:33:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__BUF_8%VNB 5 7 11 25
r40 7 25 1.30208e-05 $w=9.6e-06 $l=1e-09 $layer=MET1_cond $X=4.8 $Y=0.057
+ $X2=4.8 $Y2=0.058
r41 7 11 0.000742187 $w=9.6e-06 $l=5.7e-08 $layer=MET1_cond $X=4.8 $Y=0.057
+ $X2=4.8 $Y2=0
r42 5 11 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r43 5 11 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_8%VPB 4 6 14 21
r82 10 21 0.000742187 $w=9.6e-06 $l=5.7e-08 $layer=MET1_cond $X=4.8 $Y=4.07
+ $X2=4.8 $Y2=4.013
r83 10 14 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=9.36 $Y=4.07
+ $X2=9.36 $Y2=4.07
r84 9 14 594.995 $w=1.68e-07 $l=9.12e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=9.36 $Y2=4.07
r85 9 10 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r86 6 21 1.30208e-05 $w=9.6e-06 $l=1e-09 $layer=MET1_cond $X=4.8 $Y=4.012
+ $X2=4.8 $Y2=4.013
r87 4 14 18.2 $w=1.7e-07 $l=9.4024e-06 $layer=licon1_NTAP_notbjt $count=10 $X=0
+ $Y=3.985 $X2=9.36 $Y2=4.07
r88 4 9 18.2 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=10 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_8%A 3 5 7 8 10 12 15 17 19 22 24 25 26 27 28 37
c71 15 0 1.75696e-19 $X=1.82 $Y=2.965
r72 36 37 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.82 $Y=1.815 $X2=2.6
+ $Y2=1.815
r73 34 36 9.0955 $w=5e-07 $l=8.5e-08 $layer=POLY_cond $X=1.735 $Y=1.815 $X2=1.82
+ $Y2=1.815
r74 27 28 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.697
+ $X2=2.16 $Y2=1.697
r75 27 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.735
+ $Y=1.73 $X2=1.735 $Y2=1.73
r76 26 27 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.697
+ $X2=1.68 $Y2=1.697
r77 25 26 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.697
+ $X2=1.2 $Y2=1.697
r78 20 37 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.6 $Y=2.065 $X2=2.6
+ $Y2=1.815
r79 20 22 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=2.6 $Y=2.065 $X2=2.6
+ $Y2=2.965
r80 17 37 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.6 $Y=1.565 $X2=2.6
+ $Y2=1.815
r81 17 19 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.6 $Y=1.565 $X2=2.6
+ $Y2=1.08
r82 13 36 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.82 $Y=2.065 $X2=1.82
+ $Y2=1.815
r83 13 15 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=1.82 $Y=2.065 $X2=1.82
+ $Y2=2.965
r84 10 36 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.82 $Y=1.565 $X2=1.82
+ $Y2=1.815
r85 10 12 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.82 $Y=1.565 $X2=1.82
+ $Y2=1.08
r86 9 24 5.30422 $w=5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.03 $Y=1.815 $X2=0.77
+ $Y2=1.815
r87 8 34 17.656 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.815 $X2=1.735
+ $Y2=1.815
r88 8 9 57.7832 $w=5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.57 $Y=1.815 $X2=1.03
+ $Y2=1.815
r89 5 24 20.4101 $w=5e-07 $l=2.54951e-07 $layer=POLY_cond $X=0.78 $Y=1.565
+ $X2=0.77 $Y2=1.815
r90 5 7 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.78 $Y=1.565 $X2=0.78
+ $Y2=1.08
r91 1 24 20.4101 $w=5e-07 $l=2.54951e-07 $layer=POLY_cond $X=0.76 $Y=2.065
+ $X2=0.77 $Y2=1.815
r92 1 3 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=0.76 $Y=2.065 $X2=0.76
+ $Y2=2.965
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_8%A_45_443# 1 2 3 4 15 17 19 22 24 26 29 31 33
+ 36 38 40 43 45 47 50 52 54 57 59 61 64 66 68 71 74 77 81 85 91 94 96 99 102
+ 103 104 107 109 119
c223 96 0 1.75696e-19 $X=2.51 $Y=2.095
c224 57 0 1.2129e-19 $X=8.06 $Y=1.08
r225 118 119 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=8.06 $Y=1.855
+ $X2=8.84 $Y2=1.855
r226 117 118 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.28 $Y=1.855
+ $X2=8.06 $Y2=1.855
r227 116 117 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=6.5 $Y=1.855
+ $X2=7.28 $Y2=1.855
r228 115 116 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=5.72 $Y=1.855
+ $X2=6.5 $Y2=1.855
r229 114 115 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=4.94 $Y=1.855
+ $X2=5.72 $Y2=1.855
r230 113 114 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=4.16 $Y=1.855
+ $X2=4.94 $Y2=1.855
r231 112 113 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.38 $Y=1.855
+ $X2=4.16 $Y2=1.855
r232 100 112 9.0955 $w=5e-07 $l=8.5e-08 $layer=POLY_cond $X=3.295 $Y=1.855
+ $X2=3.38 $Y2=1.855
r233 99 100 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.295
+ $Y=1.79 $X2=3.295 $Y2=1.79
r234 97 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.79
+ $X2=2.51 $Y2=1.79
r235 97 99 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.595 $Y=1.79
+ $X2=3.295 $Y2=1.79
r236 96 104 2.66603 $w=3.6e-07 $l=2.28583e-07 $layer=LI1_cond $X=2.51 $Y=2.095
+ $X2=2.32 $Y2=2.18
r237 95 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=1.955
+ $X2=2.51 $Y2=1.79
r238 95 96 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.51 $Y=1.955
+ $X2=2.51 $Y2=2.095
r239 94 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=1.625
+ $X2=2.51 $Y2=1.79
r240 93 107 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=1.4
+ $X2=2.51 $Y2=1.315
r241 93 94 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.51 $Y=1.4
+ $X2=2.51 $Y2=1.625
r242 89 107 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.21 $Y=1.315
+ $X2=2.51 $Y2=1.315
r243 89 91 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=2.21 $Y=1.23
+ $X2=2.21 $Y2=0.895
r244 85 87 22.1818 $w=5.48e-07 $l=1.02e-06 $layer=LI1_cond $X=2.32 $Y=2.34
+ $X2=2.32 $Y2=3.36
r245 83 104 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.32 $Y=2.265
+ $X2=2.32 $Y2=2.18
r246 83 85 1.63102 $w=5.48e-07 $l=7.5e-08 $layer=LI1_cond $X=2.32 $Y=2.265
+ $X2=2.32 $Y2=2.34
r247 82 103 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.435 $Y=2.18
+ $X2=0.34 $Y2=2.18
r248 81 104 4.14084 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.045 $Y=2.18
+ $X2=2.32 $Y2=2.18
r249 81 82 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=2.045 $Y=2.18
+ $X2=0.435 $Y2=2.18
r250 77 79 59.5407 $w=1.88e-07 $l=1.02e-06 $layer=LI1_cond $X=0.34 $Y=2.36
+ $X2=0.34 $Y2=3.38
r251 75 103 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.34 $Y=2.265
+ $X2=0.34 $Y2=2.18
r252 75 77 5.54545 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=0.34 $Y=2.265
+ $X2=0.34 $Y2=2.36
r253 74 103 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.34 $Y=2.095
+ $X2=0.34 $Y2=2.18
r254 74 102 36.1914 $w=1.88e-07 $l=6.2e-07 $layer=LI1_cond $X=0.34 $Y=2.095
+ $X2=0.34 $Y2=1.475
r255 69 102 5.66915 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=0.35 $Y=1.37
+ $X2=0.35 $Y2=1.475
r256 69 71 21.1255 $w=2.08e-07 $l=4e-07 $layer=LI1_cond $X=0.35 $Y=1.37 $X2=0.35
+ $Y2=0.97
r257 66 119 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.84 $Y=2.105
+ $X2=8.84 $Y2=1.855
r258 66 68 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.84 $Y=2.105 $X2=8.84
+ $Y2=2.965
r259 62 119 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.84 $Y=1.605
+ $X2=8.84 $Y2=1.855
r260 62 64 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=8.84 $Y=1.605
+ $X2=8.84 $Y2=1.08
r261 59 118 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.06 $Y=2.105
+ $X2=8.06 $Y2=1.855
r262 59 61 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.06 $Y=2.105 $X2=8.06
+ $Y2=2.965
r263 55 118 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.06 $Y=1.605
+ $X2=8.06 $Y2=1.855
r264 55 57 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=8.06 $Y=1.605
+ $X2=8.06 $Y2=1.08
r265 52 117 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.28 $Y=2.105
+ $X2=7.28 $Y2=1.855
r266 52 54 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.28 $Y=2.105 $X2=7.28
+ $Y2=2.965
r267 48 117 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.28 $Y=1.605
+ $X2=7.28 $Y2=1.855
r268 48 50 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=7.28 $Y=1.605
+ $X2=7.28 $Y2=1.08
r269 45 116 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.5 $Y=2.105 $X2=6.5
+ $Y2=1.855
r270 45 47 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.5 $Y=2.105 $X2=6.5
+ $Y2=2.965
r271 41 116 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.5 $Y=1.605 $X2=6.5
+ $Y2=1.855
r272 41 43 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=6.5 $Y=1.605 $X2=6.5
+ $Y2=1.08
r273 38 115 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.72 $Y=2.105
+ $X2=5.72 $Y2=1.855
r274 38 40 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.72 $Y=2.105 $X2=5.72
+ $Y2=2.965
r275 34 115 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.72 $Y=1.605
+ $X2=5.72 $Y2=1.855
r276 34 36 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=5.72 $Y=1.605
+ $X2=5.72 $Y2=1.08
r277 31 114 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.94 $Y=2.105
+ $X2=4.94 $Y2=1.855
r278 31 33 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.94 $Y=2.105 $X2=4.94
+ $Y2=2.965
r279 27 114 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.94 $Y=1.605
+ $X2=4.94 $Y2=1.855
r280 27 29 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.94 $Y=1.605
+ $X2=4.94 $Y2=1.08
r281 24 113 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.16 $Y=2.105
+ $X2=4.16 $Y2=1.855
r282 24 26 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.16 $Y=2.105 $X2=4.16
+ $Y2=2.965
r283 20 113 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.16 $Y=1.605
+ $X2=4.16 $Y2=1.855
r284 20 22 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.16 $Y=1.605
+ $X2=4.16 $Y2=1.08
r285 17 112 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.38 $Y=2.105
+ $X2=3.38 $Y2=1.855
r286 17 19 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.38 $Y=2.105 $X2=3.38
+ $Y2=2.965
r287 13 112 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.38 $Y=1.605
+ $X2=3.38 $Y2=1.855
r288 13 15 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.38 $Y=1.605
+ $X2=3.38 $Y2=1.08
r289 4 87 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=2.07
+ $Y=2.215 $X2=2.21 $Y2=3.36
r290 4 85 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.07
+ $Y=2.215 $X2=2.21 $Y2=2.34
r291 3 79 300 $w=1.7e-07 $l=1.22591e-06 $layer=licon1_PDIFF $count=2 $X=0.225
+ $Y=2.215 $X2=0.35 $Y2=3.38
r292 3 77 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.225
+ $Y=2.215 $X2=0.35 $Y2=2.36
r293 2 91 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=2.07
+ $Y=0.705 $X2=2.21 $Y2=0.895
r294 1 71 91 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=2 $X=0.245
+ $Y=0.705 $X2=0.37 $Y2=0.97
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_8%VPWR 1 2 3 4 5 6 19 21 23 25 29 31 36 38 40
+ 42 43 46 56 68 80 90 105 108
r123 104 105 14.2225 $w=3.18e-07 $l=3.25e-07 $layer=LI1_cond $X=9.23 $Y=3.635
+ $X2=8.905 $Y2=3.635
r124 100 101 1.3664 $w=1.248e-06 $l=1.4e-07 $layer=LI1_cond $X=1.24 $Y=3.57
+ $X2=1.24 $Y2=3.71
r125 96 98 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=1.42 $Y=3.63
+ $X2=1.78 $Y2=3.63
r126 94 96 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.7 $Y=3.63
+ $X2=1.42 $Y2=3.63
r127 93 100 0.0976 $w=1.248e-06 $l=1e-08 $layer=LI1_cond $X=1.24 $Y=3.56
+ $X2=1.24 $Y2=3.57
r128 93 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.78 $Y=3.56
+ $X2=1.78 $Y2=3.56
r129 93 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.42 $Y=3.56
+ $X2=1.42 $Y2=3.56
r130 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.7 $Y=3.56
+ $X2=0.7 $Y2=3.56
r131 90 93 9.8576 $w=1.248e-06 $l=1.01e-06 $layer=LI1_cond $X=1.24 $Y=2.55
+ $X2=1.24 $Y2=3.56
r132 86 108 0.506755 $w=3.7e-07 $l=1.32e-06 $layer=MET1_cond $X=8.03 $Y=3.63
+ $X2=9.35 $Y2=3.63
r133 84 86 0.274492 $w=3.7e-07 $l=7.15e-07 $layer=MET1_cond $X=7.315 $Y=3.63
+ $X2=8.03 $Y2=3.63
r134 83 88 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=7.67 $Y=3.56
+ $X2=7.67 $Y2=3.57
r135 83 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.03 $Y=3.56
+ $X2=8.03 $Y2=3.56
r136 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.315 $Y=3.56
+ $X2=7.315 $Y2=3.56
r137 80 83 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=7.67 $Y=2.55
+ $X2=7.67 $Y2=3.56
r138 76 84 0.3244 $w=3.7e-07 $l=8.45e-07 $layer=MET1_cond $X=6.47 $Y=3.63
+ $X2=7.315 $Y2=3.63
r139 74 76 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=6.11 $Y=3.63
+ $X2=6.47 $Y2=3.63
r140 72 74 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=5.75 $Y=3.63
+ $X2=6.11 $Y2=3.63
r141 71 78 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=6.11 $Y=3.56
+ $X2=6.11 $Y2=3.57
r142 71 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.47 $Y=3.56
+ $X2=6.47 $Y2=3.56
r143 71 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.11 $Y=3.56
+ $X2=6.11 $Y2=3.56
r144 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=3.56
+ $X2=5.75 $Y2=3.56
r145 68 71 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=6.11 $Y=2.55
+ $X2=6.11 $Y2=3.56
r146 64 72 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=4.91 $Y=3.63
+ $X2=5.75 $Y2=3.63
r147 60 62 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=4.19 $Y=3.63
+ $X2=4.55 $Y2=3.63
r148 59 66 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=4.55 $Y=3.56
+ $X2=4.55 $Y2=3.57
r149 59 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.91 $Y=3.56
+ $X2=4.91 $Y2=3.56
r150 59 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.55 $Y=3.56
+ $X2=4.55 $Y2=3.56
r151 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.19 $Y=3.56
+ $X2=4.19 $Y2=3.56
r152 56 59 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=4.55 $Y=2.55
+ $X2=4.55 $Y2=3.56
r153 52 60 0.374308 $w=3.7e-07 $l=9.75e-07 $layer=MET1_cond $X=3.215 $Y=3.63
+ $X2=4.19 $Y2=3.63
r154 50 52 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=2.855 $Y=3.63
+ $X2=3.215 $Y2=3.63
r155 50 98 0.412698 $w=3.7e-07 $l=1.075e-06 $layer=MET1_cond $X=2.855 $Y=3.63
+ $X2=1.78 $Y2=3.63
r156 49 54 0.178519 $w=6.68e-07 $l=1e-08 $layer=LI1_cond $X=3.1 $Y=3.56 $X2=3.1
+ $Y2=3.57
r157 49 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.215 $Y=3.56
+ $X2=3.215 $Y2=3.56
r158 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.855 $Y=3.56
+ $X2=2.855 $Y2=3.56
r159 46 49 18.0304 $w=6.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.1 $Y=2.55
+ $X2=3.1 $Y2=3.56
r160 43 64 0.0422296 $w=3.7e-07 $l=1.1e-07 $layer=MET1_cond $X=4.8 $Y=3.63
+ $X2=4.91 $Y2=3.63
r161 43 62 0.0959764 $w=3.7e-07 $l=2.5e-07 $layer=MET1_cond $X=4.8 $Y=3.63
+ $X2=4.55 $Y2=3.63
r162 41 88 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=7.67 $Y=3.625
+ $X2=7.67 $Y2=3.57
r163 41 42 3.33002 $w=8.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.67 $Y=3.625
+ $X2=7.67 $Y2=3.71
r164 39 78 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6.11 $Y=3.625
+ $X2=6.11 $Y2=3.57
r165 39 40 3.33002 $w=8.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.11 $Y=3.625
+ $X2=6.11 $Y2=3.71
r166 37 66 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=4.55 $Y=3.625
+ $X2=4.55 $Y2=3.57
r167 37 38 3.33002 $w=8.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=3.625
+ $X2=4.55 $Y2=3.71
r168 35 54 0.981855 $w=6.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.1 $Y=3.625
+ $X2=3.1 $Y2=3.57
r169 35 36 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=3.625 $X2=3.1
+ $Y2=3.71
r170 31 34 21.18 $w=3.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.32 $Y=2.55 $X2=9.32
+ $Y2=3.23
r171 29 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.35 $Y=3.56
+ $X2=9.35 $Y2=3.56
r172 29 104 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=9.32 $Y=3.635
+ $X2=9.23 $Y2=3.635
r173 29 34 7.63104 $w=3.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.32 $Y=3.475
+ $X2=9.32 $Y2=3.23
r174 28 42 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=8.115 $Y=3.71
+ $X2=7.67 $Y2=3.71
r175 28 105 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.115 $Y=3.71
+ $X2=8.905 $Y2=3.71
r176 26 40 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=6.555 $Y=3.71
+ $X2=6.11 $Y2=3.71
r177 25 42 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=7.225 $Y=3.71
+ $X2=7.67 $Y2=3.71
r178 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.225 $Y=3.71
+ $X2=6.555 $Y2=3.71
r179 24 38 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=4.995 $Y=3.71
+ $X2=4.55 $Y2=3.71
r180 23 40 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=5.665 $Y=3.71
+ $X2=6.11 $Y2=3.71
r181 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.665 $Y=3.71
+ $X2=4.995 $Y2=3.71
r182 22 36 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.435 $Y=3.71
+ $X2=3.1 $Y2=3.71
r183 21 38 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=4.105 $Y=3.71
+ $X2=4.55 $Y2=3.71
r184 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.105 $Y=3.71
+ $X2=3.435 $Y2=3.71
r185 20 101 13.277 $w=1.7e-07 $l=6.25e-07 $layer=LI1_cond $X=1.865 $Y=3.71
+ $X2=1.24 $Y2=3.71
r186 19 36 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.765 $Y=3.71
+ $X2=3.1 $Y2=3.71
r187 19 20 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.765 $Y=3.71
+ $X2=1.865 $Y2=3.71
r188 6 104 600 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=1 $X=9.09
+ $Y=2.215 $X2=9.23 $Y2=3.57
r189 6 34 400 $w=1.7e-07 $l=1.08274e-06 $layer=licon1_PDIFF $count=1 $X=9.09
+ $Y=2.215 $X2=9.23 $Y2=3.23
r190 6 31 400 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=9.09
+ $Y=2.215 $X2=9.23 $Y2=2.55
r191 5 88 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=7.53
+ $Y=2.215 $X2=7.67 $Y2=3.57
r192 5 80 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=7.53
+ $Y=2.215 $X2=7.67 $Y2=2.55
r193 4 78 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=5.97
+ $Y=2.215 $X2=6.11 $Y2=3.57
r194 4 68 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=5.97
+ $Y=2.215 $X2=6.11 $Y2=2.55
r195 3 66 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=4.41
+ $Y=2.215 $X2=4.55 $Y2=3.57
r196 3 56 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=4.41
+ $Y=2.215 $X2=4.55 $Y2=2.55
r197 2 54 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=2.85
+ $Y=2.215 $X2=2.99 $Y2=3.57
r198 2 46 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=2.85
+ $Y=2.215 $X2=2.99 $Y2=2.55
r199 1 100 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=2.215 $X2=1.15 $Y2=3.57
r200 1 90 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=2.215 $X2=1.15 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_8%X 1 2 3 4 5 6 7 8 27 33 35 36 37 38 41 47 49
+ 51 55 61 63 65 67 68 69 71 72 73 74 77 78 79 80 81 82 83 93 106
r100 103 106 2.37457 $w=6.78e-07 $l=1.35e-07 $layer=LI1_cond $X=8.625 $Y=2.205
+ $X2=8.625 $Y2=2.34
r101 83 118 4.44576 $w=5.9e-07 $l=2.15e-07 $layer=LI1_cond $X=8.625 $Y=3.145
+ $X2=8.625 $Y2=3.36
r102 83 104 4.82163 $w=6.8e-07 $l=2.55e-07 $layer=LI1_cond $X=8.625 $Y=3.145
+ $X2=8.625 $Y2=2.89
r103 82 104 2.02278 $w=6.78e-07 $l=1.15e-07 $layer=LI1_cond $X=8.625 $Y=2.775
+ $X2=8.625 $Y2=2.89
r104 81 82 6.50807 $w=6.78e-07 $l=3.7e-07 $layer=LI1_cond $X=8.625 $Y=2.405
+ $X2=8.625 $Y2=2.775
r105 81 106 1.14331 $w=6.78e-07 $l=6.5e-08 $layer=LI1_cond $X=8.625 $Y=2.405
+ $X2=8.625 $Y2=2.34
r106 80 103 2.14437 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=8.625 $Y=2.12
+ $X2=8.625 $Y2=2.205
r107 79 80 16.3847 $w=2.28e-07 $l=3.27e-07 $layer=LI1_cond $X=8.85 $Y=1.665
+ $X2=8.85 $Y2=1.992
r108 78 79 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.85 $Y=1.295
+ $X2=8.85 $Y2=1.665
r109 77 93 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=0.89 $X2=8.85
+ $Y2=0.975
r110 77 78 15.1822 $w=2.28e-07 $l=3.03e-07 $layer=LI1_cond $X=8.85 $Y=0.992
+ $X2=8.85 $Y2=1.295
r111 77 93 0.851806 $w=2.28e-07 $l=1.7e-08 $layer=LI1_cond $X=8.85 $Y=0.992
+ $X2=8.85 $Y2=0.975
r112 70 76 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.555 $Y=0.89
+ $X2=8.45 $Y2=0.89
r113 69 77 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.735 $Y=0.89
+ $X2=8.85 $Y2=0.89
r114 69 70 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.735 $Y=0.89
+ $X2=8.555 $Y2=0.89
r115 67 76 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=0.975
+ $X2=8.45 $Y2=0.89
r116 67 68 34.329 $w=2.08e-07 $l=6.5e-07 $layer=LI1_cond $X=8.45 $Y=0.975
+ $X2=8.45 $Y2=1.625
r117 66 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.055 $Y=2.12
+ $X2=6.89 $Y2=2.12
r118 65 80 5.03717 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=8.285 $Y=2.12
+ $X2=8.625 $Y2=2.12
r119 65 66 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=8.285 $Y=2.12
+ $X2=7.055 $Y2=2.12
r120 64 74 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.995 $Y=1.71
+ $X2=6.89 $Y2=1.71
r121 63 68 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.345 $Y=1.71
+ $X2=8.45 $Y2=1.625
r122 63 64 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=8.345 $Y=1.71
+ $X2=6.995 $Y2=1.71
r123 59 74 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.625
+ $X2=6.89 $Y2=1.71
r124 59 61 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=6.89 $Y=1.625
+ $X2=6.89 $Y2=0.97
r125 55 57 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=6.89 $Y=2.34
+ $X2=6.89 $Y2=3.36
r126 53 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=2.205
+ $X2=6.89 $Y2=2.12
r127 53 55 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.89 $Y=2.205
+ $X2=6.89 $Y2=2.34
r128 52 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.495 $Y=2.12
+ $X2=5.33 $Y2=2.12
r129 51 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=2.12
+ $X2=6.89 $Y2=2.12
r130 51 52 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=6.725 $Y=2.12
+ $X2=5.495 $Y2=2.12
r131 50 72 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.435 $Y=1.71
+ $X2=5.33 $Y2=1.71
r132 49 74 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.785 $Y=1.71
+ $X2=6.89 $Y2=1.71
r133 49 50 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=6.785 $Y=1.71
+ $X2=5.435 $Y2=1.71
r134 45 72 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.33 $Y=1.625
+ $X2=5.33 $Y2=1.71
r135 45 47 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=5.33 $Y=1.625
+ $X2=5.33 $Y2=0.97
r136 41 43 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=5.33 $Y=2.34
+ $X2=5.33 $Y2=3.36
r137 39 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.33 $Y=2.205
+ $X2=5.33 $Y2=2.12
r138 39 41 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.33 $Y=2.205
+ $X2=5.33 $Y2=2.34
r139 37 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=2.12
+ $X2=5.33 $Y2=2.12
r140 37 38 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=5.165 $Y=2.12
+ $X2=3.935 $Y2=2.12
r141 35 72 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.225 $Y=1.71
+ $X2=5.33 $Y2=1.71
r142 35 36 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=5.225 $Y=1.71
+ $X2=3.875 $Y2=1.71
r143 31 36 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.77 $Y=1.625
+ $X2=3.875 $Y2=1.71
r144 31 33 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=3.77 $Y=1.625
+ $X2=3.77 $Y2=0.97
r145 27 29 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3.77 $Y=2.34
+ $X2=3.77 $Y2=3.36
r146 25 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.77 $Y=2.205
+ $X2=3.935 $Y2=2.12
r147 25 27 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.77 $Y=2.205
+ $X2=3.77 $Y2=2.34
r148 8 118 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=8.31
+ $Y=2.215 $X2=8.45 $Y2=3.36
r149 8 106 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=8.31
+ $Y=2.215 $X2=8.45 $Y2=2.34
r150 7 57 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=6.75
+ $Y=2.215 $X2=6.89 $Y2=3.36
r151 7 55 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=6.75
+ $Y=2.215 $X2=6.89 $Y2=2.34
r152 6 43 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=5.19
+ $Y=2.215 $X2=5.33 $Y2=3.36
r153 6 41 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=5.19
+ $Y=2.215 $X2=5.33 $Y2=2.34
r154 5 29 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=3.63
+ $Y=2.215 $X2=3.77 $Y2=3.36
r155 5 27 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=3.63
+ $Y=2.215 $X2=3.77 $Y2=2.34
r156 4 76 91 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=2 $X=8.31
+ $Y=0.705 $X2=8.45 $Y2=0.97
r157 3 61 91 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=2 $X=6.75
+ $Y=0.705 $X2=6.89 $Y2=0.97
r158 2 47 91 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=2 $X=5.19
+ $Y=0.705 $X2=5.33 $Y2=0.97
r159 1 33 91 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=2 $X=3.63
+ $Y=0.705 $X2=3.77 $Y2=0.97
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_8%VGND 1 2 3 4 5 6 19 31 33 44 46 55 61 65 71
+ 75 81 83 85 86
c87 85 0 1.2129e-19 $X=9.42 $Y=0.465
r88 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.42 $Y=0.465
+ $X2=9.42 $Y2=0.465
r89 81 83 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=8.175 $Y=0.465
+ $X2=8.975 $Y2=0.465
r90 80 86 0.529789 $w=3.7e-07 $l=1.38e-06 $layer=MET1_cond $X=8.04 $Y=0.44
+ $X2=9.42 $Y2=0.44
r91 79 81 12.8638 $w=1.063e-06 $l=1.35e-07 $layer=LI1_cond $X=8.04 $Y=0.912
+ $X2=8.175 $Y2=0.912
r92 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.04 $Y=0.465
+ $X2=8.04 $Y2=0.465
r93 77 79 4.2385 $w=1.063e-06 $l=3.7e-07 $layer=LI1_cond $X=7.67 $Y=0.912
+ $X2=8.04 $Y2=0.912
r94 74 80 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.32 $Y=0.44
+ $X2=8.04 $Y2=0.44
r95 73 77 4.00939 $w=1.063e-06 $l=3.5e-07 $layer=LI1_cond $X=7.32 $Y=0.912
+ $X2=7.67 $Y2=0.912
r96 73 75 13.0929 $w=1.063e-06 $l=1.55e-07 $layer=LI1_cond $X=7.32 $Y=0.912
+ $X2=7.165 $Y2=0.912
r97 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.32 $Y=0.465
+ $X2=7.32 $Y2=0.465
r98 71 75 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.615 $Y=0.465
+ $X2=7.165 $Y2=0.465
r99 70 74 0.3244 $w=3.7e-07 $l=8.45e-07 $layer=MET1_cond $X=6.475 $Y=0.44
+ $X2=7.32 $Y2=0.44
r100 69 71 12.9211 $w=1.063e-06 $l=1.4e-07 $layer=LI1_cond $X=6.475 $Y=0.912
+ $X2=6.615 $Y2=0.912
r101 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.475 $Y=0.465
+ $X2=6.475 $Y2=0.465
r102 67 69 4.18122 $w=1.063e-06 $l=3.65e-07 $layer=LI1_cond $X=6.11 $Y=0.912
+ $X2=6.475 $Y2=0.912
r103 64 70 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.755 $Y=0.44
+ $X2=6.475 $Y2=0.44
r104 63 67 4.06667 $w=1.063e-06 $l=3.55e-07 $layer=LI1_cond $X=5.755 $Y=0.912
+ $X2=6.11 $Y2=0.912
r105 63 65 13.0357 $w=1.063e-06 $l=1.5e-07 $layer=LI1_cond $X=5.755 $Y=0.912
+ $X2=5.605 $Y2=0.912
r106 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.755 $Y=0.465
+ $X2=5.755 $Y2=0.465
r107 61 65 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.055 $Y=0.465
+ $X2=5.605 $Y2=0.465
r108 59 61 13.3793 $w=1.063e-06 $l=1.8e-07 $layer=LI1_cond $X=4.875 $Y=0.912
+ $X2=5.055 $Y2=0.912
r109 57 59 3.723 $w=1.063e-06 $l=3.25e-07 $layer=LI1_cond $X=4.55 $Y=0.912
+ $X2=4.875 $Y2=0.912
r110 53 57 4.52488 $w=1.063e-06 $l=3.95e-07 $layer=LI1_cond $X=4.155 $Y=0.912
+ $X2=4.55 $Y2=0.912
r111 53 55 12.5774 $w=1.063e-06 $l=1.1e-07 $layer=LI1_cond $X=4.155 $Y=0.912
+ $X2=4.045 $Y2=0.912
r112 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.155 $Y=0.465
+ $X2=4.155 $Y2=0.465
r113 49 54 0.28601 $w=3.7e-07 $l=7.45e-07 $layer=MET1_cond $X=3.41 $Y=0.44
+ $X2=4.155 $Y2=0.44
r114 47 49 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.69 $Y=0.44
+ $X2=3.41 $Y2=0.44
r115 46 51 7.36341 $w=7.87e-07 $l=4.75e-07 $layer=LI1_cond $X=3.05 $Y=0.465
+ $X2=3.05 $Y2=0.94
r116 46 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.41 $Y=0.465
+ $X2=3.41 $Y2=0.465
r117 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.69 $Y=0.465
+ $X2=2.69 $Y2=0.465
r118 43 47 0.32632 $w=3.7e-07 $l=8.5e-07 $layer=MET1_cond $X=1.84 $Y=0.44
+ $X2=2.69 $Y2=0.44
r119 42 44 11.907 $w=1.003e-06 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=0.882
+ $X2=1.925 $Y2=0.882
r120 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.84 $Y=0.465
+ $X2=1.84 $Y2=0.465
r121 40 42 7.64776 $w=1.003e-06 $l=6.3e-07 $layer=LI1_cond $X=1.21 $Y=0.882
+ $X2=1.84 $Y2=0.882
r122 37 43 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=0.76 $Y=0.44
+ $X2=1.84 $Y2=0.44
r123 36 40 5.46269 $w=1.003e-06 $l=4.5e-07 $layer=LI1_cond $X=0.76 $Y=0.882
+ $X2=1.21 $Y2=0.882
r124 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.76 $Y=0.465
+ $X2=0.76 $Y2=0.465
r125 33 64 0.36663 $w=3.7e-07 $l=9.55e-07 $layer=MET1_cond $X=4.8 $Y=0.44
+ $X2=5.755 $Y2=0.44
r126 33 54 0.247619 $w=3.7e-07 $l=6.45e-07 $layer=MET1_cond $X=4.8 $Y=0.44
+ $X2=4.155 $Y2=0.44
r127 33 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.875 $Y=0.465
+ $X2=4.875 $Y2=0.465
r128 29 85 5.23838 $w=2.18e-07 $l=1e-07 $layer=LI1_cond $X=9.32 $Y=0.49 $X2=9.42
+ $Y2=0.49
r129 29 83 18.6977 $w=2.18e-07 $l=3.45e-07 $layer=LI1_cond $X=9.32 $Y=0.49
+ $X2=8.975 $Y2=0.49
r130 29 31 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.32 $Y=0.6 $X2=9.32
+ $Y2=0.94
r131 22 46 10.0992 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=3.495 $Y=0.465
+ $X2=3.05 $Y2=0.465
r132 22 55 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.495 $Y=0.465
+ $X2=4.045 $Y2=0.465
r133 19 46 10.0992 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=2.605 $Y=0.465
+ $X2=3.05 $Y2=0.465
r134 19 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.605 $Y=0.465
+ $X2=1.925 $Y2=0.465
r135 6 31 91 $w=1.7e-07 $l=3.04672e-07 $layer=licon1_NDIFF $count=2 $X=9.09
+ $Y=0.705 $X2=9.25 $Y2=0.94
r136 5 77 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=7.53
+ $Y=0.705 $X2=7.67 $Y2=0.94
r137 4 67 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=5.97
+ $Y=0.705 $X2=6.11 $Y2=0.94
r138 3 57 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=4.41
+ $Y=0.705 $X2=4.55 $Y2=0.94
r139 2 51 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.705 $X2=2.99 $Y2=0.94
r140 1 40 91 $w=1.7e-07 $l=3.1229e-07 $layer=licon1_NDIFF $count=2 $X=1.03
+ $Y=0.705 $X2=1.21 $Y2=0.94
.ends

