* File: sky130_fd_sc_hvl__nand2_1.pxi.spice
* Created: Fri Aug 28 09:37:57 2020
* 
x_PM_SKY130_FD_SC_HVL__NAND2_1%VNB N_VNB_M1000_b VNB N_VNB_c_4_p VNB
+ PM_SKY130_FD_SC_HVL__NAND2_1%VNB
x_PM_SKY130_FD_SC_HVL__NAND2_1%VPB N_VPB_M1003_b VPB N_VPB_c_17_p VPB
+ PM_SKY130_FD_SC_HVL__NAND2_1%VPB
x_PM_SKY130_FD_SC_HVL__NAND2_1%B B B N_B_M1000_g N_B_c_36_n N_B_M1003_g
+ PM_SKY130_FD_SC_HVL__NAND2_1%B
x_PM_SKY130_FD_SC_HVL__NAND2_1%A N_A_M1001_g N_A_M1002_g A N_A_c_57_n
+ PM_SKY130_FD_SC_HVL__NAND2_1%A
x_PM_SKY130_FD_SC_HVL__NAND2_1%VPWR N_VPWR_M1003_s N_VPWR_M1002_d VPWR
+ N_VPWR_c_83_n N_VPWR_c_86_n N_VPWR_c_89_n PM_SKY130_FD_SC_HVL__NAND2_1%VPWR
x_PM_SKY130_FD_SC_HVL__NAND2_1%Y N_Y_M1001_d N_Y_M1003_d N_Y_c_105_n N_Y_c_106_n
+ N_Y_c_107_n N_Y_c_109_n Y PM_SKY130_FD_SC_HVL__NAND2_1%Y
x_PM_SKY130_FD_SC_HVL__NAND2_1%VGND N_VGND_M1000_s VGND N_VGND_c_142_n
+ PM_SKY130_FD_SC_HVL__NAND2_1%VGND
cc_1 N_VNB_M1000_b N_B_M1000_g 0.0902632f $X=-0.33 $Y=-0.265 $X2=0.915 $Y2=0.93
cc_2 N_VNB_M1000_b N_B_c_36_n 0.0234138f $X=-0.33 $Y=-0.265 $X2=0.85 $Y2=1.77
cc_3 N_VNB_M1000_b N_A_M1001_g 0.0543483f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_4 N_VNB_c_4_p N_A_M1001_g 0.00216445f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_5 N_VNB_M1000_b N_A_c_57_n 0.0878958f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_M1000_b N_Y_c_105_n 0.00161077f $X=-0.33 $Y=-0.265 $X2=0.85 $Y2=1.77
cc_7 N_VNB_M1000_b N_Y_c_106_n 0.00920162f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_8 N_VNB_M1000_b N_Y_c_107_n 0.0333398f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_c_4_p N_Y_c_107_n 7.98908e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_10 N_VNB_M1000_b N_Y_c_109_n 0.00304516f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_11 N_VNB_M1000_b VGND 0.0655937f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_12 N_VNB_c_4_p VGND 0.256671f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_13 N_VNB_M1000_b N_VGND_c_142_n 0.118788f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_14 N_VNB_c_4_p N_VGND_c_142_n 0.0037122f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_15 N_VPB_M1003_b N_B_M1000_g 0.0651567f $X=-0.33 $Y=1.885 $X2=0.915 $Y2=0.93
cc_16 VPB N_B_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.915 $Y2=0.93
cc_17 N_VPB_c_17_p N_B_M1000_g 0.0152133f $X=2.16 $Y=4.07 $X2=0.915 $Y2=0.93
cc_18 N_VPB_M1003_b N_B_c_36_n 0.00834617f $X=-0.33 $Y=1.885 $X2=0.85 $Y2=1.77
cc_19 N_VPB_M1003_b N_A_M1002_g 0.0408055f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_20 VPB N_A_M1002_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_21 N_VPB_c_17_p N_A_M1002_g 0.0160007f $X=2.16 $Y=4.07 $X2=0 $Y2=0
cc_22 N_VPB_M1003_b N_A_c_57_n 0.0447105f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_23 N_VPB_M1003_b N_VPWR_c_83_n 0.0826422f $X=-0.33 $Y=1.885 $X2=0.85 $Y2=1.77
cc_24 VPB N_VPWR_c_83_n 0.00355415f $X=0 $Y=3.955 $X2=0.85 $Y2=1.77
cc_25 N_VPB_c_17_p N_VPWR_c_83_n 0.0486145f $X=2.16 $Y=4.07 $X2=0.85 $Y2=1.77
cc_26 N_VPB_M1003_b N_VPWR_c_86_n 0.0599588f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_86_n 0.00229469f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_28 N_VPB_c_17_p N_VPWR_c_86_n 0.0299474f $X=2.16 $Y=4.07 $X2=0 $Y2=0
cc_29 N_VPB_M1003_b N_VPWR_c_89_n 0.0447872f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_89_n 0.254901f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_31 N_VPB_c_17_p N_VPWR_c_89_n 0.0107625f $X=2.16 $Y=4.07 $X2=0 $Y2=0
cc_32 N_VPB_M1003_b N_Y_c_105_n 0.00403398f $X=-0.33 $Y=1.885 $X2=0.85 $Y2=1.77
cc_33 VPB N_Y_c_105_n 8.01732e-19 $X=0 $Y=3.955 $X2=0.85 $Y2=1.77
cc_34 N_VPB_c_17_p N_Y_c_105_n 0.0130099f $X=2.16 $Y=4.07 $X2=0.85 $Y2=1.77
cc_35 N_B_M1000_g N_A_M1001_g 0.109336f $X=0.915 $Y=0.93 $X2=0 $Y2=0
cc_36 N_B_M1000_g N_A_M1002_g 0.0160832f $X=0.915 $Y=0.93 $X2=0 $Y2=0
cc_37 N_B_c_36_n N_A_c_57_n 2.87671e-19 $X=0.85 $Y=1.77 $X2=0 $Y2=0
cc_38 N_B_M1000_g N_VPWR_c_83_n 0.0800809f $X=0.915 $Y=0.93 $X2=0.24 $Y2=0
cc_39 N_B_c_36_n N_VPWR_c_83_n 0.0593454f $X=0.85 $Y=1.77 $X2=0.24 $Y2=0
cc_40 N_B_M1000_g N_VPWR_c_89_n 0.00832591f $X=0.915 $Y=0.93 $X2=1.2 $Y2=0.058
cc_41 N_B_M1000_g N_Y_c_105_n 0.0096147f $X=0.915 $Y=0.93 $X2=0 $Y2=0
cc_42 N_B_c_36_n N_Y_c_105_n 0.0170467f $X=0.85 $Y=1.77 $X2=0 $Y2=0
cc_43 N_B_M1000_g N_Y_c_107_n 3.99224e-19 $X=0.915 $Y=0.93 $X2=0 $Y2=0
cc_44 N_B_M1000_g N_Y_c_109_n 0.00199143f $X=0.915 $Y=0.93 $X2=0 $Y2=0
cc_45 N_B_c_36_n N_Y_c_109_n 0.0109158f $X=0.85 $Y=1.77 $X2=0 $Y2=0
cc_46 N_B_M1000_g Y 8.67381e-19 $X=0.915 $Y=0.93 $X2=0 $Y2=0
cc_47 N_B_M1000_g N_VGND_c_142_n 0.0790812f $X=0.915 $Y=0.93 $X2=0 $Y2=0
cc_48 N_B_c_36_n N_VGND_c_142_n 0.0666291f $X=0.85 $Y=1.77 $X2=0 $Y2=0
cc_49 N_A_M1002_g N_VPWR_c_83_n 6.71148e-19 $X=1.695 $Y=2.965 $X2=0.24 $Y2=0
cc_50 N_A_M1002_g N_VPWR_c_86_n 0.0788889f $X=1.695 $Y=2.965 $X2=0 $Y2=0
cc_51 A N_VPWR_c_86_n 0.0144202f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_52 N_A_c_57_n N_VPWR_c_86_n 0.0103641f $X=2.11 $Y=1.69 $X2=0 $Y2=0
cc_53 N_A_M1002_g N_VPWR_c_89_n 0.011025f $X=1.695 $Y=2.965 $X2=1.2 $Y2=0.058
cc_54 N_A_M1002_g N_Y_c_105_n 0.0311988f $X=1.695 $Y=2.965 $X2=0 $Y2=0
cc_55 A N_Y_c_105_n 0.00478116f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_56 N_A_c_57_n N_Y_c_105_n 0.0224603f $X=2.11 $Y=1.69 $X2=0 $Y2=0
cc_57 N_A_M1001_g N_Y_c_106_n 0.0183129f $X=1.625 $Y=0.93 $X2=0 $Y2=0
cc_58 A N_Y_c_106_n 0.0147557f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_59 N_A_c_57_n N_Y_c_106_n 0.0103473f $X=2.11 $Y=1.69 $X2=0 $Y2=0
cc_60 N_A_M1001_g N_Y_c_107_n 0.0191905f $X=1.625 $Y=0.93 $X2=0 $Y2=0
cc_61 A N_Y_c_109_n 0.0126108f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_62 N_A_c_57_n N_Y_c_109_n 0.0311182f $X=2.11 $Y=1.69 $X2=0 $Y2=0
cc_63 N_A_M1001_g Y 0.00729931f $X=1.625 $Y=0.93 $X2=0 $Y2=0
cc_64 N_A_c_57_n Y 0.0077608f $X=2.11 $Y=1.69 $X2=0 $Y2=0
cc_65 N_A_M1001_g VGND 0.020998f $X=1.625 $Y=0.93 $X2=0 $Y2=0
cc_66 N_A_M1001_g N_VGND_c_142_n 0.0312783f $X=1.625 $Y=0.93 $X2=0 $Y2=0
cc_67 N_VPWR_c_89_n N_Y_M1003_d 0.00221032f $X=2.135 $Y=3.59 $X2=0 $Y2=0
cc_68 N_VPWR_c_83_n N_Y_c_105_n 0.0677867f $X=0.525 $Y=2.34 $X2=0.24 $Y2=4.07
cc_69 N_VPWR_c_86_n N_Y_c_105_n 0.107316f $X=2.085 $Y=2.34 $X2=0.24 $Y2=4.07
cc_70 N_VPWR_c_89_n N_Y_c_105_n 0.0306945f $X=2.135 $Y=3.59 $X2=0.24 $Y2=4.07
cc_71 N_VPWR_c_86_n N_Y_c_109_n 0.0043611f $X=2.085 $Y=2.34 $X2=1.2 $Y2=4.013
cc_72 N_Y_c_106_n VGND 0.00817002f $X=2.015 $Y=1.175 $X2=0 $Y2=0
cc_73 N_Y_c_107_n VGND 0.0214014f $X=2.015 $Y=0.68 $X2=0 $Y2=0
cc_74 N_Y_c_106_n N_VGND_c_142_n 0.0133884f $X=2.015 $Y=1.175 $X2=0 $Y2=0
cc_75 N_Y_c_107_n N_VGND_c_142_n 0.0219255f $X=2.015 $Y=0.68 $X2=0 $Y2=0
cc_76 N_Y_c_109_n N_VGND_c_142_n 0.0143171f $X=1.687 $Y=1.525 $X2=0 $Y2=0
