* File: sky130_fd_sc_hvl__inv_1.pex.spice
* Created: Wed Sep  2 09:06:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__INV_1%VNB 5 7 11 25
r10 7 25 8.85771e-05 $w=1.44e-06 $l=1e-09 $layer=MET1_cond $X=0.72 $Y=0.057
+ $X2=0.72 $Y2=0.058
r11 7 11 0.00504889 $w=1.44e-06 $l=5.7e-08 $layer=MET1_cond $X=0.72 $Y=0.057
+ $X2=0.72 $Y2=0
r12 5 11 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r13 5 11 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_1%VPB 4 6 14 21
r16 10 21 0.00504889 $w=1.44e-06 $l=5.7e-08 $layer=MET1_cond $X=0.72 $Y=4.07
+ $X2=0.72 $Y2=4.013
r17 10 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=4.07 $X2=1.2
+ $Y2=4.07
r18 9 14 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=1.2
+ $Y2=4.07
r19 9 10 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r20 6 21 8.85771e-05 $w=1.44e-06 $l=1e-09 $layer=MET1_cond $X=0.72 $Y=4.012
+ $X2=0.72 $Y2=4.013
r21 4 14 121.333 $w=1.7e-07 $l=1.24177e-06 $layer=licon1_NTAP_notbjt $count=1
+ $X=0 $Y=3.985 $X2=1.2 $Y2=4.07
r22 4 9 121.333 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_1%A 3 7 9 10 14
r22 14 17 32.4104 $w=5.2e-07 $l=3.15e-07 $layer=POLY_cond $X=0.745 $Y=1.77
+ $X2=0.745 $Y2=2.085
r23 14 16 36.5261 $w=5.2e-07 $l=3.55e-07 $layer=POLY_cond $X=0.745 $Y=1.77
+ $X2=0.745 $Y2=1.415
r24 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.77 $X2=0.67 $Y2=1.77
r25 10 15 1.49668 $w=3.83e-07 $l=5e-08 $layer=LI1_cond $X=0.72 $Y=1.742 $X2=0.67
+ $Y2=1.742
r26 9 15 12.8714 $w=3.83e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=1.742
+ $X2=0.67 $Y2=1.742
r27 7 16 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.755 $Y=0.91 $X2=0.755
+ $Y2=1.415
r28 3 17 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.735 $Y=2.965
+ $X2=0.735 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_1%VPWR 1 4 7
r11 10 12 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.565 $Y=3.59
+ $X2=0.565 $Y2=3.59
r12 7 10 25.3406 $w=5.88e-07 $l=1.25e-06 $layer=LI1_cond $X=0.385 $Y=2.34
+ $X2=0.385 $Y2=3.59
r13 4 12 0.0595053 $w=3.7e-07 $l=1.55e-07 $layer=MET1_cond $X=0.72 $Y=3.63
+ $X2=0.565 $Y2=3.63
r14 1 10 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.2
+ $Y=2.215 $X2=0.345 $Y2=3.59
r15 1 7 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.2
+ $Y=2.215 $X2=0.345 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_1%Y 1 2 7 8 9 10 11 12 13 24 36
r18 34 36 1.13748 $w=3.83e-07 $l=3.8e-08 $layer=LI1_cond $X=1.152 $Y=2.367
+ $X2=1.152 $Y2=2.405
r19 13 43 13.3204 $w=3.83e-07 $l=4.45e-07 $layer=LI1_cond $X=1.152 $Y=3.145
+ $X2=1.152 $Y2=3.59
r20 12 13 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.152 $Y=2.775
+ $X2=1.152 $Y2=3.145
r21 11 34 0.808207 $w=3.83e-07 $l=2.7e-08 $layer=LI1_cond $X=1.152 $Y=2.34
+ $X2=1.152 $Y2=2.367
r22 11 47 5.20661 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.152 $Y=2.34
+ $X2=1.152 $Y2=2.175
r23 11 12 10.387 $w=3.83e-07 $l=3.47e-07 $layer=LI1_cond $X=1.152 $Y=2.428
+ $X2=1.152 $Y2=2.775
r24 11 36 0.688472 $w=3.83e-07 $l=2.3e-08 $layer=LI1_cond $X=1.152 $Y=2.428
+ $X2=1.152 $Y2=2.405
r25 10 47 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.18 $Y=2.035
+ $X2=1.18 $Y2=2.175
r26 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=1.665
+ $X2=1.18 $Y2=2.035
r27 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=1.295 $X2=1.18
+ $Y2=1.665
r28 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=0.925 $X2=1.18
+ $Y2=1.295
r29 7 24 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.18 $Y=0.925
+ $X2=1.18 $Y2=0.66
r30 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=2.215 $X2=1.125 $Y2=2.34
r31 2 43 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=2.215 $X2=1.125 $Y2=3.59
r32 1 24 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.005
+ $Y=0.535 $X2=1.145 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_1%VGND 1 4 7
r11 7 11 3.64905 $w=5.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.385 $Y=0.48
+ $X2=0.385 $Y2=0.66
r12 7 8 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.565 $Y=0.48
+ $X2=0.565 $Y2=0.48
r13 4 8 0.0595053 $w=3.7e-07 $l=1.55e-07 $layer=MET1_cond $X=0.72 $Y=0.44
+ $X2=0.565 $Y2=0.44
r14 1 11 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.22
+ $Y=0.535 $X2=0.365 $Y2=0.66
.ends

