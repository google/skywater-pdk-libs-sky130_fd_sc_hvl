* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__buf_2 A VGND VNB VPB VPWR X
*.PININFO A:I VGND:I VNB:I VPB:I VPWR:I X:O
MMIN1 Ab A VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MMIN2 X Ab VNB nhv m=2 w=0.75 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MMIP1 Ab A VPB phv m=1 w=0.75 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MMIP2 X Ab VPB phv m=2 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_hvl__buf_2
