* File: sky130_fd_sc_hvl__lsbuflv2hv_1.spice
* Created: Wed Sep  2 09:07:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__lsbuflv2hv_1.pex.spice"
.subckt sky130_fd_sc_hvl__lsbuflv2hv_1  VNB VPB LVPWR A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* LVPWR	LVPWR
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_A_M1014_g N_A_404_1133#_M1014_s N_VNB_M1014_b NSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2478 PD=1.12 PS=2.27 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1015 N_A_772_151#_M1015_d N_A_404_1133#_M1015_g N_VGND_M1014_d N_VNB_M1014_b
+ NSHORT L=0.15 W=0.84 AD=0.2478 AS=0.1176 PD=2.27 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_A_404_1133#_M1002_g N_A_504_1221#_M1002_s N_VNB_M1014_b
+ NHV L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 M=1 R=3
+ SA=250000 SB=250003 A=0.75 P=4 MULT=1
MM1003 N_VGND_M1003_d N_A_404_1133#_M1003_g N_A_504_1221#_M1002_s N_VNB_M1014_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001
+ SB=250002 A=0.75 P=4 MULT=1
MM1008 N_VGND_M1003_d N_A_404_1133#_M1008_g N_A_504_1221#_M1008_s N_VNB_M1014_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002
+ SB=250002 A=0.75 P=4 MULT=1
MM1010 N_VGND_M1010_d N_A_404_1133#_M1010_g N_A_504_1221#_M1008_s N_VNB_M1014_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002
+ SB=250001 A=0.75 P=4 MULT=1
MM1011 N_VGND_M1010_d N_A_404_1133#_M1011_g N_A_504_1221#_M1011_s N_VNB_M1014_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 M=1 R=3
+ SA=250003 SB=250000 A=0.75 P=4 MULT=1
MM1000 N_A_1197_107#_M1000_d N_A_772_151#_M1000_g N_VGND_M1000_s N_VNB_M1014_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 M=1 R=3
+ SA=250000 SB=250003 A=0.75 P=4 MULT=1
MM1007 N_A_1197_107#_M1000_d N_A_772_151#_M1007_g N_VGND_M1007_s N_VNB_M1014_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001
+ SB=250002 A=0.75 P=4 MULT=1
MM1009 N_A_1197_107#_M1009_d N_A_772_151#_M1009_g N_VGND_M1007_s N_VNB_M1014_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002
+ SB=250002 A=0.75 P=4 MULT=1
MM1012 N_A_1197_107#_M1009_d N_A_772_151#_M1012_g N_VGND_M1012_s N_VNB_M1014_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002
+ SB=250001 A=0.75 P=4 MULT=1
MM1019 N_A_1197_107#_M1019_d N_A_772_151#_M1019_g N_VGND_M1012_s N_VNB_M1014_b
+ NHV L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 M=1 R=3
+ SA=250003 SB=250000 A=0.75 P=4 MULT=1
MM1016 N_VGND_M1016_d N_A_504_1221#_M1016_g N_A_1711_885#_M1016_s N_VNB_M1014_b
+ NHV L=0.5 W=0.75 AD=0.121875 AS=0.19875 PD=1.075 PS=2.03 NRD=6.8286 NRS=0 M=1
+ R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1005 N_X_M1005_d N_A_1711_885#_M1005_g N_VGND_M1016_d N_VNB_M1014_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.121875 PD=2.03 PS=1.075 NRD=0 NRS=0 M=1 R=1.5 SA=250001
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1004 N_LVPWR_M1004_d N_A_M1004_g N_A_404_1133#_M1004_s N_LVPWR_M1004_b PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2478 PD=1.12 PS=2.27 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1017 N_A_772_151#_M1017_d N_A_404_1133#_M1017_g N_LVPWR_M1004_d
+ N_LVPWR_M1004_b PHIGHVT L=0.15 W=0.84 AD=0.2478 AS=0.1176 PD=2.27 PS=1.12
+ NRD=0 NRS=0 M=1 R=5.6 SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1018 N_VPWR_M1018_d N_A_504_1221#_M1018_g N_A_1197_107#_M1018_s N_VPB_M1018_b
+ PHV L=1 W=0.42 AD=0.1113 AS=0.1365 PD=1.37 PS=1.49 NRD=0 NRS=0 M=1 R=0.42
+ SA=500000 SB=500000 A=0.42 P=2.84 MULT=1
MM1006 N_VPWR_M1006_d N_A_1197_107#_M1006_g N_A_504_1221#_M1006_s N_VPB_M1018_b
+ PHV L=1 W=0.42 AD=0.2142 AS=0.2142 PD=1.99 PS=1.99 NRD=14.7643 NRS=14.7643 M=1
+ R=0.42 SA=500000 SB=500000 A=0.42 P=2.84 MULT=1
MM1013 N_VPWR_M1013_d N_A_504_1221#_M1013_g N_A_1711_885#_M1013_s N_VPB_M1018_b
+ PHV L=0.5 W=1.5 AD=0.24375 AS=0.3975 PD=1.825 PS=3.53 NRD=5.7109 NRS=0 M=1 R=3
+ SA=250000 SB=250001 A=0.75 P=4 MULT=1
MM1001 N_X_M1001_d N_A_1711_885#_M1001_g N_VPWR_M1013_d N_VPB_M1018_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.24375 PD=3.53 PS=1.825 NRD=0 NRS=0 M=1 R=3 SA=250001
+ SB=250000 A=0.75 P=4 MULT=1
DX20_noxref N_VNB_M1014_b N_VPB_X20_noxref_D1 NWDIODE A=4.9381 P=11
DX21_noxref N_VNB_M1014_b N_LVPWR_M1004_b NWDIODE A=3.54585 P=7.69
DX22_noxref N_VNB_M1014_b N_VPB_M1018_b NWDIODE A=17.8956 P=17.85
*
.include "sky130_fd_sc_hvl__lsbuflv2hv_1.pxi.spice"
*
.ends
*
*
