/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_HVL__UDP_ISOLATCHHV_PP_PLG_S_TB_V
`define SKY130_FD_SC_HVL__UDP_ISOLATCHHV_PP_PLG_S_TB_V

/**
 * udp_isolatchhv_pp$PLG$S: Power isolating latch (for HV). Includes
 *                          VPWR, LVPWR, and VGND power pins with
 *                          active high sleep pin (SLEEP).
 *
 * Autogenerated test bench.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

`include "sky130_fd_sc_hvl__udp_isolatchhv_pp_plg_s.v"

module top();

    // Inputs are registered
    reg UDP_IN;
    reg VPWR;
    reg LVPWR;
    reg VGND;
    reg SLEEP;

    // Outputs are wires
    wire UDP_OUT;

    initial
    begin
        // Initial state is x for all inputs.
        LVPWR  = 1'bX;
        SLEEP  = 1'bX;
        UDP_IN = 1'bX;
        VGND   = 1'bX;
        VPWR   = 1'bX;

        #20   LVPWR  = 1'b0;
        #40   SLEEP  = 1'b0;
        #60   UDP_IN = 1'b0;
        #80   VGND   = 1'b0;
        #100  VPWR   = 1'b0;
        #120  LVPWR  = 1'b1;
        #140  SLEEP  = 1'b1;
        #160  UDP_IN = 1'b1;
        #180  VGND   = 1'b1;
        #200  VPWR   = 1'b1;
        #220  LVPWR  = 1'b0;
        #240  SLEEP  = 1'b0;
        #260  UDP_IN = 1'b0;
        #280  VGND   = 1'b0;
        #300  VPWR   = 1'b0;
        #320  VPWR   = 1'b1;
        #340  VGND   = 1'b1;
        #360  UDP_IN = 1'b1;
        #380  SLEEP  = 1'b1;
        #400  LVPWR  = 1'b1;
        #420  VPWR   = 1'bx;
        #440  VGND   = 1'bx;
        #460  UDP_IN = 1'bx;
        #480  SLEEP  = 1'bx;
        #500  LVPWR  = 1'bx;
    end

    sky130_fd_sc_hvl__udp_isolatchhv_pp$PLG$S dut (.UDP_IN(UDP_IN), .VPWR(VPWR), .LVPWR(LVPWR), .VGND(VGND), .SLEEP(SLEEP), .UDP_OUT(UDP_OUT));

endmodule

`default_nettype wire
`endif  // SKY130_FD_SC_HVL__UDP_ISOLATCHHV_PP_PLG_S_TB_V
