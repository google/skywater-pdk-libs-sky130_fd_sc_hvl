# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__probec_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__probec_p_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  3.375000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.580000 2.245000 1.815000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.520000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.410000 1.445000 3.590000 2.625000 ;
        RECT 5.010000 1.445000 6.190000 2.625000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.290000  1.235000 6.310000 2.835000 ;
        RECT 4.710000 -0.365000 6.310000 1.235000 ;
        RECT 4.710000  2.835000 6.310000 4.435000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 7.910000 -0.365000 10.410000 1.235000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 9.600000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 9.600000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 9.600000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 9.930000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 7.910000 2.835000 10.410000 4.435000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.985000 9.600000 4.155000 ;
      RECT 0.245000  0.805000 0.455000 1.475000 ;
      RECT 0.245000  1.475000 0.435000 2.095000 ;
      RECT 0.245000  2.095000 2.595000 2.265000 ;
      RECT 0.245000  2.265000 0.435000 3.545000 ;
      RECT 0.615000  2.445000 1.865000 3.625000 ;
      RECT 0.615000  3.625000 9.505000 3.795000 ;
      RECT 0.675000  0.380000 9.505000 0.550000 ;
      RECT 0.675000  0.550000 1.925000 1.385000 ;
      RECT 2.045000  2.265000 2.595000 3.445000 ;
      RECT 2.105000  0.730000 2.315000 1.230000 ;
      RECT 2.105000  1.230000 2.595000 1.400000 ;
      RECT 2.425000  1.400000 2.595000 1.625000 ;
      RECT 2.425000  1.625000 3.380000 1.955000 ;
      RECT 2.425000  1.955000 2.595000 2.095000 ;
      RECT 2.605000  0.550000 3.495000 0.760000 ;
      RECT 2.765000  0.760000 3.495000 1.445000 ;
      RECT 2.765000  2.385000 3.435000 3.625000 ;
      RECT 3.605000  1.955000 8.965000 2.205000 ;
      RECT 3.605000  2.205000 3.935000 3.445000 ;
      RECT 3.665000  0.805000 3.875000 1.625000 ;
      RECT 3.665000  1.625000 8.965000 1.955000 ;
      RECT 4.045000  0.550000 5.055000 1.445000 ;
      RECT 4.105000  2.385000 4.995000 3.625000 ;
      RECT 5.165000  2.205000 5.495000 3.445000 ;
      RECT 5.225000  0.805000 5.435000 1.625000 ;
      RECT 5.605000  0.550000 6.615000 1.445000 ;
      RECT 5.665000  2.385000 6.555000 3.625000 ;
      RECT 6.725000  2.205000 7.055000 3.445000 ;
      RECT 6.785000  0.805000 6.995000 1.625000 ;
      RECT 7.165000  0.550000 8.175000 1.445000 ;
      RECT 7.225000  2.385000 8.115000 3.625000 ;
      RECT 8.285000  2.205000 8.965000 3.230000 ;
      RECT 8.285000  3.230000 8.735000 3.445000 ;
      RECT 8.345000  0.805000 8.965000 1.625000 ;
      RECT 8.905000  3.475000 9.505000 3.625000 ;
      RECT 8.975000  0.550000 9.505000 0.600000 ;
      RECT 9.135000  0.600000 9.505000 1.445000 ;
      RECT 9.135000  2.385000 9.505000 3.475000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.615000  3.475000 0.785000 3.645000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.975000  3.475000 1.145000 3.645000 ;
      RECT 1.035000  0.380000 1.205000 0.550000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.335000  3.475000 1.505000 3.645000 ;
      RECT 1.395000  0.380000 1.565000 0.550000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.695000  3.475000 1.865000 3.645000 ;
      RECT 1.755000  0.380000 1.925000 0.550000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.605000  0.380000 2.775000 0.550000 ;
      RECT 2.770000  3.475000 2.940000 3.645000 ;
      RECT 2.965000  0.380000 3.135000 0.550000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.130000  3.475000 3.300000 3.645000 ;
      RECT 3.325000  0.380000 3.495000 0.550000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.070000  0.380000 4.240000 0.550000 ;
      RECT 4.105000  3.475000 4.275000 3.645000 ;
      RECT 4.430000  0.380000 4.600000 0.550000 ;
      RECT 4.465000  3.475000 4.635000 3.645000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.790000  0.380000 4.960000 0.550000 ;
      RECT 4.825000  3.475000 4.995000 3.645000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.985000 5.605000 4.155000 ;
      RECT 5.620000  1.950000 5.790000 2.120000 ;
      RECT 5.665000  3.475000 5.835000 3.645000 ;
      RECT 5.670000  0.380000 5.840000 0.550000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.985000 6.085000 4.155000 ;
      RECT 5.980000  1.950000 6.150000 2.120000 ;
      RECT 6.025000  3.475000 6.195000 3.645000 ;
      RECT 6.030000  0.380000 6.200000 0.550000 ;
      RECT 6.385000  3.475000 6.555000 3.645000 ;
      RECT 6.390000  0.380000 6.560000 0.550000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.985000 6.565000 4.155000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.985000 7.045000 4.155000 ;
      RECT 7.230000  3.475000 7.400000 3.645000 ;
      RECT 7.235000  0.380000 7.405000 0.550000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.595000  0.380000 7.765000 0.550000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 7.945000  3.475000 8.115000 3.645000 ;
      RECT 7.955000  0.380000 8.125000 0.550000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.985000 8.485000 4.155000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.985000 8.965000 4.155000 ;
      RECT 8.975000  0.380000 9.145000 0.550000 ;
      RECT 9.265000  3.475000 9.435000 3.645000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.985000 9.445000 4.155000 ;
      RECT 9.335000  0.380000 9.505000 0.550000 ;
    LAYER met1 ;
      RECT 0.000000 0.255000 9.600000 0.305000 ;
      RECT 0.000000 0.305000 9.920000 0.565000 ;
      RECT 0.000000 0.565000 9.600000 0.625000 ;
      RECT 0.000000 3.445000 9.600000 3.505000 ;
      RECT 0.000000 3.505000 9.920000 3.765000 ;
      RECT 0.000000 3.765000 9.600000 3.815000 ;
      RECT 5.560000 1.905000 6.210000 2.165000 ;
    LAYER met2 ;
      RECT 5.440000 1.895000 6.210000 2.175000 ;
      RECT 9.215000 0.285000 9.985000 0.565000 ;
      RECT 9.215000 3.505000 9.985000 3.785000 ;
    LAYER met3 ;
      RECT 2.835000 1.875000 3.615000 2.195000 ;
      RECT 5.435000 1.870000 6.215000 2.200000 ;
      RECT 9.210000 0.260000 9.990000 0.590000 ;
      RECT 9.210000 3.480000 9.990000 3.810000 ;
    LAYER met4 ;
      RECT 9.010000 -0.155000 10.190000 1.025000 ;
      RECT 9.010000  3.045000 10.190000 4.225000 ;
    LAYER via ;
      RECT 5.600000 1.905000 5.860000 2.165000 ;
      RECT 5.920000 1.905000 6.180000 2.165000 ;
      RECT 9.310000 0.305000 9.570000 0.565000 ;
      RECT 9.310000 3.505000 9.570000 3.765000 ;
      RECT 9.630000 0.305000 9.890000 0.565000 ;
      RECT 9.630000 3.505000 9.890000 3.765000 ;
    LAYER via2 ;
      RECT 5.485000 1.895000 5.765000 2.175000 ;
      RECT 5.885000 1.895000 6.165000 2.175000 ;
      RECT 9.260000 0.285000 9.540000 0.565000 ;
      RECT 9.260000 3.505000 9.540000 3.785000 ;
      RECT 9.660000 0.285000 9.940000 0.565000 ;
      RECT 9.660000 3.505000 9.940000 3.785000 ;
    LAYER via3 ;
      RECT 2.865000 1.875000 3.185000 2.195000 ;
      RECT 3.265000 1.875000 3.585000 2.195000 ;
      RECT 5.465000 1.875000 5.785000 2.195000 ;
      RECT 5.865000 1.875000 6.185000 2.195000 ;
      RECT 9.240000 0.265000 9.560000 0.585000 ;
      RECT 9.240000 3.485000 9.560000 3.805000 ;
      RECT 9.640000 0.265000 9.960000 0.585000 ;
      RECT 9.640000 3.485000 9.960000 3.805000 ;
  END
END sky130_fd_sc_hvl__probec_p_8
END LIBRARY
