* File: sky130_fd_sc_hvl__buf_32.pxi.spice
* Created: Wed Sep  2 09:04:12 2020
* 
x_PM_SKY130_FD_SC_HVL__BUF_32%VNB N_VNB_M1008_b VNB N_VNB_c_2_p VNB VNB
+ PM_SKY130_FD_SC_HVL__BUF_32%VNB
x_PM_SKY130_FD_SC_HVL__BUF_32%VPB N_VPB_M1000_b VPB N_VPB_c_156_p N_VPB_c_157_p
+ VPB VPB PM_SKY130_FD_SC_HVL__BUF_32%VPB
x_PM_SKY130_FD_SC_HVL__BUF_32%A N_A_c_411_n N_A_M1008_g N_A_M1000_g N_A_c_413_n
+ N_A_M1012_g N_A_M1001_g N_A_c_415_n N_A_M1027_g N_A_M1006_g N_A_c_417_n
+ N_A_M1028_g N_A_M1016_g N_A_c_419_n N_A_M1032_g N_A_M1019_g N_A_c_421_n
+ N_A_M1043_g N_A_M1035_g N_A_c_423_n N_A_M1051_g N_A_M1039_g N_A_c_425_n
+ N_A_M1069_g N_A_M1049_g N_A_c_427_n N_A_M1074_g N_A_M1064_g N_A_c_429_n
+ N_A_M1081_g N_A_M1070_g A A A A A A A N_A_c_431_n N_A_c_432_n
+ PM_SKY130_FD_SC_HVL__BUF_32%A
x_PM_SKY130_FD_SC_HVL__BUF_32%A_183_141# N_A_183_141#_M1008_s
+ N_A_183_141#_M1027_s N_A_183_141#_M1032_s N_A_183_141#_M1051_s
+ N_A_183_141#_M1074_s N_A_183_141#_M1000_s N_A_183_141#_M1006_s
+ N_A_183_141#_M1019_s N_A_183_141#_M1039_s N_A_183_141#_M1064_s
+ N_A_183_141#_c_614_n N_A_183_141#_M1002_g N_A_183_141#_M1004_g
+ N_A_183_141#_c_616_n N_A_183_141#_M1003_g N_A_183_141#_M1011_g
+ N_A_183_141#_c_618_n N_A_183_141#_M1005_g N_A_183_141#_M1013_g
+ N_A_183_141#_c_620_n N_A_183_141#_M1007_g N_A_183_141#_M1017_g
+ N_A_183_141#_c_622_n N_A_183_141#_M1009_g N_A_183_141#_M1018_g
+ N_A_183_141#_c_624_n N_A_183_141#_M1010_g N_A_183_141#_M1020_g
+ N_A_183_141#_c_626_n N_A_183_141#_M1014_g N_A_183_141#_M1021_g
+ N_A_183_141#_c_628_n N_A_183_141#_M1015_g N_A_183_141#_M1022_g
+ N_A_183_141#_c_630_n N_A_183_141#_M1025_g N_A_183_141#_M1023_g
+ N_A_183_141#_c_632_n N_A_183_141#_M1031_g N_A_183_141#_M1024_g
+ N_A_183_141#_c_634_n N_A_183_141#_M1038_g N_A_183_141#_M1026_g
+ N_A_183_141#_c_636_n N_A_183_141#_M1040_g N_A_183_141#_M1029_g
+ N_A_183_141#_c_638_n N_A_183_141#_M1044_g N_A_183_141#_M1030_g
+ N_A_183_141#_c_640_n N_A_183_141#_M1047_g N_A_183_141#_M1033_g
+ N_A_183_141#_c_642_n N_A_183_141#_M1048_g N_A_183_141#_M1034_g
+ N_A_183_141#_c_644_n N_A_183_141#_M1052_g N_A_183_141#_M1036_g
+ N_A_183_141#_c_646_n N_A_183_141#_M1053_g N_A_183_141#_M1037_g
+ N_A_183_141#_c_648_n N_A_183_141#_M1056_g N_A_183_141#_M1041_g
+ N_A_183_141#_c_650_n N_A_183_141#_M1057_g N_A_183_141#_M1042_g
+ N_A_183_141#_c_652_n N_A_183_141#_M1058_g N_A_183_141#_M1045_g
+ N_A_183_141#_c_654_n N_A_183_141#_M1061_g N_A_183_141#_M1046_g
+ N_A_183_141#_c_656_n N_A_183_141#_M1062_g N_A_183_141#_M1050_g
+ N_A_183_141#_c_658_n N_A_183_141#_M1067_g N_A_183_141#_M1054_g
+ N_A_183_141#_c_660_n N_A_183_141#_M1068_g N_A_183_141#_M1055_g
+ N_A_183_141#_c_662_n N_A_183_141#_M1071_g N_A_183_141#_M1059_g
+ N_A_183_141#_c_664_n N_A_183_141#_M1072_g N_A_183_141#_M1060_g
+ N_A_183_141#_c_666_n N_A_183_141#_M1076_g N_A_183_141#_M1063_g
+ N_A_183_141#_c_668_n N_A_183_141#_M1077_g N_A_183_141#_M1065_g
+ N_A_183_141#_c_670_n N_A_183_141#_M1078_g N_A_183_141#_M1066_g
+ N_A_183_141#_c_672_n N_A_183_141#_M1079_g N_A_183_141#_M1073_g
+ N_A_183_141#_c_674_n N_A_183_141#_M1082_g N_A_183_141#_M1075_g
+ N_A_183_141#_c_676_n N_A_183_141#_M1083_g N_A_183_141#_M1080_g
+ N_A_183_141#_c_678_n N_A_183_141#_c_797_n N_A_183_141#_c_819_n
+ N_A_183_141#_c_823_n N_A_183_141#_c_826_n N_A_183_141#_c_830_n
+ N_A_183_141#_c_679_n N_A_183_141#_c_800_n N_A_183_141#_c_837_n
+ N_A_183_141#_c_841_n N_A_183_141#_c_803_n N_A_183_141#_c_680_n
+ N_A_183_141#_c_849_n N_A_183_141#_c_851_n N_A_183_141#_c_681_n
+ N_A_183_141#_c_806_n N_A_183_141#_c_860_n N_A_183_141#_c_865_n
+ N_A_183_141#_c_809_n N_A_183_141#_c_682_n N_A_183_141#_c_877_n
+ N_A_183_141#_c_881_n N_A_183_141#_c_884_n N_A_183_141#_c_887_n
+ N_A_183_141#_c_683_n N_A_183_141#_c_684_n N_A_183_141#_c_685_n
+ N_A_183_141#_c_686_n N_A_183_141#_c_687_n N_A_183_141#_c_688_n
+ N_A_183_141#_c_689_n N_A_183_141#_c_690_n N_A_183_141#_c_691_n
+ N_A_183_141#_c_692_n N_A_183_141#_c_693_n N_A_183_141#_c_694_n
+ N_A_183_141#_c_695_n N_A_183_141#_c_696_n N_A_183_141#_c_697_n
+ N_A_183_141#_c_698_n N_A_183_141#_c_699_n
+ PM_SKY130_FD_SC_HVL__BUF_32%A_183_141#
x_PM_SKY130_FD_SC_HVL__BUF_32%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_M1016_d
+ N_VPWR_M1035_d N_VPWR_M1049_d N_VPWR_M1070_d N_VPWR_M1011_d N_VPWR_M1017_d
+ N_VPWR_M1020_d N_VPWR_M1022_d N_VPWR_M1024_d N_VPWR_M1029_d N_VPWR_M1033_d
+ N_VPWR_M1036_d N_VPWR_M1041_d N_VPWR_M1045_d N_VPWR_M1050_d N_VPWR_M1055_d
+ N_VPWR_M1060_d N_VPWR_M1065_d N_VPWR_M1073_d N_VPWR_M1080_d VPWR
+ N_VPWR_c_1410_n N_VPWR_c_1413_n N_VPWR_c_1415_n N_VPWR_c_1417_n
+ N_VPWR_c_1419_n N_VPWR_c_1421_n N_VPWR_c_1423_n N_VPWR_c_1426_n
+ N_VPWR_c_1429_n N_VPWR_c_1432_n N_VPWR_c_1435_n N_VPWR_c_1438_n
+ N_VPWR_c_1441_n N_VPWR_c_1444_n N_VPWR_c_1447_n N_VPWR_c_1450_n
+ N_VPWR_c_1453_n N_VPWR_c_1456_n N_VPWR_c_1459_n N_VPWR_c_1462_n
+ N_VPWR_c_1465_n N_VPWR_c_1468_n N_VPWR_c_1471_n VPWR
+ PM_SKY130_FD_SC_HVL__BUF_32%VPWR
x_PM_SKY130_FD_SC_HVL__BUF_32%X N_X_M1002_d N_X_M1005_d N_X_M1009_d N_X_M1014_d
+ N_X_M1025_d N_X_M1038_d N_X_M1044_d N_X_M1048_d N_X_M1053_d N_X_M1057_d
+ N_X_M1061_d N_X_M1067_d N_X_M1071_d N_X_M1076_d N_X_M1078_d N_X_M1082_d
+ N_X_M1004_s N_X_M1013_s N_X_M1018_s N_X_M1021_s N_X_M1023_s N_X_M1026_s
+ N_X_M1030_s N_X_M1034_s N_X_M1037_s N_X_M1042_s N_X_M1046_s N_X_M1054_s
+ N_X_M1059_s N_X_M1063_s N_X_M1066_s N_X_M1075_s X N_X_c_1741_n N_X_c_1744_n
+ N_X_c_1747_n N_X_c_1750_n N_X_c_1753_n N_X_c_1756_n N_X_c_1759_n N_X_c_1762_n
+ N_X_c_1765_n N_X_c_1768_n N_X_c_1771_n N_X_c_1774_n N_X_c_1777_n N_X_c_1780_n
+ N_X_c_1783_n N_X_c_1786_n N_X_c_1916_n X PM_SKY130_FD_SC_HVL__BUF_32%X
x_PM_SKY130_FD_SC_HVL__BUF_32%VGND N_VGND_M1008_d N_VGND_M1012_d N_VGND_M1028_d
+ N_VGND_M1043_d N_VGND_M1069_d N_VGND_M1081_d N_VGND_M1003_s N_VGND_M1007_s
+ N_VGND_M1010_s N_VGND_M1015_s N_VGND_M1031_s N_VGND_M1040_s N_VGND_M1047_s
+ N_VGND_M1052_s N_VGND_M1056_s N_VGND_M1058_s N_VGND_M1062_s N_VGND_M1068_s
+ N_VGND_M1072_s N_VGND_M1077_s N_VGND_M1079_s N_VGND_M1083_s VGND
+ N_VGND_c_2075_n N_VGND_c_2077_n N_VGND_c_2079_n N_VGND_c_2081_n
+ N_VGND_c_2083_n N_VGND_c_2085_n N_VGND_c_2087_n N_VGND_c_2089_n
+ N_VGND_c_2091_n N_VGND_c_2093_n N_VGND_c_2095_n N_VGND_c_2097_n
+ N_VGND_c_2099_n N_VGND_c_2101_n N_VGND_c_2103_n N_VGND_c_2105_n
+ N_VGND_c_2107_n N_VGND_c_2109_n N_VGND_c_2111_n N_VGND_c_2113_n
+ N_VGND_c_2115_n N_VGND_c_2117_n N_VGND_c_2119_n VGND
+ PM_SKY130_FD_SC_HVL__BUF_32%VGND
cc_1 N_VNB_M1008_b N_A_c_411_n 0.0468242f $X=-0.33 $Y=-0.265 $X2=0.665 $Y2=1.565
cc_2 N_VNB_c_2_p N_A_c_411_n 0.00104452f $X=33.36 $Y=0 $X2=0.665 $Y2=1.565
cc_3 N_VNB_M1008_b N_A_c_413_n 0.0390915f $X=-0.33 $Y=-0.265 $X2=1.445 $Y2=1.565
cc_4 N_VNB_c_2_p N_A_c_413_n 5.62728e-19 $X=33.36 $Y=0 $X2=1.445 $Y2=1.565
cc_5 N_VNB_M1008_b N_A_c_415_n 0.0405965f $X=-0.33 $Y=-0.265 $X2=2.225 $Y2=1.565
cc_6 N_VNB_c_2_p N_A_c_415_n 9.48159e-19 $X=33.36 $Y=0 $X2=2.225 $Y2=1.565
cc_7 N_VNB_M1008_b N_A_c_417_n 0.0400608f $X=-0.33 $Y=-0.265 $X2=3.005 $Y2=1.565
cc_8 N_VNB_c_2_p N_A_c_417_n 7.93986e-19 $X=33.36 $Y=0 $X2=3.005 $Y2=1.565
cc_9 N_VNB_M1008_b N_A_c_419_n 0.0397162f $X=-0.33 $Y=-0.265 $X2=3.785 $Y2=1.565
cc_10 N_VNB_c_2_p N_A_c_419_n 6.97629e-19 $X=33.36 $Y=0 $X2=3.785 $Y2=1.565
cc_11 N_VNB_M1008_b N_A_c_421_n 0.0382538f $X=-0.33 $Y=-0.265 $X2=4.565
+ $Y2=1.565
cc_12 N_VNB_c_2_p N_A_c_421_n 4.85642e-19 $X=33.36 $Y=0 $X2=4.565 $Y2=1.565
cc_13 N_VNB_M1008_b N_A_c_423_n 0.0399935f $X=-0.33 $Y=-0.265 $X2=5.345
+ $Y2=1.565
cc_14 N_VNB_c_2_p N_A_c_423_n 0.00102524f $X=33.36 $Y=0 $X2=5.345 $Y2=1.565
cc_15 N_VNB_M1008_b N_A_c_425_n 0.0390701f $X=-0.33 $Y=-0.265 $X2=6.125
+ $Y2=1.565
cc_16 N_VNB_c_2_p N_A_c_425_n 7.93986e-19 $X=33.36 $Y=0 $X2=6.125 $Y2=1.565
cc_17 N_VNB_M1008_b N_A_c_427_n 0.0387251f $X=-0.33 $Y=-0.265 $X2=6.905
+ $Y2=1.565
cc_18 N_VNB_c_2_p N_A_c_427_n 6.97629e-19 $X=33.36 $Y=0 $X2=6.905 $Y2=1.565
cc_19 N_VNB_M1008_b N_A_c_429_n 0.0406269f $X=-0.33 $Y=-0.265 $X2=7.685
+ $Y2=1.565
cc_20 N_VNB_c_2_p N_A_c_429_n 4.81788e-19 $X=33.36 $Y=0 $X2=7.685 $Y2=1.565
cc_21 N_VNB_M1008_b N_A_c_431_n 0.0094895f $X=-0.33 $Y=-0.265 $X2=4.465 $Y2=1.73
cc_22 N_VNB_M1008_b N_A_c_432_n 0.309862f $X=-0.33 $Y=-0.265 $X2=7.685 $Y2=1.815
cc_23 N_VNB_M1008_b N_A_183_141#_c_614_n 0.046867f $X=-0.33 $Y=-0.265 $X2=3.785
+ $Y2=1.08
cc_24 N_VNB_c_2_p N_A_183_141#_c_614_n 0.00183079f $X=33.36 $Y=0 $X2=3.785
+ $Y2=1.08
cc_25 N_VNB_M1008_b N_A_183_141#_c_616_n 0.039525f $X=-0.33 $Y=-0.265 $X2=4.565
+ $Y2=1.08
cc_26 N_VNB_c_2_p N_A_183_141#_c_616_n 7.55443e-19 $X=33.36 $Y=0 $X2=4.565
+ $Y2=1.08
cc_27 N_VNB_M1008_b N_A_183_141#_c_618_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=5.345
+ $Y2=1.08
cc_28 N_VNB_c_2_p N_A_183_141#_c_618_n 7.55443e-19 $X=33.36 $Y=0 $X2=5.345
+ $Y2=1.08
cc_29 N_VNB_M1008_b N_A_183_141#_c_620_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=6.125
+ $Y2=1.08
cc_30 N_VNB_c_2_p N_A_183_141#_c_620_n 7.55443e-19 $X=33.36 $Y=0 $X2=6.125
+ $Y2=1.08
cc_31 N_VNB_M1008_b N_A_183_141#_c_622_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=6.905
+ $Y2=1.08
cc_32 N_VNB_c_2_p N_A_183_141#_c_622_n 7.55443e-19 $X=33.36 $Y=0 $X2=6.905
+ $Y2=1.08
cc_33 N_VNB_M1008_b N_A_183_141#_c_624_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=7.685
+ $Y2=1.08
cc_34 N_VNB_c_2_p N_A_183_141#_c_624_n 7.55443e-19 $X=33.36 $Y=0 $X2=7.685
+ $Y2=1.08
cc_35 N_VNB_M1008_b N_A_183_141#_c_626_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=1.595
+ $Y2=1.58
cc_36 N_VNB_c_2_p N_A_183_141#_c_626_n 7.55443e-19 $X=33.36 $Y=0 $X2=1.595
+ $Y2=1.58
cc_37 N_VNB_M1008_b N_A_183_141#_c_628_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_38 N_VNB_c_2_p N_A_183_141#_c_628_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_39 N_VNB_M1008_b N_A_183_141#_c_630_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0.385
+ $Y2=1.73
cc_40 N_VNB_c_2_p N_A_183_141#_c_630_n 7.55443e-19 $X=33.36 $Y=0 $X2=0.385
+ $Y2=1.73
cc_41 N_VNB_M1008_b N_A_183_141#_c_632_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=4.465
+ $Y2=1.815
cc_42 N_VNB_c_2_p N_A_183_141#_c_632_n 7.55443e-19 $X=33.36 $Y=0 $X2=4.465
+ $Y2=1.815
cc_43 N_VNB_M1008_b N_A_183_141#_c_634_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=7.685
+ $Y2=1.815
cc_44 N_VNB_c_2_p N_A_183_141#_c_634_n 7.55443e-19 $X=33.36 $Y=0 $X2=7.685
+ $Y2=1.815
cc_45 N_VNB_M1008_b N_A_183_141#_c_636_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_c_2_p N_A_183_141#_c_636_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_47 N_VNB_M1008_b N_A_183_141#_c_638_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=3.12
+ $Y2=1.697
cc_48 N_VNB_c_2_p N_A_183_141#_c_638_n 7.55443e-19 $X=33.36 $Y=0 $X2=3.12
+ $Y2=1.697
cc_49 N_VNB_M1008_b N_A_183_141#_c_640_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_c_2_p N_A_183_141#_c_640_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_51 N_VNB_M1008_b N_A_183_141#_c_642_n 0.0395229f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_52 N_VNB_c_2_p N_A_183_141#_c_642_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_53 N_VNB_M1008_b N_A_183_141#_c_644_n 0.0410269f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_54 N_VNB_c_2_p N_A_183_141#_c_644_n 0.00106379f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_55 N_VNB_M1008_b N_A_183_141#_c_646_n 0.0448195f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_56 N_VNB_c_2_p N_A_183_141#_c_646_n 0.00183465f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_57 N_VNB_M1008_b N_A_183_141#_c_648_n 0.039525f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_58 N_VNB_c_2_p N_A_183_141#_c_648_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_59 N_VNB_M1008_b N_A_183_141#_c_650_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_60 N_VNB_c_2_p N_A_183_141#_c_650_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_61 N_VNB_M1008_b N_A_183_141#_c_652_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_62 N_VNB_c_2_p N_A_183_141#_c_652_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_63 N_VNB_M1008_b N_A_183_141#_c_654_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_64 N_VNB_c_2_p N_A_183_141#_c_654_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_65 N_VNB_M1008_b N_A_183_141#_c_656_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_66 N_VNB_c_2_p N_A_183_141#_c_656_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_67 N_VNB_M1008_b N_A_183_141#_c_658_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_68 N_VNB_c_2_p N_A_183_141#_c_658_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_69 N_VNB_M1008_b N_A_183_141#_c_660_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_70 N_VNB_c_2_p N_A_183_141#_c_660_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_71 N_VNB_M1008_b N_A_183_141#_c_662_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_72 N_VNB_c_2_p N_A_183_141#_c_662_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_73 N_VNB_M1008_b N_A_183_141#_c_664_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_74 N_VNB_c_2_p N_A_183_141#_c_664_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_75 N_VNB_M1008_b N_A_183_141#_c_666_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_76 N_VNB_c_2_p N_A_183_141#_c_666_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_77 N_VNB_M1008_b N_A_183_141#_c_668_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_78 N_VNB_c_2_p N_A_183_141#_c_668_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_79 N_VNB_M1008_b N_A_183_141#_c_670_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_80 N_VNB_c_2_p N_A_183_141#_c_670_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_81 N_VNB_M1008_b N_A_183_141#_c_672_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_82 N_VNB_c_2_p N_A_183_141#_c_672_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_83 N_VNB_M1008_b N_A_183_141#_c_674_n 0.0395229f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_84 N_VNB_c_2_p N_A_183_141#_c_674_n 7.55443e-19 $X=33.36 $Y=0 $X2=0 $Y2=0
cc_85 N_VNB_M1008_b N_A_183_141#_c_676_n 0.997928f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_86 N_VNB_c_2_p N_A_183_141#_c_676_n 0.00106379f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_87 N_VNB_M1008_b N_A_183_141#_c_678_n 0.00340102f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_88 N_VNB_M1008_b N_A_183_141#_c_679_n 0.00388959f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_89 N_VNB_M1008_b N_A_183_141#_c_680_n 0.00250789f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_90 N_VNB_M1008_b N_A_183_141#_c_681_n 0.00381091f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_91 N_VNB_M1008_b N_A_183_141#_c_682_n 0.00250789f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_92 N_VNB_M1008_b N_A_183_141#_c_683_n 0.00120049f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_93 N_VNB_M1008_b N_A_183_141#_c_684_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_94 N_VNB_M1008_b N_A_183_141#_c_685_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_95 N_VNB_M1008_b N_A_183_141#_c_686_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_96 N_VNB_M1008_b N_A_183_141#_c_687_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_97 N_VNB_M1008_b N_A_183_141#_c_688_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_98 N_VNB_M1008_b N_A_183_141#_c_689_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_99 N_VNB_M1008_b N_A_183_141#_c_690_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_100 N_VNB_M1008_b N_A_183_141#_c_691_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_101 N_VNB_M1008_b N_A_183_141#_c_692_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_102 N_VNB_M1008_b N_A_183_141#_c_693_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_103 N_VNB_M1008_b N_A_183_141#_c_694_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_104 N_VNB_M1008_b N_A_183_141#_c_695_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_105 N_VNB_M1008_b N_A_183_141#_c_696_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_106 N_VNB_M1008_b N_A_183_141#_c_697_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_107 N_VNB_M1008_b N_A_183_141#_c_698_n 0.040604f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_108 N_VNB_M1008_b N_A_183_141#_c_699_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_109 N_VNB_M1008_b N_VGND_c_2075_n 0.0613833f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_110 N_VNB_c_2_p N_VGND_c_2075_n 0.00138265f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_111 N_VNB_M1008_b N_VGND_c_2077_n 0.0415829f $X=-0.33 $Y=-0.265 $X2=3.515
+ $Y2=1.58
cc_112 N_VNB_c_2_p N_VGND_c_2077_n 0.00234213f $X=33.36 $Y=0 $X2=3.515 $Y2=1.58
cc_113 N_VNB_M1008_b N_VGND_c_2079_n 0.0399392f $X=-0.33 $Y=-0.265 $X2=0.385
+ $Y2=1.73
cc_114 N_VNB_c_2_p N_VGND_c_2079_n 0.0023214f $X=33.36 $Y=0 $X2=0.385 $Y2=1.73
cc_115 N_VNB_M1008_b N_VGND_c_2081_n 0.0397337f $X=-0.33 $Y=-0.265 $X2=4.465
+ $Y2=1.73
cc_116 N_VNB_c_2_p N_VGND_c_2081_n 0.00230841f $X=33.36 $Y=0 $X2=4.465 $Y2=1.73
cc_117 N_VNB_M1008_b N_VGND_c_2083_n 0.039938f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_118 N_VNB_c_2_p N_VGND_c_2083_n 0.0023214f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_119 N_VNB_M1008_b N_VGND_c_2085_n 0.039901f $X=-0.33 $Y=-0.265 $X2=2.64
+ $Y2=1.697
cc_120 N_VNB_c_2_p N_VGND_c_2085_n 0.00230355f $X=33.36 $Y=0 $X2=2.64 $Y2=1.697
cc_121 N_VNB_M1008_b N_VGND_c_2087_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_122 N_VNB_c_2_p N_VGND_c_2087_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_123 N_VNB_M1008_b N_VGND_c_2089_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_124 N_VNB_c_2_p N_VGND_c_2089_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_125 N_VNB_M1008_b N_VGND_c_2091_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_126 N_VNB_c_2_p N_VGND_c_2091_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_127 N_VNB_M1008_b N_VGND_c_2093_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_128 N_VNB_c_2_p N_VGND_c_2093_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_129 N_VNB_M1008_b N_VGND_c_2095_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_130 N_VNB_c_2_p N_VGND_c_2095_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_131 N_VNB_M1008_b N_VGND_c_2097_n 0.039901f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_132 N_VNB_c_2_p N_VGND_c_2097_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_133 N_VNB_M1008_b N_VGND_c_2099_n 0.0256175f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_134 N_VNB_c_2_p N_VGND_c_2099_n 0.00136968f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_135 N_VNB_M1008_b N_VGND_c_2101_n 0.039901f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_136 N_VNB_c_2_p N_VGND_c_2101_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_137 N_VNB_M1008_b N_VGND_c_2103_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_138 N_VNB_c_2_p N_VGND_c_2103_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_139 N_VNB_M1008_b N_VGND_c_2105_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_140 N_VNB_c_2_p N_VGND_c_2105_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_141 N_VNB_M1008_b N_VGND_c_2107_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_142 N_VNB_c_2_p N_VGND_c_2107_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_143 N_VNB_M1008_b N_VGND_c_2109_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_144 N_VNB_c_2_p N_VGND_c_2109_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_145 N_VNB_M1008_b N_VGND_c_2111_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_146 N_VNB_c_2_p N_VGND_c_2111_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_147 N_VNB_M1008_b N_VGND_c_2113_n 0.039901f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_148 N_VNB_c_2_p N_VGND_c_2113_n 0.00230355f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_149 N_VNB_M1008_b N_VGND_c_2115_n 0.0684821f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_150 N_VNB_c_2_p N_VGND_c_2115_n 0.00136968f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_151 N_VNB_M1008_b N_VGND_c_2117_n 0.466f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_152 N_VNB_c_2_p N_VGND_c_2117_n 3.59503f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_153 N_VNB_M1008_b N_VGND_c_2119_n 0.042773f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_154 N_VNB_c_2_p N_VGND_c_2119_n 0.00238667f $X=33.36 $Y=0 $X2=0 $Y2=0
cc_155 N_VPB_M1000_b N_A_M1000_g 0.0430944f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=2.965
cc_156 N_VPB_c_156_p N_A_M1000_g 0.0157621f $X=33.36 $Y=4.07 $X2=0.665 $Y2=2.965
cc_157 N_VPB_c_157_p N_A_M1000_g 0.00970178f $X=33.36 $Y=4.07 $X2=0.665
+ $Y2=2.965
cc_158 N_VPB_M1000_b N_A_M1001_g 0.0352958f $X=-0.33 $Y=1.885 $X2=1.445
+ $Y2=2.965
cc_159 N_VPB_c_156_p N_A_M1001_g 0.0157169f $X=33.36 $Y=4.07 $X2=1.445 $Y2=2.965
cc_160 N_VPB_c_157_p N_A_M1001_g 0.00970178f $X=33.36 $Y=4.07 $X2=1.445
+ $Y2=2.965
cc_161 N_VPB_M1000_b N_A_M1006_g 0.0352691f $X=-0.33 $Y=1.885 $X2=2.225
+ $Y2=2.965
cc_162 N_VPB_c_156_p N_A_M1006_g 0.0159522f $X=33.36 $Y=4.07 $X2=2.225 $Y2=2.965
cc_163 N_VPB_c_157_p N_A_M1006_g 0.00970178f $X=33.36 $Y=4.07 $X2=2.225
+ $Y2=2.965
cc_164 N_VPB_M1000_b N_A_M1016_g 0.0352958f $X=-0.33 $Y=1.885 $X2=3.005
+ $Y2=2.965
cc_165 N_VPB_c_156_p N_A_M1016_g 0.0154933f $X=33.36 $Y=4.07 $X2=3.005 $Y2=2.965
cc_166 N_VPB_c_157_p N_A_M1016_g 0.00970178f $X=33.36 $Y=4.07 $X2=3.005
+ $Y2=2.965
cc_167 N_VPB_M1000_b N_A_M1019_g 0.0352669f $X=-0.33 $Y=1.885 $X2=3.785
+ $Y2=2.965
cc_168 N_VPB_c_156_p N_A_M1019_g 0.0159373f $X=33.36 $Y=4.07 $X2=3.785 $Y2=2.965
cc_169 N_VPB_c_157_p N_A_M1019_g 0.00970178f $X=33.36 $Y=4.07 $X2=3.785
+ $Y2=2.965
cc_170 N_VPB_M1000_b N_A_M1035_g 0.0352958f $X=-0.33 $Y=1.885 $X2=4.565
+ $Y2=2.965
cc_171 N_VPB_c_156_p N_A_M1035_g 0.0157169f $X=33.36 $Y=4.07 $X2=4.565 $Y2=2.965
cc_172 N_VPB_c_157_p N_A_M1035_g 0.00970178f $X=33.36 $Y=4.07 $X2=4.565
+ $Y2=2.965
cc_173 N_VPB_M1000_b N_A_M1039_g 0.0352691f $X=-0.33 $Y=1.885 $X2=5.345
+ $Y2=2.965
cc_174 N_VPB_c_156_p N_A_M1039_g 0.0159522f $X=33.36 $Y=4.07 $X2=5.345 $Y2=2.965
cc_175 N_VPB_c_157_p N_A_M1039_g 0.00970178f $X=33.36 $Y=4.07 $X2=5.345
+ $Y2=2.965
cc_176 N_VPB_M1000_b N_A_M1049_g 0.0352958f $X=-0.33 $Y=1.885 $X2=6.125
+ $Y2=2.965
cc_177 N_VPB_c_156_p N_A_M1049_g 0.0154933f $X=33.36 $Y=4.07 $X2=6.125 $Y2=2.965
cc_178 N_VPB_c_157_p N_A_M1049_g 0.00970178f $X=33.36 $Y=4.07 $X2=6.125
+ $Y2=2.965
cc_179 N_VPB_M1000_b N_A_M1064_g 0.0352669f $X=-0.33 $Y=1.885 $X2=6.905
+ $Y2=2.965
cc_180 N_VPB_c_156_p N_A_M1064_g 0.0159373f $X=33.36 $Y=4.07 $X2=6.905 $Y2=2.965
cc_181 N_VPB_c_157_p N_A_M1064_g 0.00970178f $X=33.36 $Y=4.07 $X2=6.905
+ $Y2=2.965
cc_182 N_VPB_M1000_b N_A_M1070_g 0.0392745f $X=-0.33 $Y=1.885 $X2=7.685
+ $Y2=2.965
cc_183 N_VPB_c_156_p N_A_M1070_g 0.0157169f $X=33.36 $Y=4.07 $X2=7.685 $Y2=2.965
cc_184 N_VPB_c_157_p N_A_M1070_g 0.00970178f $X=33.36 $Y=4.07 $X2=7.685
+ $Y2=2.965
cc_185 N_VPB_M1000_b N_A_c_432_n 0.192917f $X=-0.33 $Y=1.885 $X2=7.685 $Y2=1.815
cc_186 N_VPB_M1000_b N_A_183_141#_M1004_g 0.0443277f $X=-0.33 $Y=1.885 $X2=4.565
+ $Y2=1.565
cc_187 N_VPB_c_156_p N_A_183_141#_M1004_g 0.0191204f $X=33.36 $Y=4.07 $X2=4.565
+ $Y2=1.565
cc_188 N_VPB_c_157_p N_A_183_141#_M1004_g 0.00970178f $X=33.36 $Y=4.07 $X2=4.565
+ $Y2=1.565
cc_189 N_VPB_M1000_b N_A_183_141#_M1011_g 0.040726f $X=-0.33 $Y=1.885 $X2=5.345
+ $Y2=1.565
cc_190 N_VPB_c_156_p N_A_183_141#_M1011_g 0.0157621f $X=33.36 $Y=4.07 $X2=5.345
+ $Y2=1.565
cc_191 N_VPB_c_157_p N_A_183_141#_M1011_g 0.00970178f $X=33.36 $Y=4.07 $X2=5.345
+ $Y2=1.565
cc_192 N_VPB_M1000_b N_A_183_141#_M1013_g 0.040726f $X=-0.33 $Y=1.885 $X2=6.125
+ $Y2=1.565
cc_193 N_VPB_c_156_p N_A_183_141#_M1013_g 0.0157621f $X=33.36 $Y=4.07 $X2=6.125
+ $Y2=1.565
cc_194 N_VPB_c_157_p N_A_183_141#_M1013_g 0.00970178f $X=33.36 $Y=4.07 $X2=6.125
+ $Y2=1.565
cc_195 N_VPB_M1000_b N_A_183_141#_M1017_g 0.040726f $X=-0.33 $Y=1.885 $X2=6.905
+ $Y2=1.565
cc_196 N_VPB_c_156_p N_A_183_141#_M1017_g 0.0157621f $X=33.36 $Y=4.07 $X2=6.905
+ $Y2=1.565
cc_197 N_VPB_c_157_p N_A_183_141#_M1017_g 0.00970178f $X=33.36 $Y=4.07 $X2=6.905
+ $Y2=1.565
cc_198 N_VPB_M1000_b N_A_183_141#_M1018_g 0.040726f $X=-0.33 $Y=1.885 $X2=7.685
+ $Y2=1.565
cc_199 N_VPB_c_156_p N_A_183_141#_M1018_g 0.0157621f $X=33.36 $Y=4.07 $X2=7.685
+ $Y2=1.565
cc_200 N_VPB_c_157_p N_A_183_141#_M1018_g 0.00970178f $X=33.36 $Y=4.07 $X2=7.685
+ $Y2=1.565
cc_201 N_VPB_M1000_b N_A_183_141#_M1020_g 0.040726f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_202 N_VPB_c_156_p N_A_183_141#_M1020_g 0.0157621f $X=33.36 $Y=4.07 $X2=0.635
+ $Y2=1.58
cc_203 N_VPB_c_157_p N_A_183_141#_M1020_g 0.00970178f $X=33.36 $Y=4.07 $X2=0.635
+ $Y2=1.58
cc_204 N_VPB_M1000_b N_A_183_141#_M1021_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_205 N_VPB_c_156_p N_A_183_141#_M1021_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_206 N_VPB_c_157_p N_A_183_141#_M1021_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_207 N_VPB_M1000_b N_A_183_141#_M1022_g 0.040726f $X=-0.33 $Y=1.885 $X2=0.385
+ $Y2=1.815
cc_208 N_VPB_c_156_p N_A_183_141#_M1022_g 0.0157621f $X=33.36 $Y=4.07 $X2=0.385
+ $Y2=1.815
cc_209 N_VPB_c_157_p N_A_183_141#_M1022_g 0.00970178f $X=33.36 $Y=4.07 $X2=0.385
+ $Y2=1.815
cc_210 N_VPB_M1000_b N_A_183_141#_M1023_g 0.040726f $X=-0.33 $Y=1.885 $X2=3.005
+ $Y2=1.815
cc_211 N_VPB_c_156_p N_A_183_141#_M1023_g 0.0157621f $X=33.36 $Y=4.07 $X2=3.005
+ $Y2=1.815
cc_212 N_VPB_c_157_p N_A_183_141#_M1023_g 0.00970178f $X=33.36 $Y=4.07 $X2=3.005
+ $Y2=1.815
cc_213 N_VPB_M1000_b N_A_183_141#_M1024_g 0.040726f $X=-0.33 $Y=1.885 $X2=6.125
+ $Y2=1.815
cc_214 N_VPB_c_156_p N_A_183_141#_M1024_g 0.0157621f $X=33.36 $Y=4.07 $X2=6.125
+ $Y2=1.815
cc_215 N_VPB_c_157_p N_A_183_141#_M1024_g 0.00970178f $X=33.36 $Y=4.07 $X2=6.125
+ $Y2=1.815
cc_216 N_VPB_M1000_b N_A_183_141#_M1026_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_217 N_VPB_c_156_p N_A_183_141#_M1026_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_218 N_VPB_c_157_p N_A_183_141#_M1026_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_219 N_VPB_M1000_b N_A_183_141#_M1029_g 0.040726f $X=-0.33 $Y=1.885 $X2=2.64
+ $Y2=1.697
cc_220 N_VPB_c_156_p N_A_183_141#_M1029_g 0.0157621f $X=33.36 $Y=4.07 $X2=2.64
+ $Y2=1.697
cc_221 N_VPB_c_157_p N_A_183_141#_M1029_g 0.00970178f $X=33.36 $Y=4.07 $X2=2.64
+ $Y2=1.697
cc_222 N_VPB_M1000_b N_A_183_141#_M1030_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_223 N_VPB_c_156_p N_A_183_141#_M1030_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_224 N_VPB_c_157_p N_A_183_141#_M1030_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_225 N_VPB_M1000_b N_A_183_141#_M1033_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_226 N_VPB_c_156_p N_A_183_141#_M1033_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_227 N_VPB_c_157_p N_A_183_141#_M1033_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_228 N_VPB_M1000_b N_A_183_141#_M1034_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_229 N_VPB_c_156_p N_A_183_141#_M1034_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_230 N_VPB_c_157_p N_A_183_141#_M1034_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_231 N_VPB_M1000_b N_A_183_141#_M1036_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_232 N_VPB_c_156_p N_A_183_141#_M1036_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_233 N_VPB_c_157_p N_A_183_141#_M1036_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_234 N_VPB_M1000_b N_A_183_141#_M1037_g 0.0407837f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_235 N_VPB_c_156_p N_A_183_141#_M1037_g 0.0191024f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_236 N_VPB_c_157_p N_A_183_141#_M1037_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_237 N_VPB_M1000_b N_A_183_141#_M1041_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_238 N_VPB_c_156_p N_A_183_141#_M1041_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_239 N_VPB_c_157_p N_A_183_141#_M1041_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_240 N_VPB_M1000_b N_A_183_141#_M1042_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_241 N_VPB_c_156_p N_A_183_141#_M1042_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_242 N_VPB_c_157_p N_A_183_141#_M1042_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_243 N_VPB_M1000_b N_A_183_141#_M1045_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_244 N_VPB_c_156_p N_A_183_141#_M1045_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_245 N_VPB_c_157_p N_A_183_141#_M1045_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_246 N_VPB_M1000_b N_A_183_141#_M1046_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_247 N_VPB_c_156_p N_A_183_141#_M1046_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_248 N_VPB_c_157_p N_A_183_141#_M1046_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_249 N_VPB_M1000_b N_A_183_141#_M1050_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_250 N_VPB_c_156_p N_A_183_141#_M1050_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_251 N_VPB_c_157_p N_A_183_141#_M1050_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_252 N_VPB_M1000_b N_A_183_141#_M1054_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_253 N_VPB_c_156_p N_A_183_141#_M1054_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_254 N_VPB_c_157_p N_A_183_141#_M1054_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_255 N_VPB_M1000_b N_A_183_141#_M1055_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_256 N_VPB_c_156_p N_A_183_141#_M1055_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_257 N_VPB_c_157_p N_A_183_141#_M1055_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_258 N_VPB_M1000_b N_A_183_141#_M1059_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_259 N_VPB_c_156_p N_A_183_141#_M1059_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_260 N_VPB_c_157_p N_A_183_141#_M1059_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_261 N_VPB_M1000_b N_A_183_141#_M1060_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_262 N_VPB_c_156_p N_A_183_141#_M1060_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_263 N_VPB_c_157_p N_A_183_141#_M1060_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_264 N_VPB_M1000_b N_A_183_141#_M1063_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_265 N_VPB_c_156_p N_A_183_141#_M1063_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_266 N_VPB_c_157_p N_A_183_141#_M1063_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_267 N_VPB_M1000_b N_A_183_141#_M1065_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_268 N_VPB_c_156_p N_A_183_141#_M1065_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_269 N_VPB_c_157_p N_A_183_141#_M1065_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_270 N_VPB_M1000_b N_A_183_141#_M1066_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_271 N_VPB_c_156_p N_A_183_141#_M1066_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_272 N_VPB_c_157_p N_A_183_141#_M1066_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_273 N_VPB_M1000_b N_A_183_141#_M1073_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_274 N_VPB_c_156_p N_A_183_141#_M1073_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_275 N_VPB_c_157_p N_A_183_141#_M1073_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_276 N_VPB_M1000_b N_A_183_141#_M1075_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_277 N_VPB_c_156_p N_A_183_141#_M1075_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_278 N_VPB_c_157_p N_A_183_141#_M1075_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_279 N_VPB_M1000_b N_A_183_141#_c_676_n 0.407373f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_280 N_VPB_M1000_b N_A_183_141#_M1080_g 0.0502706f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_281 N_VPB_c_156_p N_A_183_141#_M1080_g 0.0157621f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_282 N_VPB_c_157_p N_A_183_141#_M1080_g 0.00970178f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_283 N_VPB_M1000_b N_A_183_141#_c_797_n 0.00168525f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_284 N_VPB_c_156_p N_A_183_141#_c_797_n 0.0160222f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_285 N_VPB_c_157_p N_A_183_141#_c_797_n 0.00105499f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_286 N_VPB_M1000_b N_A_183_141#_c_800_n 0.00161463f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_287 N_VPB_c_156_p N_A_183_141#_c_800_n 0.0159826f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_288 N_VPB_c_157_p N_A_183_141#_c_800_n 0.00107233f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_289 N_VPB_M1000_b N_A_183_141#_c_803_n 0.00173328f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_290 N_VPB_c_156_p N_A_183_141#_c_803_n 0.0180171f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_291 N_VPB_c_157_p N_A_183_141#_c_803_n 0.00122962f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_292 N_VPB_M1000_b N_A_183_141#_c_806_n 0.00161463f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_293 N_VPB_c_156_p N_A_183_141#_c_806_n 0.0159826f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_294 N_VPB_c_157_p N_A_183_141#_c_806_n 0.00107233f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_295 N_VPB_M1000_b N_A_183_141#_c_809_n 0.00173328f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_296 N_VPB_c_156_p N_A_183_141#_c_809_n 0.0180171f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_297 N_VPB_c_157_p N_A_183_141#_c_809_n 0.00122962f $X=33.36 $Y=4.07 $X2=0
+ $Y2=0
cc_298 N_VPB_M1000_b N_A_183_141#_c_683_n 0.00159506f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_299 N_VPB_M1000_b N_VPWR_c_1410_n 0.0644578f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_300 N_VPB_c_156_p N_VPWR_c_1410_n 0.0289697f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_301 N_VPB_c_157_p N_VPWR_c_1410_n 0.00219871f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_302 N_VPB_c_156_p N_VPWR_c_1413_n 0.0306445f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_303 N_VPB_c_157_p N_VPWR_c_1413_n 0.00361083f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_304 N_VPB_c_156_p N_VPWR_c_1415_n 0.0306445f $X=33.36 $Y=4.07 $X2=1.445
+ $Y2=1.815
cc_305 N_VPB_c_157_p N_VPWR_c_1415_n 0.00361083f $X=33.36 $Y=4.07 $X2=1.445
+ $Y2=1.815
cc_306 N_VPB_c_156_p N_VPWR_c_1417_n 0.0306445f $X=33.36 $Y=4.07 $X2=7.685
+ $Y2=1.815
cc_307 N_VPB_c_157_p N_VPWR_c_1417_n 0.00361083f $X=33.36 $Y=4.07 $X2=7.685
+ $Y2=1.815
cc_308 N_VPB_c_156_p N_VPWR_c_1419_n 0.0306445f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_309 N_VPB_c_157_p N_VPWR_c_1419_n 0.00361083f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_310 N_VPB_c_156_p N_VPWR_c_1421_n 0.0315613f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_311 N_VPB_c_157_p N_VPWR_c_1421_n 0.00318367f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_312 N_VPB_M1000_b N_VPWR_c_1423_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_313 N_VPB_c_156_p N_VPWR_c_1423_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_314 N_VPB_c_157_p N_VPWR_c_1423_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_315 N_VPB_M1000_b N_VPWR_c_1426_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_316 N_VPB_c_156_p N_VPWR_c_1426_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_317 N_VPB_c_157_p N_VPWR_c_1426_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_318 N_VPB_M1000_b N_VPWR_c_1429_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_319 N_VPB_c_156_p N_VPWR_c_1429_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_320 N_VPB_c_157_p N_VPWR_c_1429_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_321 N_VPB_M1000_b N_VPWR_c_1432_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_322 N_VPB_c_156_p N_VPWR_c_1432_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_323 N_VPB_c_157_p N_VPWR_c_1432_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_324 N_VPB_M1000_b N_VPWR_c_1435_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_325 N_VPB_c_156_p N_VPWR_c_1435_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_326 N_VPB_c_157_p N_VPWR_c_1435_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_327 N_VPB_M1000_b N_VPWR_c_1438_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_328 N_VPB_c_156_p N_VPWR_c_1438_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_329 N_VPB_c_157_p N_VPWR_c_1438_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_330 N_VPB_M1000_b N_VPWR_c_1441_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_331 N_VPB_c_156_p N_VPWR_c_1441_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_332 N_VPB_c_157_p N_VPWR_c_1441_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_333 N_VPB_M1000_b N_VPWR_c_1444_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_334 N_VPB_c_156_p N_VPWR_c_1444_n 0.0269193f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_335 N_VPB_c_157_p N_VPWR_c_1444_n 0.00204836f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_336 N_VPB_M1000_b N_VPWR_c_1447_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_337 N_VPB_c_156_p N_VPWR_c_1447_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_338 N_VPB_c_157_p N_VPWR_c_1447_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_339 N_VPB_M1000_b N_VPWR_c_1450_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_340 N_VPB_c_156_p N_VPWR_c_1450_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_341 N_VPB_c_157_p N_VPWR_c_1450_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_342 N_VPB_M1000_b N_VPWR_c_1453_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_343 N_VPB_c_156_p N_VPWR_c_1453_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_344 N_VPB_c_157_p N_VPWR_c_1453_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_345 N_VPB_M1000_b N_VPWR_c_1456_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_346 N_VPB_c_156_p N_VPWR_c_1456_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_347 N_VPB_c_157_p N_VPWR_c_1456_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_348 N_VPB_M1000_b N_VPWR_c_1459_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_349 N_VPB_c_156_p N_VPWR_c_1459_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_350 N_VPB_c_157_p N_VPWR_c_1459_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_351 N_VPB_M1000_b N_VPWR_c_1462_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_352 N_VPB_c_156_p N_VPWR_c_1462_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_353 N_VPB_c_157_p N_VPWR_c_1462_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_354 N_VPB_M1000_b N_VPWR_c_1465_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_355 N_VPB_c_156_p N_VPWR_c_1465_n 0.0445179f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_356 N_VPB_c_157_p N_VPWR_c_1465_n 0.00377602f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_357 N_VPB_M1000_b N_VPWR_c_1468_n 0.0633596f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_358 N_VPB_c_156_p N_VPWR_c_1468_n 0.0270143f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_359 N_VPB_c_157_p N_VPWR_c_1468_n 0.00200674f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_360 N_VPB_M1000_b N_VPWR_c_1471_n 0.0851249f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_361 N_VPB_c_156_p N_VPWR_c_1471_n 0.146635f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_362 N_VPB_c_157_p N_VPWR_c_1471_n 3.55827f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_363 N_VPB_M1000_b N_X_c_1741_n 0.00125033f $X=-0.33 $Y=1.885 $X2=6.905
+ $Y2=1.815
cc_364 N_VPB_c_156_p N_X_c_1741_n 0.0171423f $X=33.36 $Y=4.07 $X2=6.905
+ $Y2=1.815
cc_365 N_VPB_c_157_p N_X_c_1741_n 0.00108855f $X=33.36 $Y=4.07 $X2=6.905
+ $Y2=1.815
cc_366 N_VPB_M1000_b N_X_c_1744_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_367 N_VPB_c_156_p N_X_c_1744_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_368 N_VPB_c_157_p N_X_c_1744_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_369 N_VPB_M1000_b N_X_c_1747_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_370 N_VPB_c_156_p N_X_c_1747_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_371 N_VPB_c_157_p N_X_c_1747_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_372 N_VPB_M1000_b N_X_c_1750_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_373 N_VPB_c_156_p N_X_c_1750_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_374 N_VPB_c_157_p N_X_c_1750_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_375 N_VPB_M1000_b N_X_c_1753_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_376 N_VPB_c_156_p N_X_c_1753_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_377 N_VPB_c_157_p N_X_c_1753_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_378 N_VPB_M1000_b N_X_c_1756_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_379 N_VPB_c_156_p N_X_c_1756_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_380 N_VPB_c_157_p N_X_c_1756_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_381 N_VPB_M1000_b N_X_c_1759_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_382 N_VPB_c_156_p N_X_c_1759_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_383 N_VPB_c_157_p N_X_c_1759_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_384 N_VPB_M1000_b N_X_c_1762_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_385 N_VPB_c_156_p N_X_c_1762_n 0.0210531f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_386 N_VPB_c_157_p N_X_c_1762_n 0.00147247f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_387 N_VPB_M1000_b N_X_c_1765_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_388 N_VPB_c_156_p N_X_c_1765_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_389 N_VPB_c_157_p N_X_c_1765_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_390 N_VPB_M1000_b N_X_c_1768_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_391 N_VPB_c_156_p N_X_c_1768_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_392 N_VPB_c_157_p N_X_c_1768_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_393 N_VPB_M1000_b N_X_c_1771_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_394 N_VPB_c_156_p N_X_c_1771_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_395 N_VPB_c_157_p N_X_c_1771_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_396 N_VPB_M1000_b N_X_c_1774_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_397 N_VPB_c_156_p N_X_c_1774_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_398 N_VPB_c_157_p N_X_c_1774_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_399 N_VPB_M1000_b N_X_c_1777_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_400 N_VPB_c_156_p N_X_c_1777_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_401 N_VPB_c_157_p N_X_c_1777_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_402 N_VPB_M1000_b N_X_c_1780_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_403 N_VPB_c_156_p N_X_c_1780_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_404 N_VPB_c_157_p N_X_c_1780_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_405 N_VPB_M1000_b N_X_c_1783_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_406 N_VPB_c_156_p N_X_c_1783_n 0.0171423f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_407 N_VPB_c_157_p N_X_c_1783_n 0.00108855f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_408 N_VPB_M1000_b N_X_c_1786_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_409 N_VPB_c_156_p N_X_c_1786_n 0.0210531f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_410 N_VPB_c_157_p N_X_c_1786_n 0.00147247f $X=33.36 $Y=4.07 $X2=0 $Y2=0
cc_411 N_A_c_429_n N_A_183_141#_c_614_n 0.0172878f $X=7.685 $Y=1.565 $X2=0 $Y2=0
cc_412 N_A_M1070_g N_A_183_141#_M1004_g 0.0172878f $X=7.685 $Y=2.965 $X2=0 $Y2=0
cc_413 N_A_c_432_n N_A_183_141#_c_676_n 0.0172878f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_414 N_A_c_411_n N_A_183_141#_c_678_n 0.012066f $X=0.665 $Y=1.565 $X2=0 $Y2=0
cc_415 N_A_M1000_g N_A_183_141#_c_797_n 0.0293976f $X=0.665 $Y=2.965 $X2=0 $Y2=0
cc_416 N_A_M1001_g N_A_183_141#_c_797_n 0.0022192f $X=1.445 $Y=2.965 $X2=0 $Y2=0
cc_417 N_A_M1001_g N_A_183_141#_c_819_n 0.0253301f $X=1.445 $Y=2.965 $X2=0 $Y2=0
cc_418 N_A_M1006_g N_A_183_141#_c_819_n 0.0218849f $X=2.225 $Y=2.965 $X2=0 $Y2=0
cc_419 N_A_c_431_n N_A_183_141#_c_819_n 0.0894665f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_420 N_A_c_432_n N_A_183_141#_c_819_n 0.0283643f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_421 N_A_M1000_g N_A_183_141#_c_823_n 0.00954688f $X=0.665 $Y=2.965 $X2=0
+ $Y2=0
cc_422 N_A_c_431_n N_A_183_141#_c_823_n 0.024153f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_423 N_A_c_432_n N_A_183_141#_c_823_n 0.013297f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_424 N_A_c_413_n N_A_183_141#_c_826_n 0.0276926f $X=1.445 $Y=1.565 $X2=0 $Y2=0
cc_425 N_A_c_415_n N_A_183_141#_c_826_n 0.0243589f $X=2.225 $Y=1.565 $X2=0 $Y2=0
cc_426 N_A_c_431_n N_A_183_141#_c_826_n 0.0824875f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_427 N_A_c_432_n N_A_183_141#_c_826_n 0.0024988f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_428 N_A_c_411_n N_A_183_141#_c_830_n 0.00653924f $X=0.665 $Y=1.565 $X2=0
+ $Y2=0
cc_429 N_A_c_431_n N_A_183_141#_c_830_n 0.0242608f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_430 N_A_c_432_n N_A_183_141#_c_830_n 0.0025699f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_431 N_A_c_415_n N_A_183_141#_c_679_n 0.0163015f $X=2.225 $Y=1.565 $X2=0 $Y2=0
cc_432 N_A_c_417_n N_A_183_141#_c_679_n 0.0139077f $X=3.005 $Y=1.565 $X2=0 $Y2=0
cc_433 N_A_M1006_g N_A_183_141#_c_800_n 0.0373895f $X=2.225 $Y=2.965 $X2=0 $Y2=0
cc_434 N_A_M1016_g N_A_183_141#_c_800_n 0.00215741f $X=3.005 $Y=2.965 $X2=0
+ $Y2=0
cc_435 N_A_M1016_g N_A_183_141#_c_837_n 0.0246803f $X=3.005 $Y=2.965 $X2=0 $Y2=0
cc_436 N_A_M1019_g N_A_183_141#_c_837_n 0.0212247f $X=3.785 $Y=2.965 $X2=0 $Y2=0
cc_437 N_A_c_431_n N_A_183_141#_c_837_n 0.0887444f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_438 N_A_c_432_n N_A_183_141#_c_837_n 0.02815f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_439 N_A_c_417_n N_A_183_141#_c_841_n 0.026264f $X=3.005 $Y=1.565 $X2=0 $Y2=0
cc_440 N_A_c_419_n N_A_183_141#_c_841_n 0.0274546f $X=3.785 $Y=1.565 $X2=0 $Y2=0
cc_441 N_A_c_431_n N_A_183_141#_c_841_n 0.0837197f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_442 N_A_c_432_n N_A_183_141#_c_841_n 0.0024988f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_443 N_A_M1016_g N_A_183_141#_c_803_n 8.05117e-19 $X=3.005 $Y=2.965 $X2=0
+ $Y2=0
cc_444 N_A_M1019_g N_A_183_141#_c_803_n 0.0361085f $X=3.785 $Y=2.965 $X2=0 $Y2=0
cc_445 N_A_M1035_g N_A_183_141#_c_803_n 0.00227089f $X=4.565 $Y=2.965 $X2=0
+ $Y2=0
cc_446 N_A_c_419_n N_A_183_141#_c_680_n 0.0119333f $X=3.785 $Y=1.565 $X2=0 $Y2=0
cc_447 N_A_c_421_n N_A_183_141#_c_849_n 0.0262613f $X=4.565 $Y=1.565 $X2=0 $Y2=0
cc_448 N_A_c_431_n N_A_183_141#_c_849_n 0.0238559f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_449 N_A_M1035_g N_A_183_141#_c_851_n 0.022437f $X=4.565 $Y=2.965 $X2=0 $Y2=0
cc_450 N_A_c_431_n N_A_183_141#_c_851_n 0.0245146f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_451 N_A_c_432_n N_A_183_141#_c_851_n 0.0129239f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_452 N_A_c_423_n N_A_183_141#_c_681_n 0.0168315f $X=5.345 $Y=1.565 $X2=0 $Y2=0
cc_453 N_A_c_425_n N_A_183_141#_c_681_n 0.0140598f $X=6.125 $Y=1.565 $X2=0 $Y2=0
cc_454 N_A_c_432_n N_A_183_141#_c_681_n 2.89984e-19 $X=7.685 $Y=1.815 $X2=0
+ $Y2=0
cc_455 N_A_M1039_g N_A_183_141#_c_806_n 0.0376701f $X=5.345 $Y=2.965 $X2=0 $Y2=0
cc_456 N_A_M1049_g N_A_183_141#_c_806_n 0.00215741f $X=6.125 $Y=2.965 $X2=0
+ $Y2=0
cc_457 N_A_c_432_n N_A_183_141#_c_806_n 4.40368e-19 $X=7.685 $Y=1.815 $X2=0
+ $Y2=0
cc_458 N_A_c_425_n N_A_183_141#_c_860_n 0.0292193f $X=6.125 $Y=1.565 $X2=0 $Y2=0
cc_459 N_A_M1049_g N_A_183_141#_c_860_n 0.021273f $X=6.125 $Y=2.965 $X2=0 $Y2=0
cc_460 N_A_c_427_n N_A_183_141#_c_860_n 0.0252525f $X=6.905 $Y=1.565 $X2=0 $Y2=0
cc_461 N_A_M1064_g N_A_183_141#_c_860_n 0.0222171f $X=6.905 $Y=2.965 $X2=0 $Y2=0
cc_462 N_A_c_432_n N_A_183_141#_c_860_n 0.0579974f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_463 N_A_c_421_n N_A_183_141#_c_865_n 0.010257f $X=4.565 $Y=1.565 $X2=0 $Y2=0
cc_464 N_A_M1035_g N_A_183_141#_c_865_n 0.00288127f $X=4.565 $Y=2.965 $X2=0
+ $Y2=0
cc_465 N_A_c_423_n N_A_183_141#_c_865_n 0.0322234f $X=5.345 $Y=1.565 $X2=0 $Y2=0
cc_466 N_A_M1039_g N_A_183_141#_c_865_n 0.0264151f $X=5.345 $Y=2.965 $X2=0 $Y2=0
cc_467 N_A_c_425_n N_A_183_141#_c_865_n 0.00299493f $X=6.125 $Y=1.565 $X2=0
+ $Y2=0
cc_468 N_A_M1049_g N_A_183_141#_c_865_n 0.00418078f $X=6.125 $Y=2.965 $X2=0
+ $Y2=0
cc_469 N_A_c_431_n N_A_183_141#_c_865_n 0.0186888f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_470 N_A_c_432_n N_A_183_141#_c_865_n 0.0706902f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_471 N_A_M1049_g N_A_183_141#_c_809_n 8.05117e-19 $X=6.125 $Y=2.965 $X2=0
+ $Y2=0
cc_472 N_A_M1064_g N_A_183_141#_c_809_n 0.0361085f $X=6.905 $Y=2.965 $X2=0 $Y2=0
cc_473 N_A_M1070_g N_A_183_141#_c_809_n 0.00227089f $X=7.685 $Y=2.965 $X2=0
+ $Y2=0
cc_474 N_A_c_427_n N_A_183_141#_c_682_n 0.0119333f $X=6.905 $Y=1.565 $X2=0 $Y2=0
cc_475 N_A_c_415_n N_A_183_141#_c_877_n 0.00255636f $X=2.225 $Y=1.565 $X2=0
+ $Y2=0
cc_476 N_A_c_417_n N_A_183_141#_c_877_n 0.00116671f $X=3.005 $Y=1.565 $X2=0
+ $Y2=0
cc_477 N_A_c_431_n N_A_183_141#_c_877_n 0.0259572f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_478 N_A_c_432_n N_A_183_141#_c_877_n 0.00257254f $X=7.685 $Y=1.815 $X2=0
+ $Y2=0
cc_479 N_A_M1006_g N_A_183_141#_c_881_n 0.00316841f $X=2.225 $Y=2.965 $X2=0
+ $Y2=0
cc_480 N_A_c_431_n N_A_183_141#_c_881_n 0.024153f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_481 N_A_c_432_n N_A_183_141#_c_881_n 0.00931804f $X=7.685 $Y=1.815 $X2=0
+ $Y2=0
cc_482 N_A_M1019_g N_A_183_141#_c_884_n 0.00354318f $X=3.785 $Y=2.965 $X2=0
+ $Y2=0
cc_483 N_A_c_431_n N_A_183_141#_c_884_n 0.0272695f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_484 N_A_c_432_n N_A_183_141#_c_884_n 0.0101992f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_485 N_A_c_419_n N_A_183_141#_c_887_n 2.98176e-19 $X=3.785 $Y=1.565 $X2=0
+ $Y2=0
cc_486 N_A_c_431_n N_A_183_141#_c_887_n 0.0165976f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_487 N_A_c_432_n N_A_183_141#_c_887_n 0.00257254f $X=7.685 $Y=1.815 $X2=0
+ $Y2=0
cc_488 N_A_c_427_n N_A_183_141#_c_683_n 0.00681705f $X=6.905 $Y=1.565 $X2=0
+ $Y2=0
cc_489 N_A_M1064_g N_A_183_141#_c_683_n 0.00320206f $X=6.905 $Y=2.965 $X2=0
+ $Y2=0
cc_490 N_A_c_429_n N_A_183_141#_c_683_n 0.00375447f $X=7.685 $Y=1.565 $X2=0
+ $Y2=0
cc_491 N_A_M1070_g N_A_183_141#_c_683_n 0.00510448f $X=7.685 $Y=2.965 $X2=0
+ $Y2=0
cc_492 N_A_c_432_n N_A_183_141#_c_683_n 0.0403801f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_493 N_A_c_429_n N_A_183_141#_c_698_n 0.00942749f $X=7.685 $Y=1.565 $X2=0
+ $Y2=0
cc_494 N_A_c_431_n N_A_183_141#_c_698_n 0.00103228f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_495 N_A_c_432_n N_A_183_141#_c_698_n 0.0183017f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_496 N_A_M1000_g N_VPWR_c_1410_n 0.0688276f $X=0.665 $Y=2.965 $X2=0 $Y2=0
cc_497 N_A_c_431_n N_VPWR_c_1410_n 0.0204297f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_498 N_A_c_432_n N_VPWR_c_1410_n 0.00594552f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_499 N_A_M1000_g N_VPWR_c_1413_n 4.82782e-19 $X=0.665 $Y=2.965 $X2=0 $Y2=0
cc_500 N_A_M1001_g N_VPWR_c_1413_n 0.0590539f $X=1.445 $Y=2.965 $X2=0 $Y2=0
cc_501 N_A_M1006_g N_VPWR_c_1413_n 0.050844f $X=2.225 $Y=2.965 $X2=0 $Y2=0
cc_502 N_A_c_432_n N_VPWR_c_1413_n 4.98839e-19 $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_503 N_A_M1006_g N_VPWR_c_1415_n 4.84763e-19 $X=2.225 $Y=2.965 $X2=0 $Y2=0
cc_504 N_A_M1016_g N_VPWR_c_1415_n 0.0609199f $X=3.005 $Y=2.965 $X2=0 $Y2=0
cc_505 N_A_M1019_g N_VPWR_c_1415_n 0.0481049f $X=3.785 $Y=2.965 $X2=0 $Y2=0
cc_506 N_A_c_432_n N_VPWR_c_1415_n 4.98839e-19 $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_507 N_A_M1019_g N_VPWR_c_1417_n 4.5995e-19 $X=3.785 $Y=2.965 $X2=0 $Y2=0
cc_508 N_A_M1035_g N_VPWR_c_1417_n 0.058787f $X=4.565 $Y=2.965 $X2=0 $Y2=0
cc_509 N_A_M1039_g N_VPWR_c_1417_n 0.0508436f $X=5.345 $Y=2.965 $X2=0 $Y2=0
cc_510 N_A_c_432_n N_VPWR_c_1417_n 4.97715e-19 $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_511 N_A_M1039_g N_VPWR_c_1419_n 4.84763e-19 $X=5.345 $Y=2.965 $X2=0 $Y2=0
cc_512 N_A_M1049_g N_VPWR_c_1419_n 0.0609199f $X=6.125 $Y=2.965 $X2=0 $Y2=0
cc_513 N_A_M1064_g N_VPWR_c_1419_n 0.0481049f $X=6.905 $Y=2.965 $X2=0 $Y2=0
cc_514 N_A_c_432_n N_VPWR_c_1419_n 4.98839e-19 $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_515 N_A_M1064_g N_VPWR_c_1421_n 5.15125e-19 $X=6.905 $Y=2.965 $X2=0 $Y2=0
cc_516 N_A_M1070_g N_VPWR_c_1421_n 0.0848573f $X=7.685 $Y=2.965 $X2=0 $Y2=0
cc_517 N_A_M1000_g N_VPWR_c_1471_n 0.0100933f $X=0.665 $Y=2.965 $X2=0 $Y2=0
cc_518 N_A_M1001_g N_VPWR_c_1471_n 0.00971346f $X=1.445 $Y=2.965 $X2=0 $Y2=0
cc_519 N_A_M1006_g N_VPWR_c_1471_n 0.0104855f $X=2.225 $Y=2.965 $X2=0 $Y2=0
cc_520 N_A_M1016_g N_VPWR_c_1471_n 0.00883212f $X=3.005 $Y=2.965 $X2=0 $Y2=0
cc_521 N_A_M1019_g N_VPWR_c_1471_n 0.0104497f $X=3.785 $Y=2.965 $X2=0 $Y2=0
cc_522 N_A_M1035_g N_VPWR_c_1471_n 0.00969553f $X=4.565 $Y=2.965 $X2=0 $Y2=0
cc_523 N_A_M1039_g N_VPWR_c_1471_n 0.0104855f $X=5.345 $Y=2.965 $X2=0 $Y2=0
cc_524 N_A_M1049_g N_VPWR_c_1471_n 0.00883212f $X=6.125 $Y=2.965 $X2=0 $Y2=0
cc_525 N_A_M1064_g N_VPWR_c_1471_n 0.0104497f $X=6.905 $Y=2.965 $X2=0 $Y2=0
cc_526 N_A_M1070_g N_VPWR_c_1471_n 0.0100929f $X=7.685 $Y=2.965 $X2=0 $Y2=0
cc_527 N_A_c_411_n N_VGND_c_2075_n 0.0413536f $X=0.665 $Y=1.565 $X2=0 $Y2=0
cc_528 N_A_c_413_n N_VGND_c_2075_n 8.88499e-19 $X=1.445 $Y=1.565 $X2=0 $Y2=0
cc_529 N_A_c_431_n N_VGND_c_2075_n 0.0309722f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_530 N_A_c_432_n N_VGND_c_2075_n 0.0048454f $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_531 N_A_c_411_n N_VGND_c_2077_n 0.00101241f $X=0.665 $Y=1.565 $X2=0 $Y2=0
cc_532 N_A_c_413_n N_VGND_c_2077_n 0.0339149f $X=1.445 $Y=1.565 $X2=0 $Y2=0
cc_533 N_A_c_415_n N_VGND_c_2077_n 0.0281515f $X=2.225 $Y=1.565 $X2=0 $Y2=0
cc_534 N_A_c_417_n N_VGND_c_2077_n 7.4453e-19 $X=3.005 $Y=1.565 $X2=0 $Y2=0
cc_535 N_A_c_415_n N_VGND_c_2079_n 7.99935e-19 $X=2.225 $Y=1.565 $X2=0 $Y2=0
cc_536 N_A_c_417_n N_VGND_c_2079_n 0.0309163f $X=3.005 $Y=1.565 $X2=0 $Y2=0
cc_537 N_A_c_419_n N_VGND_c_2079_n 0.032189f $X=3.785 $Y=1.565 $X2=0 $Y2=0
cc_538 N_A_c_421_n N_VGND_c_2079_n 5.19551e-19 $X=4.565 $Y=1.565 $X2=0 $Y2=0
cc_539 N_A_c_419_n N_VGND_c_2081_n 5.04771e-19 $X=3.785 $Y=1.565 $X2=0 $Y2=0
cc_540 N_A_c_421_n N_VGND_c_2081_n 0.0341035f $X=4.565 $Y=1.565 $X2=0 $Y2=0
cc_541 N_A_c_423_n N_VGND_c_2081_n 0.0266615f $X=5.345 $Y=1.565 $X2=0 $Y2=0
cc_542 N_A_c_425_n N_VGND_c_2081_n 7.18649e-19 $X=6.125 $Y=1.565 $X2=0 $Y2=0
cc_543 N_A_c_432_n N_VGND_c_2081_n 3.58496e-19 $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_544 N_A_c_423_n N_VGND_c_2083_n 7.99935e-19 $X=5.345 $Y=1.565 $X2=0 $Y2=0
cc_545 N_A_c_425_n N_VGND_c_2083_n 0.0308964f $X=6.125 $Y=1.565 $X2=0 $Y2=0
cc_546 N_A_c_427_n N_VGND_c_2083_n 0.0321652f $X=6.905 $Y=1.565 $X2=0 $Y2=0
cc_547 N_A_c_429_n N_VGND_c_2083_n 5.19313e-19 $X=7.685 $Y=1.565 $X2=0 $Y2=0
cc_548 N_A_c_432_n N_VGND_c_2083_n 3.59322e-19 $X=7.685 $Y=1.815 $X2=0 $Y2=0
cc_549 N_A_c_411_n N_VGND_c_2117_n 0.0127777f $X=0.665 $Y=1.565 $X2=0 $Y2=0
cc_550 N_A_c_413_n N_VGND_c_2117_n 0.00454157f $X=1.445 $Y=1.565 $X2=0 $Y2=0
cc_551 N_A_c_415_n N_VGND_c_2117_n 0.00710298f $X=2.225 $Y=1.565 $X2=0 $Y2=0
cc_552 N_A_c_417_n N_VGND_c_2117_n 0.00613925f $X=3.005 $Y=1.565 $X2=0 $Y2=0
cc_553 N_A_c_419_n N_VGND_c_2117_n 0.00553692f $X=3.785 $Y=1.565 $X2=0 $Y2=0
cc_554 N_A_c_421_n N_VGND_c_2117_n 0.00393066f $X=4.565 $Y=1.565 $X2=0 $Y2=0
cc_555 N_A_c_423_n N_VGND_c_2117_n 0.00772956f $X=5.345 $Y=1.565 $X2=0 $Y2=0
cc_556 N_A_c_425_n N_VGND_c_2117_n 0.00615492f $X=6.125 $Y=1.565 $X2=0 $Y2=0
cc_557 N_A_c_427_n N_VGND_c_2117_n 0.00553554f $X=6.905 $Y=1.565 $X2=0 $Y2=0
cc_558 N_A_c_429_n N_VGND_c_2117_n 0.00756155f $X=7.685 $Y=1.565 $X2=0 $Y2=0
cc_559 N_A_c_427_n N_VGND_c_2119_n 5.05598e-19 $X=6.905 $Y=1.565 $X2=0 $Y2=0
cc_560 N_A_c_429_n N_VGND_c_2119_n 0.0573231f $X=7.685 $Y=1.565 $X2=0 $Y2=0
cc_561 N_A_183_141#_c_819_n N_VPWR_M1001_d 0.00183555f $X=2.4 $Y=2.125 $X2=0
+ $Y2=0
cc_562 N_A_183_141#_c_837_n N_VPWR_M1016_d 0.00183555f $X=3.94 $Y=2.125 $X2=0
+ $Y2=0
cc_563 N_A_183_141#_c_865_n N_VPWR_M1035_d 0.00188202f $X=5.91 $Y=1.73 $X2=0
+ $Y2=0
cc_564 N_A_183_141#_c_860_n N_VPWR_M1049_d 0.00188651f $X=7.06 $Y=1.73 $X2=-0.33
+ $Y2=-0.265
cc_565 N_A_183_141#_c_797_n N_VPWR_c_1410_n 0.112221f $X=1.055 $Y=2.34 $X2=0
+ $Y2=0
cc_566 N_A_183_141#_c_823_n N_VPWR_c_1410_n 0.00747993f $X=1.16 $Y=2.125 $X2=0
+ $Y2=0
cc_567 N_A_183_141#_c_797_n N_VPWR_c_1413_n 0.0510355f $X=1.055 $Y=2.34 $X2=0
+ $Y2=0
cc_568 N_A_183_141#_c_819_n N_VPWR_c_1413_n 0.0591121f $X=2.4 $Y=2.125 $X2=0
+ $Y2=0
cc_569 N_A_183_141#_c_800_n N_VPWR_c_1413_n 0.0941391f $X=2.615 $Y=2.34 $X2=0
+ $Y2=0
cc_570 N_A_183_141#_c_800_n N_VPWR_c_1415_n 0.0536079f $X=2.615 $Y=2.34 $X2=0
+ $Y2=0
cc_571 N_A_183_141#_c_837_n N_VPWR_c_1415_n 0.0591121f $X=3.94 $Y=2.125 $X2=0
+ $Y2=0
cc_572 N_A_183_141#_c_803_n N_VPWR_c_1415_n 0.0948437f $X=4.175 $Y=2.34 $X2=0
+ $Y2=0
cc_573 N_A_183_141#_c_803_n N_VPWR_c_1417_n 0.0536237f $X=4.175 $Y=2.34 $X2=0
+ $Y2=0
cc_574 N_A_183_141#_c_851_n N_VPWR_c_1417_n 0.0255027f $X=4.8 $Y=2.125 $X2=0
+ $Y2=0
cc_575 N_A_183_141#_c_806_n N_VPWR_c_1417_n 0.0941391f $X=5.735 $Y=2.34 $X2=0
+ $Y2=0
cc_576 N_A_183_141#_c_865_n N_VPWR_c_1417_n 0.0359064f $X=5.91 $Y=1.73 $X2=0
+ $Y2=0
cc_577 N_A_183_141#_c_806_n N_VPWR_c_1419_n 0.0536079f $X=5.735 $Y=2.34 $X2=0
+ $Y2=0
cc_578 N_A_183_141#_c_860_n N_VPWR_c_1419_n 0.0631114f $X=7.06 $Y=1.73 $X2=0
+ $Y2=0
cc_579 N_A_183_141#_c_809_n N_VPWR_c_1419_n 0.0948437f $X=7.295 $Y=2.34 $X2=0
+ $Y2=0
cc_580 N_A_183_141#_M1004_g N_VPWR_c_1421_n 0.0514992f $X=8.705 $Y=2.965 $X2=0
+ $Y2=0
cc_581 N_A_183_141#_c_809_n N_VPWR_c_1421_n 0.0611702f $X=7.295 $Y=2.34 $X2=0
+ $Y2=0
cc_582 N_A_183_141#_c_698_n N_VPWR_c_1421_n 0.0345629f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_583 N_A_183_141#_M1004_g N_VPWR_c_1423_n 6.16464e-19 $X=8.705 $Y=2.965 $X2=0
+ $Y2=0
cc_584 N_A_183_141#_M1011_g N_VPWR_c_1423_n 0.072841f $X=9.485 $Y=2.965 $X2=0
+ $Y2=0
cc_585 N_A_183_141#_M1013_g N_VPWR_c_1423_n 0.0730293f $X=10.265 $Y=2.965 $X2=0
+ $Y2=0
cc_586 N_A_183_141#_M1017_g N_VPWR_c_1423_n 6.16464e-19 $X=11.045 $Y=2.965 $X2=0
+ $Y2=0
cc_587 N_A_183_141#_c_676_n N_VPWR_c_1423_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_588 N_A_183_141#_c_684_n N_VPWR_c_1423_n 0.0279945f $X=10.035 $Y=1.665 $X2=0
+ $Y2=0
cc_589 N_A_183_141#_c_698_n N_VPWR_c_1423_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_590 N_A_183_141#_M1013_g N_VPWR_c_1426_n 6.16464e-19 $X=10.265 $Y=2.965 $X2=0
+ $Y2=0
cc_591 N_A_183_141#_M1017_g N_VPWR_c_1426_n 0.072841f $X=11.045 $Y=2.965 $X2=0
+ $Y2=0
cc_592 N_A_183_141#_M1018_g N_VPWR_c_1426_n 0.0730293f $X=11.825 $Y=2.965 $X2=0
+ $Y2=0
cc_593 N_A_183_141#_M1020_g N_VPWR_c_1426_n 6.16464e-19 $X=12.605 $Y=2.965 $X2=0
+ $Y2=0
cc_594 N_A_183_141#_c_676_n N_VPWR_c_1426_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_595 N_A_183_141#_c_685_n N_VPWR_c_1426_n 0.0279945f $X=11.595 $Y=1.665 $X2=0
+ $Y2=0
cc_596 N_A_183_141#_c_698_n N_VPWR_c_1426_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_597 N_A_183_141#_M1018_g N_VPWR_c_1429_n 6.16464e-19 $X=11.825 $Y=2.965 $X2=0
+ $Y2=0
cc_598 N_A_183_141#_M1020_g N_VPWR_c_1429_n 0.072841f $X=12.605 $Y=2.965 $X2=0
+ $Y2=0
cc_599 N_A_183_141#_M1021_g N_VPWR_c_1429_n 0.0730293f $X=13.385 $Y=2.965 $X2=0
+ $Y2=0
cc_600 N_A_183_141#_M1022_g N_VPWR_c_1429_n 6.16464e-19 $X=14.165 $Y=2.965 $X2=0
+ $Y2=0
cc_601 N_A_183_141#_c_676_n N_VPWR_c_1429_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_602 N_A_183_141#_c_686_n N_VPWR_c_1429_n 0.0279945f $X=13.155 $Y=1.665 $X2=0
+ $Y2=0
cc_603 N_A_183_141#_c_698_n N_VPWR_c_1429_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_604 N_A_183_141#_M1021_g N_VPWR_c_1432_n 6.16464e-19 $X=13.385 $Y=2.965 $X2=0
+ $Y2=0
cc_605 N_A_183_141#_M1022_g N_VPWR_c_1432_n 0.072841f $X=14.165 $Y=2.965 $X2=0
+ $Y2=0
cc_606 N_A_183_141#_M1023_g N_VPWR_c_1432_n 0.0730293f $X=14.945 $Y=2.965 $X2=0
+ $Y2=0
cc_607 N_A_183_141#_M1024_g N_VPWR_c_1432_n 6.16464e-19 $X=15.725 $Y=2.965 $X2=0
+ $Y2=0
cc_608 N_A_183_141#_c_676_n N_VPWR_c_1432_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_609 N_A_183_141#_c_687_n N_VPWR_c_1432_n 0.0279945f $X=14.715 $Y=1.665 $X2=0
+ $Y2=0
cc_610 N_A_183_141#_c_698_n N_VPWR_c_1432_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_611 N_A_183_141#_M1023_g N_VPWR_c_1435_n 6.16464e-19 $X=14.945 $Y=2.965 $X2=0
+ $Y2=0
cc_612 N_A_183_141#_M1024_g N_VPWR_c_1435_n 0.072841f $X=15.725 $Y=2.965 $X2=0
+ $Y2=0
cc_613 N_A_183_141#_M1026_g N_VPWR_c_1435_n 0.0730293f $X=16.505 $Y=2.965 $X2=0
+ $Y2=0
cc_614 N_A_183_141#_M1029_g N_VPWR_c_1435_n 6.16464e-19 $X=17.285 $Y=2.965 $X2=0
+ $Y2=0
cc_615 N_A_183_141#_c_676_n N_VPWR_c_1435_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_616 N_A_183_141#_c_688_n N_VPWR_c_1435_n 0.0279945f $X=16.275 $Y=1.665 $X2=0
+ $Y2=0
cc_617 N_A_183_141#_c_698_n N_VPWR_c_1435_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_618 N_A_183_141#_M1026_g N_VPWR_c_1438_n 6.16464e-19 $X=16.505 $Y=2.965 $X2=0
+ $Y2=0
cc_619 N_A_183_141#_M1029_g N_VPWR_c_1438_n 0.072841f $X=17.285 $Y=2.965 $X2=0
+ $Y2=0
cc_620 N_A_183_141#_M1030_g N_VPWR_c_1438_n 0.0730293f $X=18.065 $Y=2.965 $X2=0
+ $Y2=0
cc_621 N_A_183_141#_M1033_g N_VPWR_c_1438_n 6.16464e-19 $X=18.845 $Y=2.965 $X2=0
+ $Y2=0
cc_622 N_A_183_141#_c_676_n N_VPWR_c_1438_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_623 N_A_183_141#_c_689_n N_VPWR_c_1438_n 0.0279945f $X=17.835 $Y=1.665 $X2=0
+ $Y2=0
cc_624 N_A_183_141#_c_698_n N_VPWR_c_1438_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_625 N_A_183_141#_M1030_g N_VPWR_c_1441_n 6.16464e-19 $X=18.065 $Y=2.965 $X2=0
+ $Y2=0
cc_626 N_A_183_141#_M1033_g N_VPWR_c_1441_n 0.072841f $X=18.845 $Y=2.965 $X2=0
+ $Y2=0
cc_627 N_A_183_141#_M1034_g N_VPWR_c_1441_n 0.0730293f $X=19.625 $Y=2.965 $X2=0
+ $Y2=0
cc_628 N_A_183_141#_M1036_g N_VPWR_c_1441_n 6.16464e-19 $X=20.405 $Y=2.965 $X2=0
+ $Y2=0
cc_629 N_A_183_141#_c_676_n N_VPWR_c_1441_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_630 N_A_183_141#_c_690_n N_VPWR_c_1441_n 0.0279945f $X=19.395 $Y=1.665 $X2=0
+ $Y2=0
cc_631 N_A_183_141#_c_698_n N_VPWR_c_1441_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_632 N_A_183_141#_M1034_g N_VPWR_c_1444_n 5.01535e-19 $X=19.625 $Y=2.965 $X2=0
+ $Y2=0
cc_633 N_A_183_141#_M1036_g N_VPWR_c_1444_n 0.058402f $X=20.405 $Y=2.965 $X2=0
+ $Y2=0
cc_634 N_A_183_141#_M1037_g N_VPWR_c_1444_n 0.0401385f $X=21.185 $Y=2.965 $X2=0
+ $Y2=0
cc_635 N_A_183_141#_c_676_n N_VPWR_c_1444_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_636 N_A_183_141#_c_691_n N_VPWR_c_1444_n 0.0223351f $X=20.945 $Y=1.665 $X2=0
+ $Y2=0
cc_637 N_A_183_141#_c_698_n N_VPWR_c_1444_n 0.00235405f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_638 N_A_183_141#_M1037_g N_VPWR_c_1447_n 6.16464e-19 $X=21.185 $Y=2.965 $X2=0
+ $Y2=0
cc_639 N_A_183_141#_M1041_g N_VPWR_c_1447_n 0.072841f $X=21.965 $Y=2.965 $X2=0
+ $Y2=0
cc_640 N_A_183_141#_M1042_g N_VPWR_c_1447_n 0.0730293f $X=22.745 $Y=2.965 $X2=0
+ $Y2=0
cc_641 N_A_183_141#_M1045_g N_VPWR_c_1447_n 6.16464e-19 $X=23.525 $Y=2.965 $X2=0
+ $Y2=0
cc_642 N_A_183_141#_c_676_n N_VPWR_c_1447_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_643 N_A_183_141#_c_692_n N_VPWR_c_1447_n 0.0279945f $X=22.515 $Y=1.665 $X2=0
+ $Y2=0
cc_644 N_A_183_141#_c_698_n N_VPWR_c_1447_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_645 N_A_183_141#_M1042_g N_VPWR_c_1450_n 6.16464e-19 $X=22.745 $Y=2.965 $X2=0
+ $Y2=0
cc_646 N_A_183_141#_M1045_g N_VPWR_c_1450_n 0.072841f $X=23.525 $Y=2.965 $X2=0
+ $Y2=0
cc_647 N_A_183_141#_M1046_g N_VPWR_c_1450_n 0.0730293f $X=24.305 $Y=2.965 $X2=0
+ $Y2=0
cc_648 N_A_183_141#_M1050_g N_VPWR_c_1450_n 6.16464e-19 $X=25.085 $Y=2.965 $X2=0
+ $Y2=0
cc_649 N_A_183_141#_c_676_n N_VPWR_c_1450_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_650 N_A_183_141#_c_693_n N_VPWR_c_1450_n 0.0279945f $X=24.075 $Y=1.665 $X2=0
+ $Y2=0
cc_651 N_A_183_141#_c_698_n N_VPWR_c_1450_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_652 N_A_183_141#_M1046_g N_VPWR_c_1453_n 6.16464e-19 $X=24.305 $Y=2.965 $X2=0
+ $Y2=0
cc_653 N_A_183_141#_M1050_g N_VPWR_c_1453_n 0.072841f $X=25.085 $Y=2.965 $X2=0
+ $Y2=0
cc_654 N_A_183_141#_M1054_g N_VPWR_c_1453_n 0.0730293f $X=25.865 $Y=2.965 $X2=0
+ $Y2=0
cc_655 N_A_183_141#_M1055_g N_VPWR_c_1453_n 6.16464e-19 $X=26.645 $Y=2.965 $X2=0
+ $Y2=0
cc_656 N_A_183_141#_c_676_n N_VPWR_c_1453_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_657 N_A_183_141#_c_694_n N_VPWR_c_1453_n 0.0279945f $X=25.635 $Y=1.665 $X2=0
+ $Y2=0
cc_658 N_A_183_141#_c_698_n N_VPWR_c_1453_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_659 N_A_183_141#_M1054_g N_VPWR_c_1456_n 6.16464e-19 $X=25.865 $Y=2.965 $X2=0
+ $Y2=0
cc_660 N_A_183_141#_M1055_g N_VPWR_c_1456_n 0.072841f $X=26.645 $Y=2.965 $X2=0
+ $Y2=0
cc_661 N_A_183_141#_M1059_g N_VPWR_c_1456_n 0.0730293f $X=27.425 $Y=2.965 $X2=0
+ $Y2=0
cc_662 N_A_183_141#_M1060_g N_VPWR_c_1456_n 6.16464e-19 $X=28.205 $Y=2.965 $X2=0
+ $Y2=0
cc_663 N_A_183_141#_c_676_n N_VPWR_c_1456_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_664 N_A_183_141#_c_695_n N_VPWR_c_1456_n 0.0279945f $X=27.195 $Y=1.665 $X2=0
+ $Y2=0
cc_665 N_A_183_141#_c_698_n N_VPWR_c_1456_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_666 N_A_183_141#_M1059_g N_VPWR_c_1459_n 6.16464e-19 $X=27.425 $Y=2.965 $X2=0
+ $Y2=0
cc_667 N_A_183_141#_M1060_g N_VPWR_c_1459_n 0.072841f $X=28.205 $Y=2.965 $X2=0
+ $Y2=0
cc_668 N_A_183_141#_M1063_g N_VPWR_c_1459_n 0.0730293f $X=28.985 $Y=2.965 $X2=0
+ $Y2=0
cc_669 N_A_183_141#_M1065_g N_VPWR_c_1459_n 6.16464e-19 $X=29.765 $Y=2.965 $X2=0
+ $Y2=0
cc_670 N_A_183_141#_c_676_n N_VPWR_c_1459_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_671 N_A_183_141#_c_696_n N_VPWR_c_1459_n 0.0279945f $X=28.755 $Y=1.665 $X2=0
+ $Y2=0
cc_672 N_A_183_141#_c_698_n N_VPWR_c_1459_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_673 N_A_183_141#_M1063_g N_VPWR_c_1462_n 6.16464e-19 $X=28.985 $Y=2.965 $X2=0
+ $Y2=0
cc_674 N_A_183_141#_M1065_g N_VPWR_c_1462_n 0.072841f $X=29.765 $Y=2.965 $X2=0
+ $Y2=0
cc_675 N_A_183_141#_M1066_g N_VPWR_c_1462_n 0.0730293f $X=30.545 $Y=2.965 $X2=0
+ $Y2=0
cc_676 N_A_183_141#_M1073_g N_VPWR_c_1462_n 6.16464e-19 $X=31.325 $Y=2.965 $X2=0
+ $Y2=0
cc_677 N_A_183_141#_c_676_n N_VPWR_c_1462_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_678 N_A_183_141#_c_697_n N_VPWR_c_1462_n 0.0279945f $X=30.315 $Y=1.665 $X2=0
+ $Y2=0
cc_679 N_A_183_141#_c_698_n N_VPWR_c_1462_n 0.00839812f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_680 N_A_183_141#_M1066_g N_VPWR_c_1465_n 6.16464e-19 $X=30.545 $Y=2.965 $X2=0
+ $Y2=0
cc_681 N_A_183_141#_M1073_g N_VPWR_c_1465_n 0.072841f $X=31.325 $Y=2.965 $X2=0
+ $Y2=0
cc_682 N_A_183_141#_M1075_g N_VPWR_c_1465_n 0.0750023f $X=32.105 $Y=2.965 $X2=0
+ $Y2=0
cc_683 N_A_183_141#_c_676_n N_VPWR_c_1465_n 0.00264079f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_684 N_A_183_141#_M1080_g N_VPWR_c_1465_n 6.16464e-19 $X=32.885 $Y=2.965 $X2=0
+ $Y2=0
cc_685 N_A_183_141#_c_698_n N_VPWR_c_1465_n 0.00668272f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_686 N_A_183_141#_c_699_n N_VPWR_c_1465_n 0.0279945f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_687 N_A_183_141#_M1075_g N_VPWR_c_1468_n 4.37802e-19 $X=32.105 $Y=2.965 $X2=0
+ $Y2=0
cc_688 N_A_183_141#_M1080_g N_VPWR_c_1468_n 0.0636473f $X=32.885 $Y=2.965 $X2=0
+ $Y2=0
cc_689 N_A_183_141#_M1000_s N_VPWR_c_1471_n 0.00137624f $X=0.915 $Y=2.215 $X2=0
+ $Y2=0
cc_690 N_A_183_141#_M1006_s N_VPWR_c_1471_n 0.00179328f $X=2.475 $Y=2.215 $X2=0
+ $Y2=0
cc_691 N_A_183_141#_M1019_s N_VPWR_c_1471_n 9.59196e-19 $X=4.035 $Y=2.215 $X2=0
+ $Y2=0
cc_692 N_A_183_141#_M1039_s N_VPWR_c_1471_n 0.00179328f $X=5.595 $Y=2.215 $X2=0
+ $Y2=0
cc_693 N_A_183_141#_M1064_s N_VPWR_c_1471_n 9.59196e-19 $X=7.155 $Y=2.215 $X2=0
+ $Y2=0
cc_694 N_A_183_141#_M1004_g N_VPWR_c_1471_n 0.0276818f $X=8.705 $Y=2.965 $X2=0
+ $Y2=0
cc_695 N_A_183_141#_M1011_g N_VPWR_c_1471_n 0.00965647f $X=9.485 $Y=2.965 $X2=0
+ $Y2=0
cc_696 N_A_183_141#_M1013_g N_VPWR_c_1471_n 0.00965647f $X=10.265 $Y=2.965 $X2=0
+ $Y2=0
cc_697 N_A_183_141#_M1017_g N_VPWR_c_1471_n 0.00965647f $X=11.045 $Y=2.965 $X2=0
+ $Y2=0
cc_698 N_A_183_141#_M1018_g N_VPWR_c_1471_n 0.00965647f $X=11.825 $Y=2.965 $X2=0
+ $Y2=0
cc_699 N_A_183_141#_M1020_g N_VPWR_c_1471_n 0.00965647f $X=12.605 $Y=2.965 $X2=0
+ $Y2=0
cc_700 N_A_183_141#_M1021_g N_VPWR_c_1471_n 0.00965647f $X=13.385 $Y=2.965 $X2=0
+ $Y2=0
cc_701 N_A_183_141#_M1022_g N_VPWR_c_1471_n 0.00965647f $X=14.165 $Y=2.965 $X2=0
+ $Y2=0
cc_702 N_A_183_141#_M1023_g N_VPWR_c_1471_n 0.00965647f $X=14.945 $Y=2.965 $X2=0
+ $Y2=0
cc_703 N_A_183_141#_M1024_g N_VPWR_c_1471_n 0.00965647f $X=15.725 $Y=2.965 $X2=0
+ $Y2=0
cc_704 N_A_183_141#_M1026_g N_VPWR_c_1471_n 0.00965647f $X=16.505 $Y=2.965 $X2=0
+ $Y2=0
cc_705 N_A_183_141#_M1029_g N_VPWR_c_1471_n 0.00965647f $X=17.285 $Y=2.965 $X2=0
+ $Y2=0
cc_706 N_A_183_141#_M1030_g N_VPWR_c_1471_n 0.00965647f $X=18.065 $Y=2.965 $X2=0
+ $Y2=0
cc_707 N_A_183_141#_M1033_g N_VPWR_c_1471_n 0.00965647f $X=18.845 $Y=2.965 $X2=0
+ $Y2=0
cc_708 N_A_183_141#_M1034_g N_VPWR_c_1471_n 0.00965647f $X=19.625 $Y=2.965 $X2=0
+ $Y2=0
cc_709 N_A_183_141#_M1036_g N_VPWR_c_1471_n 0.00965647f $X=20.405 $Y=2.965 $X2=0
+ $Y2=0
cc_710 N_A_183_141#_M1037_g N_VPWR_c_1471_n 0.0264237f $X=21.185 $Y=2.965 $X2=0
+ $Y2=0
cc_711 N_A_183_141#_M1041_g N_VPWR_c_1471_n 0.00965647f $X=21.965 $Y=2.965 $X2=0
+ $Y2=0
cc_712 N_A_183_141#_M1042_g N_VPWR_c_1471_n 0.00965647f $X=22.745 $Y=2.965 $X2=0
+ $Y2=0
cc_713 N_A_183_141#_M1045_g N_VPWR_c_1471_n 0.00965647f $X=23.525 $Y=2.965 $X2=0
+ $Y2=0
cc_714 N_A_183_141#_M1046_g N_VPWR_c_1471_n 0.00965647f $X=24.305 $Y=2.965 $X2=0
+ $Y2=0
cc_715 N_A_183_141#_M1050_g N_VPWR_c_1471_n 0.00965647f $X=25.085 $Y=2.965 $X2=0
+ $Y2=0
cc_716 N_A_183_141#_M1054_g N_VPWR_c_1471_n 0.00965647f $X=25.865 $Y=2.965 $X2=0
+ $Y2=0
cc_717 N_A_183_141#_M1055_g N_VPWR_c_1471_n 0.00965647f $X=26.645 $Y=2.965 $X2=0
+ $Y2=0
cc_718 N_A_183_141#_M1059_g N_VPWR_c_1471_n 0.00965647f $X=27.425 $Y=2.965 $X2=0
+ $Y2=0
cc_719 N_A_183_141#_M1060_g N_VPWR_c_1471_n 0.00965647f $X=28.205 $Y=2.965 $X2=0
+ $Y2=0
cc_720 N_A_183_141#_M1063_g N_VPWR_c_1471_n 0.00965647f $X=28.985 $Y=2.965 $X2=0
+ $Y2=0
cc_721 N_A_183_141#_M1065_g N_VPWR_c_1471_n 0.00965647f $X=29.765 $Y=2.965 $X2=0
+ $Y2=0
cc_722 N_A_183_141#_M1066_g N_VPWR_c_1471_n 0.00965647f $X=30.545 $Y=2.965 $X2=0
+ $Y2=0
cc_723 N_A_183_141#_M1073_g N_VPWR_c_1471_n 0.00965647f $X=31.325 $Y=2.965 $X2=0
+ $Y2=0
cc_724 N_A_183_141#_M1075_g N_VPWR_c_1471_n 0.00965647f $X=32.105 $Y=2.965 $X2=0
+ $Y2=0
cc_725 N_A_183_141#_M1080_g N_VPWR_c_1471_n 0.0101127f $X=32.885 $Y=2.965 $X2=0
+ $Y2=0
cc_726 N_A_183_141#_c_797_n N_VPWR_c_1471_n 0.0381773f $X=1.055 $Y=2.34 $X2=0
+ $Y2=0
cc_727 N_A_183_141#_c_800_n N_VPWR_c_1471_n 0.0394745f $X=2.615 $Y=2.34 $X2=0
+ $Y2=0
cc_728 N_A_183_141#_c_803_n N_VPWR_c_1471_n 0.043412f $X=4.175 $Y=2.34 $X2=0
+ $Y2=0
cc_729 N_A_183_141#_c_806_n N_VPWR_c_1471_n 0.0394745f $X=5.735 $Y=2.34 $X2=0
+ $Y2=0
cc_730 N_A_183_141#_c_809_n N_VPWR_c_1471_n 0.043412f $X=7.295 $Y=2.34 $X2=0
+ $Y2=0
cc_731 N_A_183_141#_c_614_n N_X_c_1741_n 0.025164f $X=8.705 $Y=1.565 $X2=0 $Y2=0
cc_732 N_A_183_141#_M1004_g N_X_c_1741_n 0.0528856f $X=8.705 $Y=2.965 $X2=0
+ $Y2=0
cc_733 N_A_183_141#_c_616_n N_X_c_1741_n 0.0191337f $X=9.485 $Y=1.565 $X2=0
+ $Y2=0
cc_734 N_A_183_141#_M1011_g N_X_c_1741_n 0.0341245f $X=9.485 $Y=2.965 $X2=0
+ $Y2=0
cc_735 N_A_183_141#_c_676_n N_X_c_1741_n 0.0432451f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_736 N_A_183_141#_c_684_n N_X_c_1741_n 0.0152142f $X=10.035 $Y=1.665 $X2=0
+ $Y2=0
cc_737 N_A_183_141#_c_698_n N_X_c_1741_n 0.0458449f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_738 N_A_183_141#_c_618_n N_X_c_1744_n 0.0191337f $X=10.265 $Y=1.565 $X2=0
+ $Y2=0
cc_739 N_A_183_141#_M1013_g N_X_c_1744_n 0.0341245f $X=10.265 $Y=2.965 $X2=0
+ $Y2=0
cc_740 N_A_183_141#_c_620_n N_X_c_1744_n 0.0191337f $X=11.045 $Y=1.565 $X2=0
+ $Y2=0
cc_741 N_A_183_141#_M1017_g N_X_c_1744_n 0.0341245f $X=11.045 $Y=2.965 $X2=0
+ $Y2=0
cc_742 N_A_183_141#_c_676_n N_X_c_1744_n 0.0384414f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_743 N_A_183_141#_c_684_n N_X_c_1744_n 0.0131079f $X=10.035 $Y=1.665 $X2=0
+ $Y2=0
cc_744 N_A_183_141#_c_685_n N_X_c_1744_n 0.0152142f $X=11.595 $Y=1.665 $X2=0
+ $Y2=0
cc_745 N_A_183_141#_c_698_n N_X_c_1744_n 0.0427559f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_746 N_A_183_141#_c_622_n N_X_c_1747_n 0.0191337f $X=11.825 $Y=1.565 $X2=0
+ $Y2=0
cc_747 N_A_183_141#_M1018_g N_X_c_1747_n 0.0341245f $X=11.825 $Y=2.965 $X2=0
+ $Y2=0
cc_748 N_A_183_141#_c_624_n N_X_c_1747_n 0.0191337f $X=12.605 $Y=1.565 $X2=0
+ $Y2=0
cc_749 N_A_183_141#_M1020_g N_X_c_1747_n 0.0341245f $X=12.605 $Y=2.965 $X2=0
+ $Y2=0
cc_750 N_A_183_141#_c_676_n N_X_c_1747_n 0.0384414f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_751 N_A_183_141#_c_685_n N_X_c_1747_n 0.0131079f $X=11.595 $Y=1.665 $X2=0
+ $Y2=0
cc_752 N_A_183_141#_c_686_n N_X_c_1747_n 0.0152142f $X=13.155 $Y=1.665 $X2=0
+ $Y2=0
cc_753 N_A_183_141#_c_698_n N_X_c_1747_n 0.0427559f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_754 N_A_183_141#_c_626_n N_X_c_1750_n 0.0191337f $X=13.385 $Y=1.565 $X2=0
+ $Y2=0
cc_755 N_A_183_141#_M1021_g N_X_c_1750_n 0.0341245f $X=13.385 $Y=2.965 $X2=0
+ $Y2=0
cc_756 N_A_183_141#_c_628_n N_X_c_1750_n 0.0191337f $X=14.165 $Y=1.565 $X2=0
+ $Y2=0
cc_757 N_A_183_141#_M1022_g N_X_c_1750_n 0.0341245f $X=14.165 $Y=2.965 $X2=0
+ $Y2=0
cc_758 N_A_183_141#_c_676_n N_X_c_1750_n 0.0384414f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_759 N_A_183_141#_c_686_n N_X_c_1750_n 0.0131079f $X=13.155 $Y=1.665 $X2=0
+ $Y2=0
cc_760 N_A_183_141#_c_687_n N_X_c_1750_n 0.0152142f $X=14.715 $Y=1.665 $X2=0
+ $Y2=0
cc_761 N_A_183_141#_c_698_n N_X_c_1750_n 0.0427559f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_762 N_A_183_141#_c_630_n N_X_c_1753_n 0.0191337f $X=14.945 $Y=1.565 $X2=0
+ $Y2=0
cc_763 N_A_183_141#_M1023_g N_X_c_1753_n 0.0341245f $X=14.945 $Y=2.965 $X2=0
+ $Y2=0
cc_764 N_A_183_141#_c_632_n N_X_c_1753_n 0.0191337f $X=15.725 $Y=1.565 $X2=0
+ $Y2=0
cc_765 N_A_183_141#_M1024_g N_X_c_1753_n 0.0341245f $X=15.725 $Y=2.965 $X2=0
+ $Y2=0
cc_766 N_A_183_141#_c_676_n N_X_c_1753_n 0.0384414f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_767 N_A_183_141#_c_687_n N_X_c_1753_n 0.0131079f $X=14.715 $Y=1.665 $X2=0
+ $Y2=0
cc_768 N_A_183_141#_c_688_n N_X_c_1753_n 0.0152142f $X=16.275 $Y=1.665 $X2=0
+ $Y2=0
cc_769 N_A_183_141#_c_698_n N_X_c_1753_n 0.0427559f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_770 N_A_183_141#_c_634_n N_X_c_1756_n 0.0191337f $X=16.505 $Y=1.565 $X2=0
+ $Y2=0
cc_771 N_A_183_141#_M1026_g N_X_c_1756_n 0.0341245f $X=16.505 $Y=2.965 $X2=0
+ $Y2=0
cc_772 N_A_183_141#_c_636_n N_X_c_1756_n 0.0191337f $X=17.285 $Y=1.565 $X2=0
+ $Y2=0
cc_773 N_A_183_141#_M1029_g N_X_c_1756_n 0.0341245f $X=17.285 $Y=2.965 $X2=0
+ $Y2=0
cc_774 N_A_183_141#_c_676_n N_X_c_1756_n 0.0384414f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_775 N_A_183_141#_c_688_n N_X_c_1756_n 0.0131079f $X=16.275 $Y=1.665 $X2=0
+ $Y2=0
cc_776 N_A_183_141#_c_689_n N_X_c_1756_n 0.0152142f $X=17.835 $Y=1.665 $X2=0
+ $Y2=0
cc_777 N_A_183_141#_c_698_n N_X_c_1756_n 0.0427559f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_778 N_A_183_141#_c_638_n N_X_c_1759_n 0.0191337f $X=18.065 $Y=1.565 $X2=0
+ $Y2=0
cc_779 N_A_183_141#_M1030_g N_X_c_1759_n 0.0341245f $X=18.065 $Y=2.965 $X2=0
+ $Y2=0
cc_780 N_A_183_141#_c_640_n N_X_c_1759_n 0.0191337f $X=18.845 $Y=1.565 $X2=0
+ $Y2=0
cc_781 N_A_183_141#_M1033_g N_X_c_1759_n 0.0341245f $X=18.845 $Y=2.965 $X2=0
+ $Y2=0
cc_782 N_A_183_141#_c_676_n N_X_c_1759_n 0.0384414f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_783 N_A_183_141#_c_689_n N_X_c_1759_n 0.0131079f $X=17.835 $Y=1.665 $X2=0
+ $Y2=0
cc_784 N_A_183_141#_c_690_n N_X_c_1759_n 0.0152142f $X=19.395 $Y=1.665 $X2=0
+ $Y2=0
cc_785 N_A_183_141#_c_698_n N_X_c_1759_n 0.0427559f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_786 N_A_183_141#_c_642_n N_X_c_1762_n 0.0193861f $X=19.625 $Y=1.565 $X2=0
+ $Y2=0
cc_787 N_A_183_141#_M1034_g N_X_c_1762_n 0.0344467f $X=19.625 $Y=2.965 $X2=0
+ $Y2=0
cc_788 N_A_183_141#_c_644_n N_X_c_1762_n 0.0226072f $X=20.405 $Y=1.565 $X2=0
+ $Y2=0
cc_789 N_A_183_141#_M1036_g N_X_c_1762_n 0.0436049f $X=20.405 $Y=2.965 $X2=0
+ $Y2=0
cc_790 N_A_183_141#_c_646_n N_X_c_1762_n 5.10774e-19 $X=21.185 $Y=1.565 $X2=0
+ $Y2=0
cc_791 N_A_183_141#_M1037_g N_X_c_1762_n 9.65539e-19 $X=21.185 $Y=2.965 $X2=0
+ $Y2=0
cc_792 N_A_183_141#_c_676_n N_X_c_1762_n 0.040836f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_793 N_A_183_141#_c_690_n N_X_c_1762_n 0.013207f $X=19.395 $Y=1.665 $X2=0
+ $Y2=0
cc_794 N_A_183_141#_c_691_n N_X_c_1762_n 0.0233521f $X=20.945 $Y=1.665 $X2=0
+ $Y2=0
cc_795 N_A_183_141#_c_698_n N_X_c_1762_n 0.0506394f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_796 N_A_183_141#_c_646_n N_X_c_1765_n 0.025182f $X=21.185 $Y=1.565 $X2=0
+ $Y2=0
cc_797 N_A_183_141#_M1037_g N_X_c_1765_n 0.0494356f $X=21.185 $Y=2.965 $X2=0
+ $Y2=0
cc_798 N_A_183_141#_c_648_n N_X_c_1765_n 0.0191337f $X=21.965 $Y=1.565 $X2=0
+ $Y2=0
cc_799 N_A_183_141#_M1041_g N_X_c_1765_n 0.0341245f $X=21.965 $Y=2.965 $X2=0
+ $Y2=0
cc_800 N_A_183_141#_c_676_n N_X_c_1765_n 0.0385516f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_801 N_A_183_141#_c_691_n N_X_c_1765_n 0.0126553f $X=20.945 $Y=1.665 $X2=0
+ $Y2=0
cc_802 N_A_183_141#_c_692_n N_X_c_1765_n 0.0152142f $X=22.515 $Y=1.665 $X2=0
+ $Y2=0
cc_803 N_A_183_141#_c_698_n N_X_c_1765_n 0.042833f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_804 N_A_183_141#_c_650_n N_X_c_1768_n 0.0191337f $X=22.745 $Y=1.565 $X2=0
+ $Y2=0
cc_805 N_A_183_141#_M1042_g N_X_c_1768_n 0.0341245f $X=22.745 $Y=2.965 $X2=0
+ $Y2=0
cc_806 N_A_183_141#_c_652_n N_X_c_1768_n 0.0191337f $X=23.525 $Y=1.565 $X2=0
+ $Y2=0
cc_807 N_A_183_141#_M1045_g N_X_c_1768_n 0.0341245f $X=23.525 $Y=2.965 $X2=0
+ $Y2=0
cc_808 N_A_183_141#_c_676_n N_X_c_1768_n 0.0384414f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_809 N_A_183_141#_c_692_n N_X_c_1768_n 0.0131079f $X=22.515 $Y=1.665 $X2=0
+ $Y2=0
cc_810 N_A_183_141#_c_693_n N_X_c_1768_n 0.0152142f $X=24.075 $Y=1.665 $X2=0
+ $Y2=0
cc_811 N_A_183_141#_c_698_n N_X_c_1768_n 0.0427559f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_812 N_A_183_141#_c_654_n N_X_c_1771_n 0.0191337f $X=24.305 $Y=1.565 $X2=0
+ $Y2=0
cc_813 N_A_183_141#_M1046_g N_X_c_1771_n 0.0341245f $X=24.305 $Y=2.965 $X2=0
+ $Y2=0
cc_814 N_A_183_141#_c_656_n N_X_c_1771_n 0.0191337f $X=25.085 $Y=1.565 $X2=0
+ $Y2=0
cc_815 N_A_183_141#_M1050_g N_X_c_1771_n 0.0341245f $X=25.085 $Y=2.965 $X2=0
+ $Y2=0
cc_816 N_A_183_141#_c_676_n N_X_c_1771_n 0.0384414f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_817 N_A_183_141#_c_693_n N_X_c_1771_n 0.0131079f $X=24.075 $Y=1.665 $X2=0
+ $Y2=0
cc_818 N_A_183_141#_c_694_n N_X_c_1771_n 0.0152142f $X=25.635 $Y=1.665 $X2=0
+ $Y2=0
cc_819 N_A_183_141#_c_698_n N_X_c_1771_n 0.0427559f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_820 N_A_183_141#_c_658_n N_X_c_1774_n 0.0191337f $X=25.865 $Y=1.565 $X2=0
+ $Y2=0
cc_821 N_A_183_141#_M1054_g N_X_c_1774_n 0.0341245f $X=25.865 $Y=2.965 $X2=0
+ $Y2=0
cc_822 N_A_183_141#_c_660_n N_X_c_1774_n 0.0191337f $X=26.645 $Y=1.565 $X2=0
+ $Y2=0
cc_823 N_A_183_141#_M1055_g N_X_c_1774_n 0.0341245f $X=26.645 $Y=2.965 $X2=0
+ $Y2=0
cc_824 N_A_183_141#_c_676_n N_X_c_1774_n 0.0384414f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_825 N_A_183_141#_c_694_n N_X_c_1774_n 0.0131079f $X=25.635 $Y=1.665 $X2=0
+ $Y2=0
cc_826 N_A_183_141#_c_695_n N_X_c_1774_n 0.0152142f $X=27.195 $Y=1.665 $X2=0
+ $Y2=0
cc_827 N_A_183_141#_c_698_n N_X_c_1774_n 0.0427559f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_828 N_A_183_141#_c_662_n N_X_c_1777_n 0.0191337f $X=27.425 $Y=1.565 $X2=0
+ $Y2=0
cc_829 N_A_183_141#_M1059_g N_X_c_1777_n 0.0341245f $X=27.425 $Y=2.965 $X2=0
+ $Y2=0
cc_830 N_A_183_141#_c_664_n N_X_c_1777_n 0.0191337f $X=28.205 $Y=1.565 $X2=0
+ $Y2=0
cc_831 N_A_183_141#_M1060_g N_X_c_1777_n 0.0341245f $X=28.205 $Y=2.965 $X2=0
+ $Y2=0
cc_832 N_A_183_141#_c_676_n N_X_c_1777_n 0.0384414f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_833 N_A_183_141#_c_695_n N_X_c_1777_n 0.0131079f $X=27.195 $Y=1.665 $X2=0
+ $Y2=0
cc_834 N_A_183_141#_c_696_n N_X_c_1777_n 0.0152142f $X=28.755 $Y=1.665 $X2=0
+ $Y2=0
cc_835 N_A_183_141#_c_698_n N_X_c_1777_n 0.0427559f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_836 N_A_183_141#_c_666_n N_X_c_1780_n 0.0191337f $X=28.985 $Y=1.565 $X2=0
+ $Y2=0
cc_837 N_A_183_141#_M1063_g N_X_c_1780_n 0.0341245f $X=28.985 $Y=2.965 $X2=0
+ $Y2=0
cc_838 N_A_183_141#_c_668_n N_X_c_1780_n 0.0191337f $X=29.765 $Y=1.565 $X2=0
+ $Y2=0
cc_839 N_A_183_141#_M1065_g N_X_c_1780_n 0.0341245f $X=29.765 $Y=2.965 $X2=0
+ $Y2=0
cc_840 N_A_183_141#_c_676_n N_X_c_1780_n 0.0384414f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_841 N_A_183_141#_c_696_n N_X_c_1780_n 0.0131079f $X=28.755 $Y=1.665 $X2=0
+ $Y2=0
cc_842 N_A_183_141#_c_697_n N_X_c_1780_n 0.0152142f $X=30.315 $Y=1.665 $X2=0
+ $Y2=0
cc_843 N_A_183_141#_c_698_n N_X_c_1780_n 0.0427559f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_844 N_A_183_141#_c_670_n N_X_c_1783_n 0.0191337f $X=30.545 $Y=1.565 $X2=0
+ $Y2=0
cc_845 N_A_183_141#_M1066_g N_X_c_1783_n 0.0341245f $X=30.545 $Y=2.965 $X2=0
+ $Y2=0
cc_846 N_A_183_141#_c_672_n N_X_c_1783_n 0.0191337f $X=31.325 $Y=1.565 $X2=0
+ $Y2=0
cc_847 N_A_183_141#_M1073_g N_X_c_1783_n 0.0341245f $X=31.325 $Y=2.965 $X2=0
+ $Y2=0
cc_848 N_A_183_141#_c_676_n N_X_c_1783_n 0.0384414f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_849 N_A_183_141#_c_697_n N_X_c_1783_n 0.0131079f $X=30.315 $Y=1.665 $X2=0
+ $Y2=0
cc_850 N_A_183_141#_c_698_n N_X_c_1783_n 0.0427559f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_851 N_A_183_141#_c_699_n N_X_c_1783_n 0.0152142f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_852 N_A_183_141#_c_674_n N_X_c_1786_n 0.0193104f $X=32.105 $Y=1.565 $X2=0
+ $Y2=0
cc_853 N_A_183_141#_M1075_g N_X_c_1786_n 0.0344467f $X=32.105 $Y=2.965 $X2=0
+ $Y2=0
cc_854 N_A_183_141#_c_676_n N_X_c_1786_n 0.0769669f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_855 N_A_183_141#_M1080_g N_X_c_1786_n 0.0494075f $X=32.885 $Y=2.965 $X2=0
+ $Y2=0
cc_856 N_A_183_141#_c_698_n N_X_c_1786_n 0.00677521f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_857 N_A_183_141#_c_699_n N_X_c_1786_n 0.0129738f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_858 N_A_183_141#_M1011_g N_X_c_1916_n 0.0101772f $X=9.485 $Y=2.965 $X2=0
+ $Y2=0
cc_859 N_A_183_141#_M1013_g N_X_c_1916_n 0.0101772f $X=10.265 $Y=2.965 $X2=0
+ $Y2=0
cc_860 N_A_183_141#_M1017_g N_X_c_1916_n 0.0101772f $X=11.045 $Y=2.965 $X2=0
+ $Y2=0
cc_861 N_A_183_141#_M1018_g N_X_c_1916_n 0.0101772f $X=11.825 $Y=2.965 $X2=0
+ $Y2=0
cc_862 N_A_183_141#_M1020_g N_X_c_1916_n 0.0101772f $X=12.605 $Y=2.965 $X2=0
+ $Y2=0
cc_863 N_A_183_141#_M1021_g N_X_c_1916_n 0.0101772f $X=13.385 $Y=2.965 $X2=0
+ $Y2=0
cc_864 N_A_183_141#_M1022_g N_X_c_1916_n 0.0101772f $X=14.165 $Y=2.965 $X2=0
+ $Y2=0
cc_865 N_A_183_141#_M1023_g N_X_c_1916_n 0.0101772f $X=14.945 $Y=2.965 $X2=0
+ $Y2=0
cc_866 N_A_183_141#_M1024_g N_X_c_1916_n 0.0101772f $X=15.725 $Y=2.965 $X2=0
+ $Y2=0
cc_867 N_A_183_141#_M1026_g N_X_c_1916_n 0.0101772f $X=16.505 $Y=2.965 $X2=0
+ $Y2=0
cc_868 N_A_183_141#_M1029_g N_X_c_1916_n 0.0101772f $X=17.285 $Y=2.965 $X2=0
+ $Y2=0
cc_869 N_A_183_141#_M1030_g N_X_c_1916_n 0.0101772f $X=18.065 $Y=2.965 $X2=0
+ $Y2=0
cc_870 N_A_183_141#_M1033_g N_X_c_1916_n 0.0101772f $X=18.845 $Y=2.965 $X2=0
+ $Y2=0
cc_871 N_A_183_141#_M1034_g N_X_c_1916_n 0.0101772f $X=19.625 $Y=2.965 $X2=0
+ $Y2=0
cc_872 N_A_183_141#_M1036_g N_X_c_1916_n 0.0101772f $X=20.405 $Y=2.965 $X2=0
+ $Y2=0
cc_873 N_A_183_141#_M1037_g N_X_c_1916_n 0.0286069f $X=21.185 $Y=2.965 $X2=0
+ $Y2=0
cc_874 N_A_183_141#_M1041_g N_X_c_1916_n 0.0101772f $X=21.965 $Y=2.965 $X2=0
+ $Y2=0
cc_875 N_A_183_141#_M1042_g N_X_c_1916_n 0.0101772f $X=22.745 $Y=2.965 $X2=0
+ $Y2=0
cc_876 N_A_183_141#_M1045_g N_X_c_1916_n 0.0101772f $X=23.525 $Y=2.965 $X2=0
+ $Y2=0
cc_877 N_A_183_141#_M1046_g N_X_c_1916_n 0.0101772f $X=24.305 $Y=2.965 $X2=0
+ $Y2=0
cc_878 N_A_183_141#_M1050_g N_X_c_1916_n 0.0101772f $X=25.085 $Y=2.965 $X2=0
+ $Y2=0
cc_879 N_A_183_141#_M1054_g N_X_c_1916_n 0.0101772f $X=25.865 $Y=2.965 $X2=0
+ $Y2=0
cc_880 N_A_183_141#_M1055_g N_X_c_1916_n 0.0101772f $X=26.645 $Y=2.965 $X2=0
+ $Y2=0
cc_881 N_A_183_141#_M1059_g N_X_c_1916_n 0.0101772f $X=27.425 $Y=2.965 $X2=0
+ $Y2=0
cc_882 N_A_183_141#_M1060_g N_X_c_1916_n 0.0101772f $X=28.205 $Y=2.965 $X2=0
+ $Y2=0
cc_883 N_A_183_141#_M1063_g N_X_c_1916_n 0.0101772f $X=28.985 $Y=2.965 $X2=0
+ $Y2=0
cc_884 N_A_183_141#_M1065_g N_X_c_1916_n 0.0101772f $X=29.765 $Y=2.965 $X2=0
+ $Y2=0
cc_885 N_A_183_141#_M1066_g N_X_c_1916_n 0.0101772f $X=30.545 $Y=2.965 $X2=0
+ $Y2=0
cc_886 N_A_183_141#_M1073_g N_X_c_1916_n 0.0101772f $X=31.325 $Y=2.965 $X2=0
+ $Y2=0
cc_887 N_A_183_141#_M1075_g N_X_c_1916_n 0.0148001f $X=32.105 $Y=2.965 $X2=0
+ $Y2=0
cc_888 N_A_183_141#_c_684_n N_X_c_1916_n 0.00241498f $X=10.035 $Y=1.665 $X2=0
+ $Y2=0
cc_889 N_A_183_141#_c_685_n N_X_c_1916_n 0.00241498f $X=11.595 $Y=1.665 $X2=0
+ $Y2=0
cc_890 N_A_183_141#_c_686_n N_X_c_1916_n 0.00241498f $X=13.155 $Y=1.665 $X2=0
+ $Y2=0
cc_891 N_A_183_141#_c_687_n N_X_c_1916_n 0.00241498f $X=14.715 $Y=1.665 $X2=0
+ $Y2=0
cc_892 N_A_183_141#_c_688_n N_X_c_1916_n 0.00241498f $X=16.275 $Y=1.665 $X2=0
+ $Y2=0
cc_893 N_A_183_141#_c_689_n N_X_c_1916_n 0.00241498f $X=17.835 $Y=1.665 $X2=0
+ $Y2=0
cc_894 N_A_183_141#_c_690_n N_X_c_1916_n 0.00241498f $X=19.395 $Y=1.665 $X2=0
+ $Y2=0
cc_895 N_A_183_141#_c_691_n N_X_c_1916_n 0.00497485f $X=20.945 $Y=1.665 $X2=0
+ $Y2=0
cc_896 N_A_183_141#_c_692_n N_X_c_1916_n 0.00241498f $X=22.515 $Y=1.665 $X2=0
+ $Y2=0
cc_897 N_A_183_141#_c_693_n N_X_c_1916_n 0.00241498f $X=24.075 $Y=1.665 $X2=0
+ $Y2=0
cc_898 N_A_183_141#_c_694_n N_X_c_1916_n 0.00241498f $X=25.635 $Y=1.665 $X2=0
+ $Y2=0
cc_899 N_A_183_141#_c_695_n N_X_c_1916_n 0.00241498f $X=27.195 $Y=1.665 $X2=0
+ $Y2=0
cc_900 N_A_183_141#_c_696_n N_X_c_1916_n 0.00241498f $X=28.755 $Y=1.665 $X2=0
+ $Y2=0
cc_901 N_A_183_141#_c_697_n N_X_c_1916_n 0.00241498f $X=30.315 $Y=1.665 $X2=0
+ $Y2=0
cc_902 N_A_183_141#_c_698_n N_X_c_1916_n 1.03594f $X=31.875 $Y=1.665 $X2=0 $Y2=0
cc_903 N_A_183_141#_c_699_n N_X_c_1916_n 0.00241498f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_904 N_A_183_141#_c_826_n N_VGND_M1012_d 0.00329714f $X=2.4 $Y=1.302 $X2=0
+ $Y2=0
cc_905 N_A_183_141#_c_841_n N_VGND_M1028_d 0.00329714f $X=4.025 $Y=1.302 $X2=0
+ $Y2=0
cc_906 N_A_183_141#_c_865_n N_VGND_M1043_d 0.00180843f $X=5.91 $Y=1.73 $X2=0
+ $Y2=0
cc_907 N_A_183_141#_c_860_n N_VGND_M1069_d 0.00181294f $X=7.06 $Y=1.73 $X2=-0.33
+ $Y2=-0.265
cc_908 N_A_183_141#_c_678_n N_VGND_c_2075_n 0.0344333f $X=1.055 $Y=0.92 $X2=0
+ $Y2=0
cc_909 N_A_183_141#_c_830_n N_VGND_c_2075_n 0.0177838f $X=1.17 $Y=1.302 $X2=0
+ $Y2=0
cc_910 N_A_183_141#_c_826_n N_VGND_c_2077_n 0.058686f $X=2.4 $Y=1.302 $X2=0
+ $Y2=0
cc_911 N_A_183_141#_c_679_n N_VGND_c_2077_n 0.0237236f $X=2.615 $Y=0.895 $X2=0
+ $Y2=0
cc_912 N_A_183_141#_c_679_n N_VGND_c_2079_n 0.0237236f $X=2.615 $Y=0.895 $X2=0
+ $Y2=0
cc_913 N_A_183_141#_c_841_n N_VGND_c_2079_n 0.0589786f $X=4.025 $Y=1.302 $X2=0
+ $Y2=0
cc_914 N_A_183_141#_c_680_n N_VGND_c_2079_n 0.0229431f $X=4.175 $Y=0.895 $X2=0
+ $Y2=0
cc_915 N_A_183_141#_c_849_n N_VGND_c_2081_n 0.0267967f $X=4.8 $Y=1.302 $X2=0
+ $Y2=0
cc_916 N_A_183_141#_c_681_n N_VGND_c_2081_n 0.0217012f $X=5.735 $Y=0.895 $X2=0
+ $Y2=0
cc_917 N_A_183_141#_c_865_n N_VGND_c_2081_n 0.033745f $X=5.91 $Y=1.73 $X2=0
+ $Y2=0
cc_918 N_A_183_141#_c_698_n N_VGND_c_2081_n 0.00142827f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_919 N_A_183_141#_c_681_n N_VGND_c_2083_n 0.0237236f $X=5.735 $Y=0.895 $X2=0
+ $Y2=0
cc_920 N_A_183_141#_c_860_n N_VGND_c_2083_n 0.0619717f $X=7.06 $Y=1.73 $X2=0
+ $Y2=0
cc_921 N_A_183_141#_c_682_n N_VGND_c_2083_n 0.0229431f $X=7.295 $Y=0.895 $X2=0
+ $Y2=0
cc_922 N_A_183_141#_c_698_n N_VGND_c_2083_n 0.00344444f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_923 N_A_183_141#_c_614_n N_VGND_c_2085_n 0.00109327f $X=8.705 $Y=1.565 $X2=0
+ $Y2=0
cc_924 N_A_183_141#_c_616_n N_VGND_c_2085_n 0.0475663f $X=9.485 $Y=1.565 $X2=0
+ $Y2=0
cc_925 N_A_183_141#_c_618_n N_VGND_c_2085_n 0.0474425f $X=10.265 $Y=1.565 $X2=0
+ $Y2=0
cc_926 N_A_183_141#_c_620_n N_VGND_c_2085_n 6.39245e-19 $X=11.045 $Y=1.565 $X2=0
+ $Y2=0
cc_927 N_A_183_141#_c_676_n N_VGND_c_2085_n 7.87968e-19 $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_928 N_A_183_141#_c_684_n N_VGND_c_2085_n 0.0413475f $X=10.035 $Y=1.665 $X2=0
+ $Y2=0
cc_929 N_A_183_141#_c_698_n N_VGND_c_2085_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_930 N_A_183_141#_c_618_n N_VGND_c_2087_n 6.39245e-19 $X=10.265 $Y=1.565 $X2=0
+ $Y2=0
cc_931 N_A_183_141#_c_620_n N_VGND_c_2087_n 0.0472746f $X=11.045 $Y=1.565 $X2=0
+ $Y2=0
cc_932 N_A_183_141#_c_622_n N_VGND_c_2087_n 0.0474425f $X=11.825 $Y=1.565 $X2=0
+ $Y2=0
cc_933 N_A_183_141#_c_624_n N_VGND_c_2087_n 6.39245e-19 $X=12.605 $Y=1.565 $X2=0
+ $Y2=0
cc_934 N_A_183_141#_c_676_n N_VGND_c_2087_n 7.87968e-19 $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_935 N_A_183_141#_c_685_n N_VGND_c_2087_n 0.0413475f $X=11.595 $Y=1.665 $X2=0
+ $Y2=0
cc_936 N_A_183_141#_c_698_n N_VGND_c_2087_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_937 N_A_183_141#_c_622_n N_VGND_c_2089_n 6.39245e-19 $X=11.825 $Y=1.565 $X2=0
+ $Y2=0
cc_938 N_A_183_141#_c_624_n N_VGND_c_2089_n 0.0472746f $X=12.605 $Y=1.565 $X2=0
+ $Y2=0
cc_939 N_A_183_141#_c_626_n N_VGND_c_2089_n 0.0474425f $X=13.385 $Y=1.565 $X2=0
+ $Y2=0
cc_940 N_A_183_141#_c_628_n N_VGND_c_2089_n 6.39245e-19 $X=14.165 $Y=1.565 $X2=0
+ $Y2=0
cc_941 N_A_183_141#_c_676_n N_VGND_c_2089_n 7.87968e-19 $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_942 N_A_183_141#_c_686_n N_VGND_c_2089_n 0.0413475f $X=13.155 $Y=1.665 $X2=0
+ $Y2=0
cc_943 N_A_183_141#_c_698_n N_VGND_c_2089_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_944 N_A_183_141#_c_626_n N_VGND_c_2091_n 6.39245e-19 $X=13.385 $Y=1.565 $X2=0
+ $Y2=0
cc_945 N_A_183_141#_c_628_n N_VGND_c_2091_n 0.0472746f $X=14.165 $Y=1.565 $X2=0
+ $Y2=0
cc_946 N_A_183_141#_c_630_n N_VGND_c_2091_n 0.0474425f $X=14.945 $Y=1.565 $X2=0
+ $Y2=0
cc_947 N_A_183_141#_c_632_n N_VGND_c_2091_n 6.39245e-19 $X=15.725 $Y=1.565 $X2=0
+ $Y2=0
cc_948 N_A_183_141#_c_676_n N_VGND_c_2091_n 7.87968e-19 $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_949 N_A_183_141#_c_687_n N_VGND_c_2091_n 0.0413475f $X=14.715 $Y=1.665 $X2=0
+ $Y2=0
cc_950 N_A_183_141#_c_698_n N_VGND_c_2091_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_951 N_A_183_141#_c_630_n N_VGND_c_2093_n 6.39245e-19 $X=14.945 $Y=1.565 $X2=0
+ $Y2=0
cc_952 N_A_183_141#_c_632_n N_VGND_c_2093_n 0.0472746f $X=15.725 $Y=1.565 $X2=0
+ $Y2=0
cc_953 N_A_183_141#_c_634_n N_VGND_c_2093_n 0.0474425f $X=16.505 $Y=1.565 $X2=0
+ $Y2=0
cc_954 N_A_183_141#_c_636_n N_VGND_c_2093_n 6.39245e-19 $X=17.285 $Y=1.565 $X2=0
+ $Y2=0
cc_955 N_A_183_141#_c_676_n N_VGND_c_2093_n 7.87968e-19 $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_956 N_A_183_141#_c_688_n N_VGND_c_2093_n 0.0413475f $X=16.275 $Y=1.665 $X2=0
+ $Y2=0
cc_957 N_A_183_141#_c_698_n N_VGND_c_2093_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_958 N_A_183_141#_c_634_n N_VGND_c_2095_n 6.39245e-19 $X=16.505 $Y=1.565 $X2=0
+ $Y2=0
cc_959 N_A_183_141#_c_636_n N_VGND_c_2095_n 0.0472746f $X=17.285 $Y=1.565 $X2=0
+ $Y2=0
cc_960 N_A_183_141#_c_638_n N_VGND_c_2095_n 0.0474425f $X=18.065 $Y=1.565 $X2=0
+ $Y2=0
cc_961 N_A_183_141#_c_640_n N_VGND_c_2095_n 6.39245e-19 $X=18.845 $Y=1.565 $X2=0
+ $Y2=0
cc_962 N_A_183_141#_c_676_n N_VGND_c_2095_n 7.87968e-19 $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_963 N_A_183_141#_c_689_n N_VGND_c_2095_n 0.0413475f $X=17.835 $Y=1.665 $X2=0
+ $Y2=0
cc_964 N_A_183_141#_c_698_n N_VGND_c_2095_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_965 N_A_183_141#_c_638_n N_VGND_c_2097_n 6.39245e-19 $X=18.065 $Y=1.565 $X2=0
+ $Y2=0
cc_966 N_A_183_141#_c_640_n N_VGND_c_2097_n 0.0472746f $X=18.845 $Y=1.565 $X2=0
+ $Y2=0
cc_967 N_A_183_141#_c_642_n N_VGND_c_2097_n 0.0477342f $X=19.625 $Y=1.565 $X2=0
+ $Y2=0
cc_968 N_A_183_141#_c_644_n N_VGND_c_2097_n 0.00109327f $X=20.405 $Y=1.565 $X2=0
+ $Y2=0
cc_969 N_A_183_141#_c_676_n N_VGND_c_2097_n 7.87968e-19 $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_970 N_A_183_141#_c_690_n N_VGND_c_2097_n 0.0413475f $X=19.395 $Y=1.665 $X2=0
+ $Y2=0
cc_971 N_A_183_141#_c_698_n N_VGND_c_2097_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_972 N_A_183_141#_c_642_n N_VGND_c_2099_n 9.4454e-19 $X=19.625 $Y=1.565 $X2=0
+ $Y2=0
cc_973 N_A_183_141#_c_644_n N_VGND_c_2099_n 0.0385917f $X=20.405 $Y=1.565 $X2=0
+ $Y2=0
cc_974 N_A_183_141#_c_646_n N_VGND_c_2099_n 0.0279616f $X=21.185 $Y=1.565 $X2=0
+ $Y2=0
cc_975 N_A_183_141#_c_676_n N_VGND_c_2099_n 7.87968e-19 $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_976 N_A_183_141#_c_691_n N_VGND_c_2099_n 0.0319273f $X=20.945 $Y=1.665 $X2=0
+ $Y2=0
cc_977 N_A_183_141#_c_698_n N_VGND_c_2099_n 0.0141551f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_978 N_A_183_141#_c_646_n N_VGND_c_2101_n 0.00109327f $X=21.185 $Y=1.565 $X2=0
+ $Y2=0
cc_979 N_A_183_141#_c_648_n N_VGND_c_2101_n 0.0475663f $X=21.965 $Y=1.565 $X2=0
+ $Y2=0
cc_980 N_A_183_141#_c_650_n N_VGND_c_2101_n 0.0474425f $X=22.745 $Y=1.565 $X2=0
+ $Y2=0
cc_981 N_A_183_141#_c_652_n N_VGND_c_2101_n 6.39245e-19 $X=23.525 $Y=1.565 $X2=0
+ $Y2=0
cc_982 N_A_183_141#_c_676_n N_VGND_c_2101_n 7.87968e-19 $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_983 N_A_183_141#_c_692_n N_VGND_c_2101_n 0.0413475f $X=22.515 $Y=1.665 $X2=0
+ $Y2=0
cc_984 N_A_183_141#_c_698_n N_VGND_c_2101_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_985 N_A_183_141#_c_650_n N_VGND_c_2103_n 6.39245e-19 $X=22.745 $Y=1.565 $X2=0
+ $Y2=0
cc_986 N_A_183_141#_c_652_n N_VGND_c_2103_n 0.0472746f $X=23.525 $Y=1.565 $X2=0
+ $Y2=0
cc_987 N_A_183_141#_c_654_n N_VGND_c_2103_n 0.0474425f $X=24.305 $Y=1.565 $X2=0
+ $Y2=0
cc_988 N_A_183_141#_c_656_n N_VGND_c_2103_n 6.39245e-19 $X=25.085 $Y=1.565 $X2=0
+ $Y2=0
cc_989 N_A_183_141#_c_676_n N_VGND_c_2103_n 7.87968e-19 $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_990 N_A_183_141#_c_693_n N_VGND_c_2103_n 0.0413475f $X=24.075 $Y=1.665 $X2=0
+ $Y2=0
cc_991 N_A_183_141#_c_698_n N_VGND_c_2103_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_992 N_A_183_141#_c_654_n N_VGND_c_2105_n 6.39245e-19 $X=24.305 $Y=1.565 $X2=0
+ $Y2=0
cc_993 N_A_183_141#_c_656_n N_VGND_c_2105_n 0.0472746f $X=25.085 $Y=1.565 $X2=0
+ $Y2=0
cc_994 N_A_183_141#_c_658_n N_VGND_c_2105_n 0.0474425f $X=25.865 $Y=1.565 $X2=0
+ $Y2=0
cc_995 N_A_183_141#_c_660_n N_VGND_c_2105_n 6.39245e-19 $X=26.645 $Y=1.565 $X2=0
+ $Y2=0
cc_996 N_A_183_141#_c_676_n N_VGND_c_2105_n 7.87968e-19 $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_997 N_A_183_141#_c_694_n N_VGND_c_2105_n 0.0413475f $X=25.635 $Y=1.665 $X2=0
+ $Y2=0
cc_998 N_A_183_141#_c_698_n N_VGND_c_2105_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_999 N_A_183_141#_c_658_n N_VGND_c_2107_n 6.39245e-19 $X=25.865 $Y=1.565 $X2=0
+ $Y2=0
cc_1000 N_A_183_141#_c_660_n N_VGND_c_2107_n 0.0472746f $X=26.645 $Y=1.565 $X2=0
+ $Y2=0
cc_1001 N_A_183_141#_c_662_n N_VGND_c_2107_n 0.0474425f $X=27.425 $Y=1.565 $X2=0
+ $Y2=0
cc_1002 N_A_183_141#_c_664_n N_VGND_c_2107_n 6.39245e-19 $X=28.205 $Y=1.565
+ $X2=0 $Y2=0
cc_1003 N_A_183_141#_c_676_n N_VGND_c_2107_n 7.87968e-19 $X=32.885 $Y=1.565
+ $X2=0 $Y2=0
cc_1004 N_A_183_141#_c_695_n N_VGND_c_2107_n 0.0413475f $X=27.195 $Y=1.665 $X2=0
+ $Y2=0
cc_1005 N_A_183_141#_c_698_n N_VGND_c_2107_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_1006 N_A_183_141#_c_662_n N_VGND_c_2109_n 6.39245e-19 $X=27.425 $Y=1.565
+ $X2=0 $Y2=0
cc_1007 N_A_183_141#_c_664_n N_VGND_c_2109_n 0.0472746f $X=28.205 $Y=1.565 $X2=0
+ $Y2=0
cc_1008 N_A_183_141#_c_666_n N_VGND_c_2109_n 0.0474425f $X=28.985 $Y=1.565 $X2=0
+ $Y2=0
cc_1009 N_A_183_141#_c_668_n N_VGND_c_2109_n 6.39245e-19 $X=29.765 $Y=1.565
+ $X2=0 $Y2=0
cc_1010 N_A_183_141#_c_676_n N_VGND_c_2109_n 7.87968e-19 $X=32.885 $Y=1.565
+ $X2=0 $Y2=0
cc_1011 N_A_183_141#_c_696_n N_VGND_c_2109_n 0.0413475f $X=28.755 $Y=1.665 $X2=0
+ $Y2=0
cc_1012 N_A_183_141#_c_698_n N_VGND_c_2109_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_1013 N_A_183_141#_c_666_n N_VGND_c_2111_n 6.39245e-19 $X=28.985 $Y=1.565
+ $X2=0 $Y2=0
cc_1014 N_A_183_141#_c_668_n N_VGND_c_2111_n 0.0472746f $X=29.765 $Y=1.565 $X2=0
+ $Y2=0
cc_1015 N_A_183_141#_c_670_n N_VGND_c_2111_n 0.0474425f $X=30.545 $Y=1.565 $X2=0
+ $Y2=0
cc_1016 N_A_183_141#_c_672_n N_VGND_c_2111_n 6.39245e-19 $X=31.325 $Y=1.565
+ $X2=0 $Y2=0
cc_1017 N_A_183_141#_c_676_n N_VGND_c_2111_n 7.87968e-19 $X=32.885 $Y=1.565
+ $X2=0 $Y2=0
cc_1018 N_A_183_141#_c_697_n N_VGND_c_2111_n 0.0413475f $X=30.315 $Y=1.665 $X2=0
+ $Y2=0
cc_1019 N_A_183_141#_c_698_n N_VGND_c_2111_n 0.0281234f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_1020 N_A_183_141#_c_670_n N_VGND_c_2113_n 6.39245e-19 $X=30.545 $Y=1.565
+ $X2=0 $Y2=0
cc_1021 N_A_183_141#_c_672_n N_VGND_c_2113_n 0.0472746f $X=31.325 $Y=1.565 $X2=0
+ $Y2=0
cc_1022 N_A_183_141#_c_674_n N_VGND_c_2113_n 0.05007f $X=32.105 $Y=1.565 $X2=0
+ $Y2=0
cc_1023 N_A_183_141#_c_676_n N_VGND_c_2113_n 0.00188124f $X=32.885 $Y=1.565
+ $X2=0 $Y2=0
cc_1024 N_A_183_141#_c_698_n N_VGND_c_2113_n 0.0248195f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_1025 N_A_183_141#_c_699_n N_VGND_c_2113_n 0.0413475f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_1026 N_A_183_141#_c_674_n N_VGND_c_2115_n 0.00109203f $X=32.105 $Y=1.565
+ $X2=0 $Y2=0
cc_1027 N_A_183_141#_c_676_n N_VGND_c_2115_n 0.0488451f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_1028 N_A_183_141#_c_614_n N_VGND_c_2117_n 0.0276587f $X=8.705 $Y=1.565 $X2=0
+ $Y2=0
cc_1029 N_A_183_141#_c_616_n N_VGND_c_2117_n 0.0109642f $X=9.485 $Y=1.565 $X2=0
+ $Y2=0
cc_1030 N_A_183_141#_c_618_n N_VGND_c_2117_n 0.0109642f $X=10.265 $Y=1.565 $X2=0
+ $Y2=0
cc_1031 N_A_183_141#_c_620_n N_VGND_c_2117_n 0.0109642f $X=11.045 $Y=1.565 $X2=0
+ $Y2=0
cc_1032 N_A_183_141#_c_622_n N_VGND_c_2117_n 0.0109642f $X=11.825 $Y=1.565 $X2=0
+ $Y2=0
cc_1033 N_A_183_141#_c_624_n N_VGND_c_2117_n 0.0109642f $X=12.605 $Y=1.565 $X2=0
+ $Y2=0
cc_1034 N_A_183_141#_c_626_n N_VGND_c_2117_n 0.0109642f $X=13.385 $Y=1.565 $X2=0
+ $Y2=0
cc_1035 N_A_183_141#_c_628_n N_VGND_c_2117_n 0.0109642f $X=14.165 $Y=1.565 $X2=0
+ $Y2=0
cc_1036 N_A_183_141#_c_630_n N_VGND_c_2117_n 0.0109642f $X=14.945 $Y=1.565 $X2=0
+ $Y2=0
cc_1037 N_A_183_141#_c_632_n N_VGND_c_2117_n 0.0109642f $X=15.725 $Y=1.565 $X2=0
+ $Y2=0
cc_1038 N_A_183_141#_c_634_n N_VGND_c_2117_n 0.0109642f $X=16.505 $Y=1.565 $X2=0
+ $Y2=0
cc_1039 N_A_183_141#_c_636_n N_VGND_c_2117_n 0.0109642f $X=17.285 $Y=1.565 $X2=0
+ $Y2=0
cc_1040 N_A_183_141#_c_638_n N_VGND_c_2117_n 0.0109642f $X=18.065 $Y=1.565 $X2=0
+ $Y2=0
cc_1041 N_A_183_141#_c_640_n N_VGND_c_2117_n 0.0109642f $X=18.845 $Y=1.565 $X2=0
+ $Y2=0
cc_1042 N_A_183_141#_c_642_n N_VGND_c_2117_n 0.0109642f $X=19.625 $Y=1.565 $X2=0
+ $Y2=0
cc_1043 N_A_183_141#_c_644_n N_VGND_c_2117_n 0.0129321f $X=20.405 $Y=1.565 $X2=0
+ $Y2=0
cc_1044 N_A_183_141#_c_646_n N_VGND_c_2117_n 0.0277186f $X=21.185 $Y=1.565 $X2=0
+ $Y2=0
cc_1045 N_A_183_141#_c_648_n N_VGND_c_2117_n 0.0109642f $X=21.965 $Y=1.565 $X2=0
+ $Y2=0
cc_1046 N_A_183_141#_c_650_n N_VGND_c_2117_n 0.0109642f $X=22.745 $Y=1.565 $X2=0
+ $Y2=0
cc_1047 N_A_183_141#_c_652_n N_VGND_c_2117_n 0.0109642f $X=23.525 $Y=1.565 $X2=0
+ $Y2=0
cc_1048 N_A_183_141#_c_654_n N_VGND_c_2117_n 0.0109642f $X=24.305 $Y=1.565 $X2=0
+ $Y2=0
cc_1049 N_A_183_141#_c_656_n N_VGND_c_2117_n 0.0109642f $X=25.085 $Y=1.565 $X2=0
+ $Y2=0
cc_1050 N_A_183_141#_c_658_n N_VGND_c_2117_n 0.0109642f $X=25.865 $Y=1.565 $X2=0
+ $Y2=0
cc_1051 N_A_183_141#_c_660_n N_VGND_c_2117_n 0.0109642f $X=26.645 $Y=1.565 $X2=0
+ $Y2=0
cc_1052 N_A_183_141#_c_662_n N_VGND_c_2117_n 0.0109642f $X=27.425 $Y=1.565 $X2=0
+ $Y2=0
cc_1053 N_A_183_141#_c_664_n N_VGND_c_2117_n 0.0109642f $X=28.205 $Y=1.565 $X2=0
+ $Y2=0
cc_1054 N_A_183_141#_c_666_n N_VGND_c_2117_n 0.0109642f $X=28.985 $Y=1.565 $X2=0
+ $Y2=0
cc_1055 N_A_183_141#_c_668_n N_VGND_c_2117_n 0.0109642f $X=29.765 $Y=1.565 $X2=0
+ $Y2=0
cc_1056 N_A_183_141#_c_670_n N_VGND_c_2117_n 0.0109642f $X=30.545 $Y=1.565 $X2=0
+ $Y2=0
cc_1057 N_A_183_141#_c_672_n N_VGND_c_2117_n 0.0109642f $X=31.325 $Y=1.565 $X2=0
+ $Y2=0
cc_1058 N_A_183_141#_c_674_n N_VGND_c_2117_n 0.0109642f $X=32.105 $Y=1.565 $X2=0
+ $Y2=0
cc_1059 N_A_183_141#_c_676_n N_VGND_c_2117_n 0.0129321f $X=32.885 $Y=1.565 $X2=0
+ $Y2=0
cc_1060 N_A_183_141#_c_678_n N_VGND_c_2117_n 0.0140143f $X=1.055 $Y=0.92 $X2=0
+ $Y2=0
cc_1061 N_A_183_141#_c_826_n N_VGND_c_2117_n 0.0124959f $X=2.4 $Y=1.302 $X2=0
+ $Y2=0
cc_1062 N_A_183_141#_c_679_n N_VGND_c_2117_n 0.0157921f $X=2.615 $Y=0.895 $X2=0
+ $Y2=0
cc_1063 N_A_183_141#_c_841_n N_VGND_c_2117_n 0.0123648f $X=4.025 $Y=1.302 $X2=0
+ $Y2=0
cc_1064 N_A_183_141#_c_680_n N_VGND_c_2117_n 0.0102287f $X=4.175 $Y=0.895 $X2=0
+ $Y2=0
cc_1065 N_A_183_141#_c_849_n N_VGND_c_2117_n 0.00615439f $X=4.8 $Y=1.302 $X2=0
+ $Y2=0
cc_1066 N_A_183_141#_c_681_n N_VGND_c_2117_n 0.0154229f $X=5.735 $Y=0.895 $X2=0
+ $Y2=0
cc_1067 N_A_183_141#_c_860_n N_VGND_c_2117_n 0.0058903f $X=7.06 $Y=1.73 $X2=0
+ $Y2=0
cc_1068 N_A_183_141#_c_865_n N_VGND_c_2117_n 0.0134192f $X=5.91 $Y=1.73 $X2=0
+ $Y2=0
cc_1069 N_A_183_141#_c_682_n N_VGND_c_2117_n 0.0102287f $X=7.295 $Y=0.895 $X2=0
+ $Y2=0
cc_1070 N_A_183_141#_c_683_n N_VGND_c_2117_n 0.00347419f $X=7.265 $Y=1.665 $X2=0
+ $Y2=0
cc_1071 N_A_183_141#_c_614_n N_VGND_c_2119_n 0.0359409f $X=8.705 $Y=1.565 $X2=0
+ $Y2=0
cc_1072 N_A_183_141#_c_698_n N_VGND_c_2119_n 0.0477715f $X=31.875 $Y=1.665 $X2=0
+ $Y2=0
cc_1073 N_VPWR_c_1421_n N_X_c_1741_n 0.0463441f $X=8.315 $Y=2.34 $X2=0 $Y2=0
cc_1074 N_VPWR_c_1423_n N_X_c_1741_n 0.117967f $X=9.875 $Y=2.34 $X2=0 $Y2=0
cc_1075 N_VPWR_c_1471_n N_X_c_1741_n 0.0415524f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1076 N_VPWR_c_1423_n N_X_c_1744_n 0.117967f $X=9.875 $Y=2.34 $X2=0 $Y2=0
cc_1077 N_VPWR_c_1426_n N_X_c_1744_n 0.117967f $X=11.435 $Y=2.34 $X2=0 $Y2=0
cc_1078 N_VPWR_c_1471_n N_X_c_1744_n 0.037804f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1079 N_VPWR_c_1426_n N_X_c_1747_n 0.117967f $X=11.435 $Y=2.34 $X2=0 $Y2=0
cc_1080 N_VPWR_c_1429_n N_X_c_1747_n 0.117967f $X=12.995 $Y=2.34 $X2=0 $Y2=0
cc_1081 N_VPWR_c_1471_n N_X_c_1747_n 0.037804f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1082 N_VPWR_c_1429_n N_X_c_1750_n 0.117967f $X=12.995 $Y=2.34 $X2=0 $Y2=0
cc_1083 N_VPWR_c_1432_n N_X_c_1750_n 0.117967f $X=14.555 $Y=2.34 $X2=0 $Y2=0
cc_1084 N_VPWR_c_1471_n N_X_c_1750_n 0.037804f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1085 N_VPWR_c_1432_n N_X_c_1753_n 0.117967f $X=14.555 $Y=2.34 $X2=0 $Y2=0
cc_1086 N_VPWR_c_1435_n N_X_c_1753_n 0.117967f $X=16.115 $Y=2.34 $X2=0 $Y2=0
cc_1087 N_VPWR_c_1471_n N_X_c_1753_n 0.037804f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1088 N_VPWR_c_1435_n N_X_c_1756_n 0.117967f $X=16.115 $Y=2.34 $X2=0 $Y2=0
cc_1089 N_VPWR_c_1438_n N_X_c_1756_n 0.117967f $X=17.675 $Y=2.34 $X2=0 $Y2=0
cc_1090 N_VPWR_c_1471_n N_X_c_1756_n 0.037804f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1091 N_VPWR_c_1438_n N_X_c_1759_n 0.117967f $X=17.675 $Y=2.34 $X2=0 $Y2=0
cc_1092 N_VPWR_c_1441_n N_X_c_1759_n 0.117967f $X=19.235 $Y=2.34 $X2=0 $Y2=0
cc_1093 N_VPWR_c_1471_n N_X_c_1759_n 0.037804f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1094 N_VPWR_c_1441_n N_X_c_1762_n 0.119317f $X=19.235 $Y=2.34 $X2=0 $Y2=0
cc_1095 N_VPWR_c_1444_n N_X_c_1762_n 0.117633f $X=20.795 $Y=2.36 $X2=0 $Y2=0
cc_1096 N_VPWR_c_1471_n N_X_c_1762_n 0.0456596f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1097 N_VPWR_c_1444_n N_X_c_1765_n 0.0469427f $X=20.795 $Y=2.36 $X2=0 $Y2=0
cc_1098 N_VPWR_c_1447_n N_X_c_1765_n 0.117967f $X=22.355 $Y=2.34 $X2=0 $Y2=0
cc_1099 N_VPWR_c_1471_n N_X_c_1765_n 0.0409539f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1100 N_VPWR_c_1447_n N_X_c_1768_n 0.117967f $X=22.355 $Y=2.34 $X2=0 $Y2=0
cc_1101 N_VPWR_c_1450_n N_X_c_1768_n 0.117967f $X=23.915 $Y=2.34 $X2=0 $Y2=0
cc_1102 N_VPWR_c_1471_n N_X_c_1768_n 0.037804f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1103 N_VPWR_c_1450_n N_X_c_1771_n 0.117967f $X=23.915 $Y=2.34 $X2=0 $Y2=0
cc_1104 N_VPWR_c_1453_n N_X_c_1771_n 0.117967f $X=25.475 $Y=2.34 $X2=0 $Y2=0
cc_1105 N_VPWR_c_1471_n N_X_c_1771_n 0.037804f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1106 N_VPWR_c_1453_n N_X_c_1774_n 0.117967f $X=25.475 $Y=2.34 $X2=0 $Y2=0
cc_1107 N_VPWR_c_1456_n N_X_c_1774_n 0.117967f $X=27.035 $Y=2.34 $X2=0 $Y2=0
cc_1108 N_VPWR_c_1471_n N_X_c_1774_n 0.037804f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1109 N_VPWR_c_1456_n N_X_c_1777_n 0.117967f $X=27.035 $Y=2.34 $X2=0 $Y2=0
cc_1110 N_VPWR_c_1459_n N_X_c_1777_n 0.117967f $X=28.595 $Y=2.34 $X2=0 $Y2=0
cc_1111 N_VPWR_c_1471_n N_X_c_1777_n 0.037804f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1112 N_VPWR_c_1459_n N_X_c_1780_n 0.117967f $X=28.595 $Y=2.34 $X2=0 $Y2=0
cc_1113 N_VPWR_c_1462_n N_X_c_1780_n 0.117967f $X=30.155 $Y=2.34 $X2=0 $Y2=0
cc_1114 N_VPWR_c_1471_n N_X_c_1780_n 0.037804f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1115 N_VPWR_c_1462_n N_X_c_1783_n 0.117967f $X=30.155 $Y=2.34 $X2=0 $Y2=0
cc_1116 N_VPWR_c_1465_n N_X_c_1783_n 0.117967f $X=31.715 $Y=2.34 $X2=0 $Y2=0
cc_1117 N_VPWR_c_1471_n N_X_c_1783_n 0.037804f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1118 N_VPWR_c_1465_n N_X_c_1786_n 0.119317f $X=31.715 $Y=2.34 $X2=0 $Y2=0
cc_1119 N_VPWR_c_1468_n N_X_c_1786_n 0.119397f $X=33.275 $Y=2.36 $X2=0 $Y2=0
cc_1120 N_VPWR_c_1471_n N_X_c_1786_n 0.0456596f $X=33.355 $Y=3.56 $X2=0 $Y2=0
cc_1121 N_VPWR_c_1421_n N_X_c_1916_n 0.00152661f $X=8.315 $Y=2.34 $X2=0 $Y2=0
cc_1122 N_VPWR_c_1423_n N_X_c_1916_n 0.0919982f $X=9.875 $Y=2.34 $X2=0 $Y2=0
cc_1123 N_VPWR_c_1426_n N_X_c_1916_n 0.0919982f $X=11.435 $Y=2.34 $X2=0 $Y2=0
cc_1124 N_VPWR_c_1429_n N_X_c_1916_n 0.0919982f $X=12.995 $Y=2.34 $X2=0 $Y2=0
cc_1125 N_VPWR_c_1432_n N_X_c_1916_n 0.0919982f $X=14.555 $Y=2.34 $X2=0 $Y2=0
cc_1126 N_VPWR_c_1435_n N_X_c_1916_n 0.0919982f $X=16.115 $Y=2.34 $X2=0 $Y2=0
cc_1127 N_VPWR_c_1438_n N_X_c_1916_n 0.0919982f $X=17.675 $Y=2.34 $X2=0 $Y2=0
cc_1128 N_VPWR_c_1441_n N_X_c_1916_n 0.0919982f $X=19.235 $Y=2.34 $X2=0 $Y2=0
cc_1129 N_VPWR_c_1444_n N_X_c_1916_n 0.0584837f $X=20.795 $Y=2.36 $X2=0 $Y2=0
cc_1130 N_VPWR_c_1447_n N_X_c_1916_n 0.0919982f $X=22.355 $Y=2.34 $X2=0 $Y2=0
cc_1131 N_VPWR_c_1450_n N_X_c_1916_n 0.0919982f $X=23.915 $Y=2.34 $X2=0 $Y2=0
cc_1132 N_VPWR_c_1453_n N_X_c_1916_n 0.0919982f $X=25.475 $Y=2.34 $X2=0 $Y2=0
cc_1133 N_VPWR_c_1456_n N_X_c_1916_n 0.0919982f $X=27.035 $Y=2.34 $X2=0 $Y2=0
cc_1134 N_VPWR_c_1459_n N_X_c_1916_n 0.0919982f $X=28.595 $Y=2.34 $X2=0 $Y2=0
cc_1135 N_VPWR_c_1462_n N_X_c_1916_n 0.0919982f $X=30.155 $Y=2.34 $X2=0 $Y2=0
cc_1136 N_VPWR_c_1465_n N_X_c_1916_n 0.0938713f $X=31.715 $Y=2.34 $X2=0 $Y2=0
cc_1137 N_VPWR_c_1468_n N_X_c_1916_n 0.00133085f $X=33.275 $Y=2.36 $X2=0 $Y2=0
cc_1138 N_VPWR_c_1468_n N_VGND_c_2115_n 0.0166422f $X=33.275 $Y=2.36 $X2=0 $Y2=0
cc_1139 N_X_c_1741_n N_VGND_c_2085_n 0.0480657f $X=9.095 $Y=0.955 $X2=0 $Y2=0
cc_1140 N_X_c_1744_n N_VGND_c_2085_n 0.0480657f $X=10.655 $Y=0.955 $X2=0 $Y2=0
cc_1141 N_X_c_1744_n N_VGND_c_2087_n 0.0480657f $X=10.655 $Y=0.955 $X2=0 $Y2=0
cc_1142 N_X_c_1747_n N_VGND_c_2087_n 0.0480657f $X=12.215 $Y=0.955 $X2=0 $Y2=0
cc_1143 N_X_c_1747_n N_VGND_c_2089_n 0.0480657f $X=12.215 $Y=0.955 $X2=0 $Y2=0
cc_1144 N_X_c_1750_n N_VGND_c_2089_n 0.0480657f $X=13.775 $Y=0.955 $X2=0 $Y2=0
cc_1145 N_X_c_1750_n N_VGND_c_2091_n 0.0480657f $X=13.775 $Y=0.955 $X2=0 $Y2=0
cc_1146 N_X_c_1753_n N_VGND_c_2091_n 0.0480657f $X=15.335 $Y=0.955 $X2=0 $Y2=0
cc_1147 N_X_c_1753_n N_VGND_c_2093_n 0.0480657f $X=15.335 $Y=0.955 $X2=0 $Y2=0
cc_1148 N_X_c_1756_n N_VGND_c_2093_n 0.0480657f $X=16.895 $Y=0.955 $X2=0 $Y2=0
cc_1149 N_X_c_1756_n N_VGND_c_2095_n 0.0480657f $X=16.895 $Y=0.955 $X2=0 $Y2=0
cc_1150 N_X_c_1759_n N_VGND_c_2095_n 0.0480657f $X=18.455 $Y=0.955 $X2=0 $Y2=0
cc_1151 N_X_c_1759_n N_VGND_c_2097_n 0.0480657f $X=18.455 $Y=0.955 $X2=0 $Y2=0
cc_1152 N_X_c_1762_n N_VGND_c_2097_n 0.0488323f $X=20.015 $Y=0.955 $X2=0 $Y2=0
cc_1153 N_X_c_1762_n N_VGND_c_2099_n 0.0478744f $X=20.015 $Y=0.955 $X2=0 $Y2=0
cc_1154 N_X_c_1765_n N_VGND_c_2099_n 0.0214076f $X=21.575 $Y=0.955 $X2=0 $Y2=0
cc_1155 N_X_c_1765_n N_VGND_c_2101_n 0.0480657f $X=21.575 $Y=0.955 $X2=0 $Y2=0
cc_1156 N_X_c_1768_n N_VGND_c_2101_n 0.0480657f $X=23.135 $Y=0.955 $X2=0 $Y2=0
cc_1157 N_X_c_1768_n N_VGND_c_2103_n 0.0480657f $X=23.135 $Y=0.955 $X2=0 $Y2=0
cc_1158 N_X_c_1771_n N_VGND_c_2103_n 0.0480657f $X=24.695 $Y=0.955 $X2=0 $Y2=0
cc_1159 N_X_c_1771_n N_VGND_c_2105_n 0.0480657f $X=24.695 $Y=0.955 $X2=0 $Y2=0
cc_1160 N_X_c_1774_n N_VGND_c_2105_n 0.0480657f $X=26.255 $Y=0.955 $X2=0 $Y2=0
cc_1161 N_X_c_1774_n N_VGND_c_2107_n 0.0480657f $X=26.255 $Y=0.955 $X2=0 $Y2=0
cc_1162 N_X_c_1777_n N_VGND_c_2107_n 0.0480657f $X=27.815 $Y=0.955 $X2=0 $Y2=0
cc_1163 N_X_c_1777_n N_VGND_c_2109_n 0.0480657f $X=27.815 $Y=0.955 $X2=0 $Y2=0
cc_1164 N_X_c_1780_n N_VGND_c_2109_n 0.0480657f $X=29.375 $Y=0.955 $X2=0 $Y2=0
cc_1165 N_X_c_1780_n N_VGND_c_2111_n 0.0480657f $X=29.375 $Y=0.955 $X2=0 $Y2=0
cc_1166 N_X_c_1783_n N_VGND_c_2111_n 0.0480657f $X=30.935 $Y=0.955 $X2=0 $Y2=0
cc_1167 N_X_c_1783_n N_VGND_c_2113_n 0.0480657f $X=30.935 $Y=0.955 $X2=0 $Y2=0
cc_1168 N_X_c_1786_n N_VGND_c_2113_n 0.0488323f $X=32.495 $Y=0.955 $X2=0 $Y2=0
cc_1169 N_X_c_1786_n N_VGND_c_2115_n 0.0557875f $X=32.495 $Y=0.955 $X2=0 $Y2=0
cc_1170 N_X_c_1741_n N_VGND_c_2117_n 0.0184011f $X=9.095 $Y=0.955 $X2=0 $Y2=0
cc_1171 N_X_c_1744_n N_VGND_c_2117_n 0.0184011f $X=10.655 $Y=0.955 $X2=0 $Y2=0
cc_1172 N_X_c_1747_n N_VGND_c_2117_n 0.0184011f $X=12.215 $Y=0.955 $X2=0 $Y2=0
cc_1173 N_X_c_1750_n N_VGND_c_2117_n 0.0184011f $X=13.775 $Y=0.955 $X2=0 $Y2=0
cc_1174 N_X_c_1753_n N_VGND_c_2117_n 0.0184011f $X=15.335 $Y=0.955 $X2=0 $Y2=0
cc_1175 N_X_c_1756_n N_VGND_c_2117_n 0.0184011f $X=16.895 $Y=0.955 $X2=0 $Y2=0
cc_1176 N_X_c_1759_n N_VGND_c_2117_n 0.0184011f $X=18.455 $Y=0.955 $X2=0 $Y2=0
cc_1177 N_X_c_1762_n N_VGND_c_2117_n 0.0223691f $X=20.015 $Y=0.955 $X2=0 $Y2=0
cc_1178 N_X_c_1765_n N_VGND_c_2117_n 0.0184011f $X=21.575 $Y=0.955 $X2=0 $Y2=0
cc_1179 N_X_c_1768_n N_VGND_c_2117_n 0.0184011f $X=23.135 $Y=0.955 $X2=0 $Y2=0
cc_1180 N_X_c_1771_n N_VGND_c_2117_n 0.0184011f $X=24.695 $Y=0.955 $X2=0 $Y2=0
cc_1181 N_X_c_1774_n N_VGND_c_2117_n 0.0184011f $X=26.255 $Y=0.955 $X2=0 $Y2=0
cc_1182 N_X_c_1777_n N_VGND_c_2117_n 0.0184011f $X=27.815 $Y=0.955 $X2=0 $Y2=0
cc_1183 N_X_c_1780_n N_VGND_c_2117_n 0.0184011f $X=29.375 $Y=0.955 $X2=0 $Y2=0
cc_1184 N_X_c_1783_n N_VGND_c_2117_n 0.0184011f $X=30.935 $Y=0.955 $X2=0 $Y2=0
cc_1185 N_X_c_1786_n N_VGND_c_2117_n 0.0223691f $X=32.495 $Y=0.955 $X2=0 $Y2=0
cc_1186 N_X_c_1741_n N_VGND_c_2119_n 0.0218845f $X=9.095 $Y=0.955 $X2=0 $Y2=0
