* File: sky130_fd_sc_hvl__dfstp_1.spice
* Created: Wed Sep  2 09:05:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__dfstp_1.pex.spice"
.subckt sky130_fd_sc_hvl__dfstp_1  VNB VPB CLK D SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_CLK_M1017_g N_A_30_131#_M1017_s N_VNB_M1017_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1029 N_A_340_593#_M1029_d N_A_30_131#_M1029_g N_VGND_M1017_d N_VNB_M1017_b NHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1027 N_A_642_107#_M1027_d N_D_M1027_g N_VGND_M1027_s N_VNB_M1017_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1006 N_A_798_107#_M1006_d N_A_30_131#_M1006_g N_A_642_107#_M1027_d
+ N_VNB_M1017_b NHV L=0.5 W=0.42 AD=0.063 AS=0.0588 PD=0.72 PS=0.7 NRD=5.4264
+ NRS=0 M=1 R=0.84 SA=250001 SB=250002 A=0.21 P=1.84 MULT=1
MM1023 A_958_107# N_A_340_593#_M1023_g N_A_798_107#_M1006_d N_VNB_M1017_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.063 PD=0.63 PS=0.72 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1003 N_VGND_M1003_d N_A_1000_81#_M1003_g A_958_107# N_VNB_M1017_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1025 A_1268_251# N_A_798_107#_M1025_g N_A_1000_81#_M1025_s N_VNB_M1017_b NHV
+ L=0.5 W=0.42 AD=0.1419 AS=0.1113 PD=1.17 PS=1.37 NRD=76.7676 NRS=0 M=1 R=0.84
+ SA=250000 SB=250003 A=0.21 P=1.84 MULT=1
MM1022 N_VGND_M1022_d N_SET_B_M1022_g A_1268_251# N_VNB_M1017_b NHV L=0.5 W=0.42
+ AD=0.0879308 AS=0.1419 PD=0.807692 PS=1.17 NRD=25.7754 NRS=76.7676 M=1 R=0.84
+ SA=250001 SB=250005 A=0.21 P=1.84 MULT=1
MM1013 A_1645_137# N_A_798_107#_M1013_g N_VGND_M1022_d N_VNB_M1017_b NHV L=0.5
+ W=0.75 AD=0.07875 AS=0.157019 PD=0.96 PS=1.44231 NRD=7.5924 NRS=0 M=1 R=1.5
+ SA=250001 SB=250003 A=0.375 P=2.5 MULT=1
MM1015 N_A_1787_137#_M1015_d N_A_340_593#_M1015_g A_1645_137# N_VNB_M1017_b NHV
+ L=0.5 W=0.75 AD=0.190192 AS=0.07875 PD=1.61538 PS=0.96 NRD=17.4762 NRS=7.5924
+ M=1 R=1.5 SA=250002 SB=250002 A=0.375 P=2.5 MULT=1
MM1018 A_1989_203# N_A_30_131#_M1018_g N_A_1787_137#_M1015_d N_VNB_M1017_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.106508 PD=0.63 PS=0.904615 NRD=13.566 NRS=31.2132
+ M=1 R=0.84 SA=250003 SB=250002 A=0.21 P=1.84 MULT=1
MM1019 A_2131_203# N_A_2031_177#_M1019_g A_1989_203# N_VNB_M1017_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=13.566 NRS=13.566 M=1 R=0.84
+ SA=250004 SB=250002 A=0.21 P=1.84 MULT=1
MM1020 N_VGND_M1020_d N_SET_B_M1020_g A_2131_203# N_VNB_M1017_b NHV L=0.5 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250005
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1007 N_A_2031_177#_M1007_d N_A_1787_137#_M1007_g N_VGND_M1020_d N_VNB_M1017_b
+ NHV L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250005 SB=250000 A=0.21 P=1.84 MULT=1
MM1004 N_VGND_M1004_d N_A_1787_137#_M1004_g N_A_2553_203#_M1004_s N_VNB_M1017_b
+ NHV L=0.5 W=0.42 AD=0.0933154 AS=0.1197 PD=0.822051 PS=1.41 NRD=31.2132 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1008 N_Q_M1008_d N_A_2553_203#_M1008_g N_VGND_M1004_d N_VNB_M1017_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.166635 PD=2.07 PS=1.46795 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1016 N_VPWR_M1016_d N_CLK_M1016_g N_A_30_131#_M1016_s N_VPB_M1016_b PHV L=0.5
+ W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1028 N_A_340_593#_M1028_d N_A_30_131#_M1028_g N_VPWR_M1016_d N_VPB_M1016_b PHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1002 N_A_642_107#_M1002_d N_D_M1002_g N_VPWR_M1002_s N_VPB_M1016_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.2247 PD=0.7 PS=1.91 NRD=0 NRS=122.775 M=1 R=0.84
+ SA=250000 SB=250008 A=0.21 P=1.84 MULT=1
MM1024 N_A_798_107#_M1024_d N_A_340_593#_M1024_g N_A_642_107#_M1002_d
+ N_VPB_M1016_b PHV L=0.5 W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=0 NRS=0
+ M=1 R=0.84 SA=250001 SB=250007 A=0.21 P=1.84 MULT=1
MM1021 A_982_529# N_A_30_131#_M1021_g N_A_798_107#_M1024_d N_VPB_M1016_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=22.729 NRS=18.1832 M=1
+ R=0.84 SA=250002 SB=250006 A=0.21 P=1.84 MULT=1
MM1000 N_VPWR_M1000_d N_A_1000_81#_M1000_g A_982_529# N_VPB_M1016_b PHV L=0.5
+ W=0.42 AD=0.0987 AS=0.0441 PD=0.89 PS=0.63 NRD=4.5458 NRS=22.729 M=1 R=0.84
+ SA=250003 SB=250005 A=0.21 P=1.84 MULT=1
MM1009 N_A_1000_81#_M1009_d N_A_798_107#_M1009_g N_VPWR_M1000_d N_VPB_M1016_b
+ PHV L=0.5 W=0.42 AD=0.0588 AS=0.0987 PD=0.7 PS=0.89 NRD=0 NRS=81.8435 M=1
+ R=0.84 SA=250004 SB=250004 A=0.21 P=1.84 MULT=1
MM1026 N_VPWR_M1026_d N_SET_B_M1026_g N_A_1000_81#_M1009_d N_VPB_M1016_b PHV
+ L=0.5 W=0.42 AD=0.0979606 AS=0.0588 PD=0.825211 PS=0.7 NRD=53.4227 NRS=0 M=1
+ R=0.84 SA=250004 SB=250004 A=0.21 P=1.84 MULT=1
MM1011 A_1653_515# N_A_798_107#_M1011_g N_VPWR_M1026_d N_VPB_M1016_b PHV L=0.5
+ W=1 AD=0.105 AS=0.233239 PD=1.21 PS=1.96479 NRD=9.5309 NRS=0 M=1 R=2 SA=250002
+ SB=250002 A=0.5 P=3 MULT=1
MM1014 N_A_1787_137#_M1014_d N_A_30_131#_M1014_g A_1653_515# N_VPB_M1016_b PHV
+ L=0.5 W=1 AD=0.286056 AS=0.105 PD=2.07042 PS=1.21 NRD=18.145 NRS=9.5309 M=1
+ R=2 SA=250003 SB=250001 A=0.5 P=3 MULT=1
MM1030 A_1989_515# N_A_340_593#_M1030_g N_A_1787_137#_M1014_d N_VPB_M1016_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.120144 PD=0.63 PS=0.869577 NRD=22.729 NRS=105.069
+ M=1 R=0.84 SA=250006 SB=250002 A=0.21 P=1.84 MULT=1
MM1031 N_VPWR_M1031_d N_A_2031_177#_M1031_g A_1989_515# N_VPB_M1016_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250007 SB=250001 A=0.21 P=1.84 MULT=1
MM1010 N_A_1787_137#_M1010_d N_SET_B_M1010_g N_VPWR_M1031_d N_VPB_M1016_b PHV
+ L=0.5 W=0.42 AD=0.11585 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250008 SB=250000 A=0.21 P=1.84 MULT=1
MM1012 N_VPWR_M1012_d N_A_1787_137#_M1012_g N_A_2031_177#_M1012_s N_VPB_M1016_b
+ PHV L=0.5 W=0.42 AD=0.1113 AS=0.1848 PD=1.37 PS=1.72 NRD=0 NRS=70.479 M=1
+ R=0.84 SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1005 N_VPWR_M1005_d N_A_1787_137#_M1005_g N_A_2553_203#_M1005_s N_VPB_M1016_b
+ PHV L=0.5 W=0.75 AD=0.148929 AS=0.19875 PD=1.17857 PS=2.03 NRD=24.1806 NRS=0
+ M=1 R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1001 N_Q_M1001_d N_A_2553_203#_M1001_g N_VPWR_M1005_d N_VPB_M1016_b PHV L=0.5
+ W=1 AD=0.265 AS=0.198571 PD=2.53 PS=1.57143 NRD=0 NRS=0 M=1 R=2 SA=250001
+ SB=250000 A=0.5 P=3 MULT=1
DX32_noxref N_VNB_M1017_b N_VPB_M1016_b NWDIODE A=39.675 P=37
*
.include "sky130_fd_sc_hvl__dfstp_1.pxi.spice"
*
.ends
*
*
