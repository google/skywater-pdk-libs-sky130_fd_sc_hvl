* File: sky130_fd_sc_hvl__dlxtp_1.pex.spice
* Created: Wed Sep  2 09:06:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__DLXTP_1%VNB 5 7 11 25
r61 7 25 1.53186e-05 $w=8.16e-06 $l=1e-09 $layer=MET1_cond $X=4.08 $Y=0.057
+ $X2=4.08 $Y2=0.058
r62 7 11 0.000873162 $w=8.16e-06 $l=5.7e-08 $layer=MET1_cond $X=4.08 $Y=0.057
+ $X2=4.08 $Y2=0
r63 5 11 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r64 5 11 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__DLXTP_1%VPB 4 6 14 21
r75 10 21 0.000873162 $w=8.16e-06 $l=5.7e-08 $layer=MET1_cond $X=4.08 $Y=4.07
+ $X2=4.08 $Y2=4.013
r76 10 14 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=7.92 $Y=4.07
+ $X2=7.92 $Y2=4.07
r77 9 14 501.048 $w=1.68e-07 $l=7.68e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=7.92 $Y2=4.07
r78 9 10 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r79 6 21 1.53186e-05 $w=8.16e-06 $l=1e-09 $layer=MET1_cond $X=4.08 $Y=4.012
+ $X2=4.08 $Y2=4.013
r80 4 14 21.4118 $w=1.7e-07 $l=7.96239e-06 $layer=licon1_NTAP_notbjt $count=8
+ $X=0 $Y=3.985 $X2=7.92 $Y2=4.07
r81 4 9 21.4118 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=8
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__DLXTP_1%GATE 3 7 9 12
r30 12 15 42.2298 $w=7.25e-07 $l=5.25e-07 $layer=POLY_cond $X=0.777 $Y=1.28
+ $X2=0.777 $Y2=1.805
r31 12 14 18.8261 $w=7.25e-07 $l=1.95e-07 $layer=POLY_cond $X=0.777 $Y=1.28
+ $X2=0.777 $Y2=1.085
r32 9 12 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.705
+ $Y=1.28 $X2=0.705 $Y2=1.28
r33 7 14 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.89 $Y=0.745 $X2=0.89
+ $Y2=1.085
r34 3 15 83.9996 $w=5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.665 $Y=2.59
+ $X2=0.665 $Y2=1.805
.ends

.subckt PM_SKY130_FD_SC_HVL__DLXTP_1%A_30_443# 1 2 9 13 16 19 21 25 26 29 30 33
+ 34 35 36 37 38 42 48 50 51 54 58 61
c142 42 0 1.663e-19 $X=4.575 $Y=1.25
c143 38 0 1.10735e-19 $X=4.41 $Y=2.615
r144 54 58 74.9041 $w=5e-07 $l=7e-07 $layer=POLY_cond $X=3.925 $Y=2.61 $X2=3.925
+ $Y2=3.31
r145 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.885
+ $Y=2.61 $X2=3.885 $Y2=2.61
r146 45 48 6.33922 $w=4.98e-07 $l=2.65e-07 $layer=LI1_cond $X=0.235 $Y=0.745
+ $X2=0.5 $Y2=0.745
r147 43 61 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.56 $Y=1.25 $X2=4.56
+ $Y2=0.745
r148 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.575
+ $Y=1.25 $X2=4.575 $Y2=1.25
r149 40 42 44.177 $w=3.28e-07 $l=1.265e-06 $layer=LI1_cond $X=4.575 $Y=2.515
+ $X2=4.575 $Y2=1.25
r150 39 53 3.28802 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=2.615
+ $X2=3.885 $Y2=2.615
r151 38 40 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=4.41 $Y=2.615
+ $X2=4.575 $Y2=2.515
r152 38 39 19.9636 $w=1.98e-07 $l=3.6e-07 $layer=LI1_cond $X=4.41 $Y=2.615
+ $X2=4.05 $Y2=2.615
r153 36 53 3.58693 $w=1.7e-07 $l=1.34164e-07 $layer=LI1_cond $X=3.965 $Y=2.715
+ $X2=3.885 $Y2=2.615
r154 36 37 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.965 $Y=2.715
+ $X2=3.965 $Y2=3.635
r155 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.88 $Y=3.72
+ $X2=3.965 $Y2=3.635
r156 34 35 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.88 $Y=3.72
+ $X2=3.19 $Y2=3.72
r157 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.105 $Y=3.635
+ $X2=3.19 $Y2=3.72
r158 32 33 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.105 $Y=2.815
+ $X2=3.105 $Y2=3.635
r159 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.02 $Y=2.73
+ $X2=3.105 $Y2=2.815
r160 30 31 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.02 $Y=2.73
+ $X2=1.78 $Y2=2.73
r161 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.695 $Y=2.645
+ $X2=1.78 $Y2=2.73
r162 28 51 4.27425 $w=2.12e-07 $l=2.35053e-07 $layer=LI1_cond $X=1.695 $Y=2.075
+ $X2=1.54 $Y2=1.905
r163 28 29 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.695 $Y=2.075
+ $X2=1.695 $Y2=2.645
r164 26 67 55.2893 $w=5.65e-07 $l=5.75e-07 $layer=POLY_cond $X=1.702 $Y=1.51
+ $X2=1.702 $Y2=2.085
r165 26 66 18.358 $w=5.65e-07 $l=1.85e-07 $layer=POLY_cond $X=1.702 $Y=1.51
+ $X2=1.702 $Y2=1.325
r166 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.705
+ $Y=1.51 $X2=1.705 $Y2=1.51
r167 23 51 4.27425 $w=2.12e-07 $l=1.27e-07 $layer=LI1_cond $X=1.667 $Y=1.905
+ $X2=1.54 $Y2=1.905
r168 23 25 17.8516 $w=2.53e-07 $l=3.95e-07 $layer=LI1_cond $X=1.667 $Y=1.905
+ $X2=1.667 $Y2=1.51
r169 22 50 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.36 $Y=1.99
+ $X2=0.235 $Y2=1.99
r170 21 51 2.15711 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=1.99
+ $X2=1.54 $Y2=1.905
r171 21 22 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=1.54 $Y=1.99
+ $X2=0.36 $Y2=1.99
r172 17 50 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=2.075
+ $X2=0.235 $Y2=1.99
r173 17 19 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=0.235 $Y=2.075
+ $X2=0.235 $Y2=2.36
r174 16 50 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=1.905
+ $X2=0.235 $Y2=1.99
r175 15 45 4.80115 $w=2.5e-07 $l=2.5e-07 $layer=LI1_cond $X=0.235 $Y=0.995
+ $X2=0.235 $Y2=0.745
r176 15 16 41.9489 $w=2.48e-07 $l=9.1e-07 $layer=LI1_cond $X=0.235 $Y=0.995
+ $X2=0.235 $Y2=1.905
r177 13 67 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.735 $Y=2.59
+ $X2=1.735 $Y2=2.085
r178 9 66 62.0634 $w=5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.67 $Y=0.745 $X2=1.67
+ $Y2=1.325
r179 2 19 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.215 $X2=0.275 $Y2=2.36
r180 1 48 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.355
+ $Y=0.535 $X2=0.5 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DLXTP_1%D 3 6 9 11 12 15 16
c48 16 0 3.56284e-20 $X=2.935 $Y=1.96
r49 15 17 18.3095 $w=5.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.035 $Y=1.96
+ $X2=3.035 $Y2=1.775
r50 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.935
+ $Y=1.96 $X2=2.935 $Y2=1.96
r51 12 16 5.26632 $w=6.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.64 $Y=2.13
+ $X2=2.935 $Y2=2.13
r52 9 11 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.07 $Y=3.31 $X2=3.07
+ $Y2=2.805
r53 6 11 27.696 $w=5.7e-07 $l=2.85e-07 $layer=POLY_cond $X=3.035 $Y=2.52
+ $X2=3.035 $Y2=2.805
r54 5 15 9.38648 $w=5.7e-07 $l=1e-07 $layer=POLY_cond $X=3.035 $Y=2.06 $X2=3.035
+ $Y2=1.96
r55 5 6 43.1778 $w=5.7e-07 $l=4.6e-07 $layer=POLY_cond $X=3.035 $Y=2.06
+ $X2=3.035 $Y2=2.52
r56 3 17 110.216 $w=5e-07 $l=1.03e-06 $layer=POLY_cond $X=3 $Y=0.745 $X2=3
+ $Y2=1.775
.ends

.subckt PM_SKY130_FD_SC_HVL__DLXTP_1%A_384_107# 1 2 9 12 13 14 15 17 22 26 31 32
+ 34 36 37
c98 14 0 1.46364e-19 $X=4.06 $Y=2.1
c99 13 0 1.5616e-19 $X=4.54 $Y=2.1
c100 9 0 1.663e-19 $X=3.78 $Y=0.745
r101 37 39 18.909 $w=5.3e-07 $l=1.85e-07 $layer=POLY_cond $X=3.795 $Y=1.545
+ $X2=3.795 $Y2=1.36
r102 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.715
+ $Y=1.545 $X2=3.715 $Y2=1.545
r103 31 32 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=2.125 $Y=2.37
+ $X2=2.125 $Y2=2.195
r104 27 34 3.22099 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.29 $Y=1.53
+ $X2=2.132 $Y2=1.53
r105 26 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=1.53
+ $X2=3.715 $Y2=1.53
r106 26 27 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=3.55 $Y=1.53
+ $X2=2.29 $Y2=1.53
r107 24 34 3.32435 $w=2.82e-07 $l=8.5e-08 $layer=LI1_cond $X=2.132 $Y=1.615
+ $X2=2.132 $Y2=1.53
r108 24 32 21.2196 $w=3.13e-07 $l=5.8e-07 $layer=LI1_cond $X=2.132 $Y=1.615
+ $X2=2.132 $Y2=2.195
r109 20 34 3.32435 $w=2.82e-07 $l=9.97246e-08 $layer=LI1_cond $X=2.1 $Y=1.445
+ $X2=2.132 $Y2=1.53
r110 20 22 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=2.1 $Y=1.445 $X2=2.1
+ $Y2=0.745
r111 15 19 65.2226 $w=5.21e-07 $l=7.12461e-07 $layer=POLY_cond $X=4.82 $Y=2.805
+ $X2=4.805 $Y2=2.1
r112 15 17 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.82 $Y=2.805 $X2=4.82
+ $Y2=3.145
r113 13 19 21.9195 $w=2.3e-07 $l=2.65e-07 $layer=POLY_cond $X=4.54 $Y=2.1
+ $X2=4.805 $Y2=2.1
r114 13 14 133.923 $w=2.3e-07 $l=4.8e-07 $layer=POLY_cond $X=4.54 $Y=2.1
+ $X2=4.06 $Y2=2.1
r115 12 14 32.7876 $w=2.3e-07 $l=3.17333e-07 $layer=POLY_cond $X=3.795 $Y=1.985
+ $X2=4.06 $Y2=2.1
r116 11 37 8.07592 $w=5.3e-07 $l=8e-08 $layer=POLY_cond $X=3.795 $Y=1.625
+ $X2=3.795 $Y2=1.545
r117 11 12 36.3416 $w=5.3e-07 $l=3.6e-07 $layer=POLY_cond $X=3.795 $Y=1.625
+ $X2=3.795 $Y2=1.985
r118 9 39 65.8086 $w=5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.78 $Y=0.745
+ $X2=3.78 $Y2=1.36
r119 2 31 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=2.215 $X2=2.125 $Y2=2.37
r120 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.535 $X2=2.06 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DLXTP_1%A_1004_81# 1 2 7 9 10 12 13 15 19 21 23 26
+ 29 30 35 39
c72 12 0 1.86045e-19 $X=5.595 $Y=1.23
r73 41 43 27.8215 $w=5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.27 $Y=1.315 $X2=5.53
+ $Y2=1.315
r74 36 43 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.53 $Y=1.565 $X2=5.53
+ $Y2=1.315
r75 30 33 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=6.19 $Y=2.27
+ $X2=6.19 $Y2=2.425
r76 29 39 168.534 $w=5e-07 $l=1.575e-06 $layer=POLY_cond $X=5.53 $Y=1.57
+ $X2=5.53 $Y2=3.145
r77 29 36 0.535029 $w=5e-07 $l=5e-09 $layer=POLY_cond $X=5.53 $Y=1.57 $X2=5.53
+ $Y2=1.565
r78 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.595
+ $Y=1.57 $X2=5.595 $Y2=1.57
r79 25 26 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.945 $Y=1.595
+ $X2=6.945 $Y2=2.185
r80 24 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.375 $Y=1.51
+ $X2=6.21 $Y2=1.51
r81 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.86 $Y=1.51
+ $X2=6.945 $Y2=1.595
r82 23 24 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=6.86 $Y=1.51
+ $X2=6.375 $Y2=1.51
r83 22 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.355 $Y=2.27
+ $X2=6.19 $Y2=2.27
r84 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.86 $Y=2.27
+ $X2=6.945 $Y2=2.185
r85 21 22 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=6.86 $Y=2.27
+ $X2=6.355 $Y2=2.27
r86 17 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.21 $Y=1.425
+ $X2=6.21 $Y2=1.51
r87 17 19 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=6.21 $Y=1.425
+ $X2=6.21 $Y2=1.075
r88 16 28 4.88517 $w=1.7e-07 $l=1.79374e-07 $layer=LI1_cond $X=5.76 $Y=1.51
+ $X2=5.595 $Y2=1.54
r89 15 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.045 $Y=1.51
+ $X2=6.21 $Y2=1.51
r90 15 16 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.045 $Y=1.51
+ $X2=5.76 $Y2=1.51
r91 13 43 6.95538 $w=5e-07 $l=6.5e-08 $layer=POLY_cond $X=5.595 $Y=1.315
+ $X2=5.53 $Y2=1.315
r92 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.595
+ $Y=1.23 $X2=5.595 $Y2=1.23
r93 10 28 2.881 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=5.595 $Y=1.425
+ $X2=5.595 $Y2=1.54
r94 10 12 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=5.595 $Y=1.425
+ $X2=5.595 $Y2=1.23
r95 7 41 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.27 $Y=1.065 $X2=5.27
+ $Y2=1.315
r96 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.27 $Y=1.065 $X2=5.27
+ $Y2=0.745
r97 2 33 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=6.045
+ $Y=2.215 $X2=6.19 $Y2=2.425
r98 1 19 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=6.085
+ $Y=0.865 $X2=6.21 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__DLXTP_1%A_806_107# 1 2 9 13 17 21 23 25 27 29 32 34
+ 38 44 46 48 53
c106 53 0 1.14976e-20 $X=7.475 $Y=1.75
c107 29 0 1.5616e-19 $X=4.92 $Y=2.98
c108 13 0 1.74548e-19 $X=6.6 $Y=1.075
r109 52 53 75.0445 $w=5.62e-07 $l=8.75e-07 $layer=POLY_cond $X=6.6 $Y=1.75
+ $X2=7.475 $Y2=1.75
r110 51 52 1.7153 $w=5.62e-07 $l=2e-08 $layer=POLY_cond $X=6.58 $Y=1.75 $X2=6.6
+ $Y2=1.75
r111 47 51 5.57473 $w=5.62e-07 $l=6.5e-08 $layer=POLY_cond $X=6.515 $Y=1.75
+ $X2=6.58 $Y2=1.75
r112 46 48 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.515 $Y=1.89
+ $X2=6.35 $Y2=1.89
r113 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.515
+ $Y=1.89 $X2=6.515 $Y2=1.89
r114 38 40 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=0.745
+ $X2=4.17 $Y2=0.83
r115 36 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.09 $Y=1.92
+ $X2=5.005 $Y2=1.92
r116 36 48 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=5.09 $Y=1.92
+ $X2=6.35 $Y2=1.92
r117 33 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=2.005
+ $X2=5.005 $Y2=1.92
r118 33 34 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=5.005 $Y=2.005
+ $X2=5.005 $Y2=2.895
r119 32 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=1.835
+ $X2=5.005 $Y2=1.92
r120 31 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.005 $Y=0.915
+ $X2=5.005 $Y2=1.835
r121 30 43 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.48 $Y=2.98
+ $X2=4.355 $Y2=2.98
r122 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.92 $Y=2.98
+ $X2=5.005 $Y2=2.895
r123 29 30 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=4.92 $Y=2.98
+ $X2=4.48 $Y2=2.98
r124 28 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=0.83
+ $X2=4.17 $Y2=0.83
r125 27 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.92 $Y=0.83
+ $X2=5.005 $Y2=0.915
r126 27 28 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.92 $Y=0.83
+ $X2=4.335 $Y2=0.83
r127 23 43 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.355 $Y=3.065
+ $X2=4.355 $Y2=2.98
r128 23 25 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=4.355 $Y=3.065
+ $X2=4.355 $Y2=3.56
r129 19 53 1.7153 $w=5.62e-07 $l=2e-08 $layer=POLY_cond $X=7.495 $Y=1.75
+ $X2=7.475 $Y2=1.75
r130 19 21 72.229 $w=5e-07 $l=6.75e-07 $layer=POLY_cond $X=7.495 $Y=1.585
+ $X2=7.495 $Y2=0.91
r131 15 53 5.60901 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=7.475 $Y=2.085
+ $X2=7.475 $Y2=1.75
r132 15 17 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=7.475 $Y=2.085
+ $X2=7.475 $Y2=2.965
r133 11 52 5.60901 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.6 $Y=1.415 $X2=6.6
+ $Y2=1.75
r134 11 13 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.6 $Y=1.415 $X2=6.6
+ $Y2=1.075
r135 7 51 5.60901 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.58 $Y=2.085
+ $X2=6.58 $Y2=1.75
r136 7 9 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.58 $Y=2.085 $X2=6.58
+ $Y2=2.425
r137 2 43 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.175
+ $Y=2.935 $X2=4.315 $Y2=3.06
r138 2 25 600 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=1 $X=4.175
+ $Y=2.935 $X2=4.315 $Y2=3.56
r139 1 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.535 $X2=4.17 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DLXTP_1%VPWR 1 2 3 4 13 16 31 35 44 51
r54 48 51 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=6.65 $Y=3.63
+ $X2=7.37 $Y2=3.63
r55 47 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.37 $Y=3.59
+ $X2=7.37 $Y2=3.59
r56 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.65 $Y=3.59
+ $X2=6.65 $Y2=3.59
r57 44 47 12.4568 $w=9.48e-07 $l=9.7e-07 $layer=LI1_cond $X=7.01 $Y=2.62
+ $X2=7.01 $Y2=3.59
r58 41 48 0.209228 $w=3.7e-07 $l=5.45e-07 $layer=MET1_cond $X=6.105 $Y=3.63
+ $X2=6.65 $Y2=3.63
r59 39 41 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.385 $Y=3.63
+ $X2=6.105 $Y2=3.63
r60 38 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.105 $Y=3.59
+ $X2=6.105 $Y2=3.59
r61 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.385 $Y=3.59
+ $X2=5.385 $Y2=3.59
r62 35 38 5.71474 $w=9.48e-07 $l=4.45e-07 $layer=LI1_cond $X=5.745 $Y=3.145
+ $X2=5.745 $Y2=3.59
r63 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.725 $Y=3.59
+ $X2=2.725 $Y2=3.59
r64 29 31 0.842309 $w=7.08e-07 $l=5e-08 $layer=LI1_cond $X=2.675 $Y=3.35
+ $X2=2.725 $Y2=3.35
r65 26 32 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.005 $Y=3.63
+ $X2=2.725 $Y2=3.63
r66 25 29 11.2869 $w=7.08e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=3.35
+ $X2=2.675 $Y2=3.35
r67 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.005 $Y=3.59
+ $X2=2.005 $Y2=3.59
r68 22 26 0.253378 $w=3.7e-07 $l=6.6e-07 $layer=MET1_cond $X=1.345 $Y=3.63
+ $X2=2.005 $Y2=3.63
r69 20 22 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.625 $Y=3.63
+ $X2=1.345 $Y2=3.63
r70 19 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.345 $Y=3.59
+ $X2=1.345 $Y2=3.59
r71 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.625 $Y=3.59
+ $X2=0.625 $Y2=3.59
r72 16 19 17.1348 $w=8.88e-07 $l=1.25e-06 $layer=LI1_cond $X=0.985 $Y=2.34
+ $X2=0.985 $Y2=3.59
r73 13 39 0.500997 $w=3.7e-07 $l=1.305e-06 $layer=MET1_cond $X=4.08 $Y=3.63
+ $X2=5.385 $Y2=3.63
r74 13 32 0.520192 $w=3.7e-07 $l=1.355e-06 $layer=MET1_cond $X=4.08 $Y=3.63
+ $X2=2.725 $Y2=3.63
r75 4 47 400 $w=1.7e-07 $l=1.49708e-06 $layer=licon1_PDIFF $count=1 $X=6.83
+ $Y=2.215 $X2=7.085 $Y2=3.59
r76 4 44 400 $w=1.7e-07 $l=5.17011e-07 $layer=licon1_PDIFF $count=1 $X=6.83
+ $Y=2.215 $X2=7.085 $Y2=2.62
r77 3 35 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.78
+ $Y=2.935 $X2=5.92 $Y2=3.145
r78 2 29 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.55
+ $Y=2.935 $X2=2.675 $Y2=3.08
r79 1 16 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.915
+ $Y=2.215 $X2=1.055 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__DLXTP_1%A_650_107# 1 2 7 9 13 15 17 18 19 22 24
r64 21 22 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=4.145 $Y=1.265
+ $X2=4.145 $Y2=2.165
r65 20 23 2.50919 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=1.18
+ $X2=3.39 $Y2=1.18
r66 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=1.18
+ $X2=4.145 $Y2=1.265
r67 19 20 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.06 $Y=1.18
+ $X2=3.555 $Y2=1.18
r68 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=2.25
+ $X2=4.145 $Y2=2.165
r69 17 18 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.06 $Y=2.25
+ $X2=3.54 $Y2=2.25
r70 13 24 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.535 $Y=3.06
+ $X2=3.535 $Y2=2.895
r71 13 15 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.535 $Y=3.06
+ $X2=3.535 $Y2=3.215
r72 11 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.455 $Y=2.335
+ $X2=3.54 $Y2=2.25
r73 11 24 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.455 $Y=2.335
+ $X2=3.455 $Y2=2.895
r74 7 23 14.0725 $w=3.3e-07 $l=3.5e-07 $layer=LI1_cond $X=3.39 $Y=0.83 $X2=3.39
+ $Y2=1.18
r75 7 9 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.39 $Y=0.83 $X2=3.39
+ $Y2=0.745
r76 2 15 600 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=2.935 $X2=3.535 $Y2=3.215
r77 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.25
+ $Y=0.535 $X2=3.39 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DLXTP_1%Q 1 2 7 8 12
r15 19 21 41.1587 $w=3.48e-07 $l=1.25e-06 $layer=LI1_cond $X=7.875 $Y=2.34
+ $X2=7.875 $Y2=3.59
r16 8 19 10.0427 $w=3.48e-07 $l=3.05e-07 $layer=LI1_cond $X=7.875 $Y=2.035
+ $X2=7.875 $Y2=2.34
r17 7 8 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=7.875 $Y=1.665
+ $X2=7.875 $Y2=2.035
r18 7 12 32.433 $w=3.48e-07 $l=9.85e-07 $layer=LI1_cond $X=7.875 $Y=1.665
+ $X2=7.875 $Y2=0.68
r19 2 21 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=7.725
+ $Y=2.215 $X2=7.865 $Y2=3.59
r20 2 19 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=7.725
+ $Y=2.215 $X2=7.865 $Y2=2.34
r21 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.745
+ $Y=0.535 $X2=7.885 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__DLXTP_1%VGND 1 2 3 4 13 16 25 32 39 43
r58 45 47 6.42105 $w=9.48e-07 $l=5e-07 $layer=LI1_cond $X=7.03 $Y=0.66 $X2=7.03
+ $Y2=1.16
r59 40 43 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=6.67 $Y=0.44
+ $X2=7.39 $Y2=0.44
r60 39 45 2.31158 $w=9.48e-07 $l=1.8e-07 $layer=LI1_cond $X=7.03 $Y=0.48
+ $X2=7.03 $Y2=0.66
r61 39 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.39 $Y=0.48
+ $X2=7.39 $Y2=0.48
r62 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.67 $Y=0.48
+ $X2=6.67 $Y2=0.48
r63 33 40 0.355112 $w=3.7e-07 $l=9.25e-07 $layer=MET1_cond $X=5.745 $Y=0.44
+ $X2=6.67 $Y2=0.44
r64 32 36 5.37222 $w=5.88e-07 $l=2.65e-07 $layer=LI1_cond $X=5.565 $Y=0.48
+ $X2=5.565 $Y2=0.745
r65 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.745 $Y=0.48
+ $X2=5.745 $Y2=0.48
r66 25 29 5.37222 $w=5.88e-07 $l=2.65e-07 $layer=LI1_cond $X=2.7 $Y=0.48 $X2=2.7
+ $Y2=0.745
r67 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.88 $Y=0.48
+ $X2=2.88 $Y2=0.48
r68 20 26 0.460686 $w=3.7e-07 $l=1.2e-06 $layer=MET1_cond $X=1.68 $Y=0.44
+ $X2=2.88 $Y2=0.44
r69 17 20 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0.44
+ $X2=1.68 $Y2=0.44
r70 16 22 3.40316 $w=9.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.32 $Y=0.48
+ $X2=1.32 $Y2=0.745
r71 16 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0.48
+ $X2=1.68 $Y2=0.48
r72 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.96 $Y=0.48
+ $X2=0.96 $Y2=0.48
r73 13 33 0.639202 $w=3.7e-07 $l=1.665e-06 $layer=MET1_cond $X=4.08 $Y=0.44
+ $X2=5.745 $Y2=0.44
r74 13 26 0.460686 $w=3.7e-07 $l=1.2e-06 $layer=MET1_cond $X=4.08 $Y=0.44
+ $X2=2.88 $Y2=0.44
r75 4 47 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=6.85
+ $Y=0.865 $X2=7.105 $Y2=1.16
r76 4 45 182 $w=1.7e-07 $l=3.42491e-07 $layer=licon1_NDIFF $count=1 $X=6.85
+ $Y=0.865 $X2=7.105 $Y2=0.66
r77 3 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.52
+ $Y=0.535 $X2=5.66 $Y2=0.745
r78 2 29 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.535 $X2=2.61 $Y2=0.745
r79 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.535 $X2=1.28 $Y2=0.745
.ends

