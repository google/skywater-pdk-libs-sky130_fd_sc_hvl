* File: sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1.pxi.spice
* Created: Fri Aug 28 09:37:35 2020
* 
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%VNB N_VNB_M1015_b VNB VNB
+ N_VNB_c_62_p VNB VNB PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%VNB
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%VPB N_VPB_X19_noxref_D1
+ N_VPB_M1008_b VPB N_VPB_c_88_n N_VPB_c_100_p N_VPB_c_89_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%VPB
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%LVPWR N_LVPWR_M1005_d
+ N_LVPWR_M1005_b N_LVPWR_c_178_p LVPWR N_LVPWR_c_175_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%LVPWR
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A N_A_c_226_n N_A_c_227_n
+ N_A_M1015_g N_A_M1005_g N_A_c_228_n A A N_A_c_230_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_573_897# N_A_573_897#_M1015_s
+ N_A_573_897#_M1005_s N_A_573_897#_c_258_n N_A_573_897#_c_259_n
+ N_A_573_897#_c_260_n N_A_573_897#_M1001_g N_A_573_897#_c_261_n
+ N_A_573_897#_M1016_g N_A_573_897#_M1017_g N_A_573_897#_c_262_n
+ N_A_573_897#_M1004_g N_A_573_897#_c_263_n N_A_573_897#_c_264_n
+ N_A_573_897#_c_265_n N_A_573_897#_c_266_n N_A_573_897#_c_281_n
+ N_A_573_897#_c_267_n N_A_573_897#_c_268_n N_A_573_897#_c_285_n
+ N_A_573_897#_c_301_n PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_573_897#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_772_151# N_A_772_151#_M1016_d
+ N_A_772_151#_M1017_d N_A_772_151#_c_340_n N_A_772_151#_M1000_g
+ N_A_772_151#_c_341_n N_A_772_151#_M1012_g N_A_772_151#_c_342_n
+ N_A_772_151#_c_343_n N_A_772_151#_c_344_n N_A_772_151#_c_352_n
+ N_A_772_151#_c_345_n N_A_772_151#_c_353_n N_A_772_151#_c_346_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_772_151#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_1400_777# N_A_1400_777#_M1010_s
+ N_A_1400_777#_M15_noxref_d N_A_1400_777#_M1008_g N_A_1400_777#_c_390_n
+ N_A_1400_777#_M1009_g N_A_1400_777#_c_394_n N_A_1400_777#_c_397_n
+ N_A_1400_777#_c_400_n N_A_1400_777#_c_429_p N_A_1400_777#_c_401_n
+ N_A_1400_777#_c_404_n PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_1400_777#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_816_1221# N_A_816_1221#_M1001_s
+ N_A_816_1221#_M1008_s N_A_816_1221#_M13_noxref_s N_A_816_1221#_M1009_s
+ N_A_816_1221#_c_460_n N_A_816_1221#_c_472_n N_A_816_1221#_M1013_g
+ N_A_816_1221#_c_461_n N_A_816_1221#_c_462_n N_A_816_1221#_M1011_g
+ N_A_816_1221#_M15_noxref_g N_A_816_1221#_c_479_n N_A_816_1221#_c_482_n
+ N_A_816_1221#_c_497_n N_A_816_1221#_c_464_n N_A_816_1221#_c_465_n
+ N_A_816_1221#_c_484_n N_A_816_1221#_c_486_n N_A_816_1221#_c_466_n
+ N_A_816_1221#_c_467_n N_A_816_1221#_c_468_n N_A_816_1221#_c_469_n
+ N_A_816_1221#_c_491_n N_A_816_1221#_c_493_n N_A_816_1221#_c_470_n
+ N_A_816_1221#_c_471_n PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_816_1221#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_1406_429# N_A_1406_429#_M1011_s
+ N_A_1406_429#_M1013_s N_A_1406_429#_c_569_n N_A_1406_429#_M1010_g
+ N_A_1406_429#_c_570_n N_A_1406_429#_M1018_g N_A_1406_429#_c_571_n
+ N_A_1406_429#_c_572_n N_A_1406_429#_c_582_n N_A_1406_429#_M17_noxref_g
+ N_A_1406_429#_M1014_g N_A_1406_429#_M1007_g N_A_1406_429#_M13_noxref_g
+ N_A_1406_429#_c_587_n N_A_1406_429#_c_575_n N_A_1406_429#_c_577_n
+ N_A_1406_429#_c_578_n N_A_1406_429#_c_579_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_1406_429#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%VPWR N_VPWR_M1008_d
+ N_VPWR_M13_noxref_d N_VPWR_M1013_d N_VPWR_M17_noxref_d VPWR VPWR
+ N_VPWR_c_670_n N_VPWR_c_672_n N_VPWR_c_675_n N_VPWR_c_668_n N_VPWR_c_683_n
+ N_VPWR_c_669_n PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%VPWR
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%X N_X_M1007_d N_X_M1014_d X X X X
+ X N_X_c_758_n X X PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%X
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%VGND N_VGND_M1001_d N_VGND_M1015_d
+ N_VGND_M1004_d N_VGND_M1000_s N_VGND_M1012_s N_VGND_M1011_d N_VGND_c_771_n
+ N_VGND_c_772_n N_VGND_c_774_n N_VGND_c_776_n N_VGND_c_778_n VGND VGND
+ N_VGND_c_780_n N_VGND_c_782_n N_VGND_c_783_n N_VGND_c_785_n N_VGND_c_786_n
+ N_VGND_c_787_n N_VGND_c_788_n N_VGND_c_790_n N_VGND_c_792_n N_VGND_c_794_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%VGND
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_1197_107# N_A_1197_107#_M1000_d
+ N_A_1197_107#_M1010_d N_A_1197_107#_M1018_d N_A_1197_107#_c_874_n
+ N_A_1197_107#_c_867_n N_A_1197_107#_c_877_n N_A_1197_107#_c_868_n
+ N_A_1197_107#_c_869_n N_A_1197_107#_c_871_n N_A_1197_107#_c_873_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_1197_107#
cc_1 N_VNB_M1015_b N_VPB_c_88_n 0.0021751f $X=-0.33 $Y=-0.265 $X2=0.24 $Y2=4.07
cc_2 N_VNB_M1015_b N_VPB_c_89_n 0.0836033f $X=-0.33 $Y=-0.265 $X2=10.8 $Y2=4.07
cc_3 N_VNB_M1015_b LVPWR 0.161501f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_4 N_VNB_M1015_b N_A_c_226_n 0.0315583f $X=-0.33 $Y=-0.265 $X2=0 $Y2=3.985
cc_5 N_VNB_M1015_b N_A_c_227_n 0.0215558f $X=-0.33 $Y=-0.265 $X2=10.56 $Y2=3.985
cc_6 N_VNB_M1015_b N_A_c_228_n 0.00851298f $X=-0.33 $Y=-0.265 $X2=-0.33
+ $Y2=1.885
cc_7 N_VNB_M1015_b A 0.0248803f $X=-0.33 $Y=-0.265 $X2=6.335 $Y2=2.465
cc_8 N_VNB_M1015_b N_A_c_230_n 0.0812462f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_M1015_b N_A_573_897#_c_258_n 0.0422114f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_10 N_VNB_M1015_b N_A_573_897#_c_259_n 0.0466102f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1015_b N_A_573_897#_c_260_n 0.041717f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1015_b N_A_573_897#_c_261_n 0.0223696f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1015_b N_A_573_897#_c_262_n 0.160696f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_M1015_b N_A_573_897#_c_263_n 0.0125974f $X=-0.33 $Y=-0.265 $X2=8.88
+ $Y2=4.07
cc_15 N_VNB_M1015_b N_A_573_897#_c_264_n 0.00411489f $X=-0.33 $Y=-0.265 $X2=10.8
+ $Y2=4.07
cc_16 N_VNB_M1015_b N_A_573_897#_c_265_n 0.164089f $X=-0.33 $Y=-0.265 $X2=10.8
+ $Y2=4.07
cc_17 N_VNB_M1015_b N_A_573_897#_c_266_n 0.035967f $X=-0.33 $Y=-0.265 $X2=10.8
+ $Y2=4.07
cc_18 N_VNB_M1015_b N_A_573_897#_c_267_n 0.00652689f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_19 N_VNB_M1015_b N_A_573_897#_c_268_n 0.0344484f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_20 N_VNB_M1015_b N_A_772_151#_c_340_n 0.0398058f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_21 N_VNB_M1015_b N_A_772_151#_c_341_n 0.129288f $X=-0.33 $Y=-0.265 $X2=-0.33
+ $Y2=1.885
cc_22 N_VNB_M1015_b N_A_772_151#_c_342_n 0.0244016f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_23 N_VNB_M1015_b N_A_772_151#_c_343_n 0.0185531f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_24 N_VNB_M1015_b N_A_772_151#_c_344_n 0.014445f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_25 N_VNB_M1015_b N_A_772_151#_c_345_n 0.0384012f $X=-0.33 $Y=-0.265 $X2=10.8
+ $Y2=4.07
cc_26 N_VNB_M1015_b N_A_772_151#_c_346_n 0.084631f $X=-0.33 $Y=-0.265 $X2=8.4
+ $Y2=4.07
cc_27 N_VNB_M1015_b N_A_1400_777#_c_390_n 0.0615692f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_28 N_VNB_M1015_b N_A_816_1221#_c_460_n 0.0390225f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_29 N_VNB_M1015_b N_A_816_1221#_c_461_n 0.00158704f $X=-0.33 $Y=-0.265 $X2=8.4
+ $Y2=4.07
cc_30 N_VNB_M1015_b N_A_816_1221#_c_462_n 0.0816521f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_31 VNB N_A_816_1221#_c_462_n 0.00181995f $X=5.52 $Y=8.08 $X2=0 $Y2=0
cc_32 N_VNB_M1015_b N_A_816_1221#_c_464_n 0.113503f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_33 N_VNB_M1015_b N_A_816_1221#_c_465_n 0.0134401f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_M1015_b N_A_816_1221#_c_466_n 0.00121379f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_35 N_VNB_M1015_b N_A_816_1221#_c_467_n 0.04975f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_36 N_VNB_M1015_b N_A_816_1221#_c_468_n 0.0287849f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_37 N_VNB_M1015_b N_A_816_1221#_c_469_n 3.65815e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_38 N_VNB_M1015_b N_A_816_1221#_c_470_n 0.0226463f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_39 N_VNB_M1015_b N_A_816_1221#_c_471_n 0.0767625f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_M1015_b N_A_1406_429#_c_569_n 0.0390089f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_41 N_VNB_M1015_b N_A_1406_429#_c_570_n 0.0412062f $X=-0.33 $Y=-0.265
+ $X2=-0.33 $Y2=1.885
cc_42 N_VNB_M1015_b N_A_1406_429#_c_571_n 0.0505781f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_M1015_b N_A_1406_429#_c_572_n 0.109193f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=3.955
cc_44 N_VNB_M1015_b N_A_1406_429#_M1007_g 0.0682348f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_45 VNB N_A_1406_429#_M1007_g 0.00161049f $X=5.52 $Y=8.08 $X2=0 $Y2=0
cc_46 N_VNB_M1015_b N_A_1406_429#_c_575_n 0.0365757f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_47 VNB N_A_1406_429#_c_575_n 7.98897e-19 $X=5.52 $Y=8.08 $X2=0 $Y2=0
cc_48 N_VNB_M1015_b N_A_1406_429#_c_577_n 0.00203039f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_49 N_VNB_M1015_b N_A_1406_429#_c_578_n 0.0377119f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_M1015_b N_A_1406_429#_c_579_n 3.1372e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_51 N_VNB_M1015_b N_VPWR_c_668_n 0.281259f $X=-0.33 $Y=-0.265 $X2=10.8
+ $Y2=4.07
cc_52 N_VNB_M1015_b N_VPWR_c_669_n 0.0985775f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_53 N_VNB_M1015_b X 0.0443485f $X=-0.33 $Y=-0.265 $X2=6.335 $Y2=2.465
cc_54 VNB X 7.98897e-19 $X=5.52 $Y=8.08 $X2=6.335 $Y2=2.465
cc_55 N_VNB_M1015_b X 0.0234434f $X=-0.33 $Y=-0.265 $X2=10.8 $Y2=4.07
cc_56 N_VNB_M1015_b N_VGND_c_771_n 0.00570671f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_57 N_VNB_M1015_b N_VGND_c_772_n 0.119953f $X=-0.33 $Y=-0.265 $X2=8.4 $Y2=4.07
cc_58 VNB N_VGND_c_772_n 0.00531562f $X=5.52 $Y=8.08 $X2=8.4 $Y2=4.07
cc_59 N_VNB_M1015_b N_VGND_c_774_n 0.0481389f $X=-0.33 $Y=-0.265 $X2=8.4
+ $Y2=4.07
cc_60 VNB N_VGND_c_774_n 0.00198821f $X=5.52 $Y=8.08 $X2=8.4 $Y2=4.07
cc_61 N_VNB_M1015_b N_VGND_c_776_n 0.118741f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_62 N_VNB_c_62_p N_VGND_c_776_n 0.00531562f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_63 N_VNB_M1015_b N_VGND_c_778_n 0.0481389f $X=-0.33 $Y=-0.265 $X2=8.88
+ $Y2=4.07
cc_64 N_VNB_c_62_p N_VGND_c_778_n 0.00198821f $X=0.24 $Y=0 $X2=8.88 $Y2=4.07
cc_65 N_VNB_M1015_b N_VGND_c_780_n 0.0262752f $X=-0.33 $Y=-0.265 $X2=5.52
+ $Y2=4.07
cc_66 N_VNB_c_62_p N_VGND_c_780_n 0.00102546f $X=0.24 $Y=0 $X2=5.52 $Y2=4.07
cc_67 N_VNB_M1015_b N_VGND_c_782_n 0.0685056f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_68 N_VNB_M1015_b N_VGND_c_783_n 0.0262752f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_69 N_VNB_c_62_p N_VGND_c_783_n 0.00102546f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_70 N_VNB_M1015_b N_VGND_c_785_n 0.0682032f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_71 N_VNB_M1015_b N_VGND_c_786_n 0.0461766f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_72 N_VNB_M1015_b N_VGND_c_787_n 0.0252816f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_73 N_VNB_M1015_b N_VGND_c_788_n 0.410759f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_74 N_VNB_c_62_p N_VGND_c_788_n 1.16909f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_75 N_VNB_M1015_b N_VGND_c_790_n 0.0294115f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_790_n 0.00159492f $X=5.52 $Y=8.08 $X2=0 $Y2=0
cc_77 N_VNB_M1015_b N_VGND_c_792_n 0.463924f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_792_n 1.17391f $X=5.52 $Y=8.08 $X2=0 $Y2=0
cc_79 N_VNB_M1015_b N_VGND_c_794_n 0.0167066f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_80 N_VNB_c_62_p N_VGND_c_794_n 8.02293e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_81 N_VNB_M1015_b N_A_1197_107#_c_867_n 0.00895108f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_82 N_VNB_M1015_b N_A_1197_107#_c_868_n 0.0260815f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_83 N_VNB_M1015_b N_A_1197_107#_c_869_n 0.118614f $X=-0.33 $Y=-0.265 $X2=8.4
+ $Y2=4.07
cc_84 N_VNB_c_62_p N_A_1197_107#_c_869_n 0.00533173f $X=0.24 $Y=0 $X2=8.4
+ $Y2=4.07
cc_85 N_VNB_M1015_b N_A_1197_107#_c_871_n 0.0265719f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_86 N_VNB_c_62_p N_A_1197_107#_c_871_n 0.00111205f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_87 N_VNB_M1015_b N_A_1197_107#_c_873_n 0.0611567f $X=-0.33 $Y=-0.265 $X2=10.8
+ $Y2=4.07
cc_88 N_VPB_c_89_n N_LVPWR_M1005_b 0.00792118f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_89 N_VPB_X19_noxref_D1 LVPWR 0.050189f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_90 N_VPB_M1008_b LVPWR 0.0292589f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_91 N_VPB_c_89_n N_LVPWR_c_175_n 0.0433246f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_92 N_VPB_c_89_n N_A_573_897#_c_264_n 0.0252548f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_93 N_VPB_M1008_b N_A_772_151#_c_341_n 0.0161105f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_94 N_VPB_M1008_b N_A_1400_777#_M1008_g 0.0174193f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_95 N_VPB_M1008_b N_A_1400_777#_c_390_n 0.0429404f $X=6.335 $Y=2.465 $X2=0
+ $Y2=8.025
cc_96 N_VPB_M1008_b N_A_1400_777#_M1009_g 0.0174383f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_97 N_VPB_M1008_b N_A_1400_777#_c_394_n 0.0129548f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_98 N_VPB_c_100_p N_A_1400_777#_c_394_n 0.0033354f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_99 N_VPB_c_89_n N_A_1400_777#_c_394_n 0.0369239f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_100 N_VPB_M1008_b N_A_1400_777#_c_397_n 0.129279f $X=6.335 $Y=2.465 $X2=10.8
+ $Y2=0
cc_101 N_VPB_c_100_p N_A_1400_777#_c_397_n 0.00781608f $X=10.8 $Y=4.07 $X2=10.8
+ $Y2=0
cc_102 N_VPB_c_89_n N_A_1400_777#_c_397_n 0.0193145f $X=10.8 $Y=4.07 $X2=10.8
+ $Y2=0
cc_103 N_VPB_M1008_b N_A_1400_777#_c_400_n 0.00473944f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_104 N_VPB_M1008_b N_A_1400_777#_c_401_n 0.0239584f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_105 N_VPB_c_100_p N_A_1400_777#_c_401_n 0.0164577f $X=10.8 $Y=4.07 $X2=0
+ $Y2=0
cc_106 N_VPB_c_89_n N_A_1400_777#_c_401_n 0.00298227f $X=10.8 $Y=4.07 $X2=0
+ $Y2=0
cc_107 N_VPB_M1008_b N_A_1400_777#_c_404_n 9.68666e-19 $X=6.335 $Y=2.465
+ $X2=0.24 $Y2=8.14
cc_108 N_VPB_M1008_b N_A_816_1221#_c_472_n 0.0205311f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_109 N_VPB_c_100_p N_A_816_1221#_c_472_n 0.00747379f $X=10.8 $Y=4.07 $X2=0
+ $Y2=0
cc_110 N_VPB_c_89_n N_A_816_1221#_c_472_n 0.0042972f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_111 N_VPB_M1008_b N_A_816_1221#_c_461_n 0.0172572f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_112 N_VPB_M1008_b N_A_816_1221#_M15_noxref_g 0.165672f $X=6.335 $Y=2.465
+ $X2=0.24 $Y2=8.14
cc_113 N_VPB_c_100_p N_A_816_1221#_M15_noxref_g 0.031589f $X=10.8 $Y=4.07
+ $X2=0.24 $Y2=8.14
cc_114 N_VPB_c_89_n N_A_816_1221#_M15_noxref_g 0.0170487f $X=10.8 $Y=4.07
+ $X2=0.24 $Y2=8.14
cc_115 N_VPB_M1008_b N_A_816_1221#_c_479_n 0.0272169f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_VPB_c_100_p N_A_816_1221#_c_479_n 0.0215907f $X=10.8 $Y=4.07 $X2=0
+ $Y2=0
cc_117 N_VPB_c_89_n N_A_816_1221#_c_479_n 0.00529755f $X=10.8 $Y=4.07 $X2=0
+ $Y2=0
cc_118 N_VPB_M1008_b N_A_816_1221#_c_482_n 0.015503f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_119 N_VPB_M1008_b N_A_816_1221#_c_464_n 0.0311141f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_VPB_M1008_b N_A_816_1221#_c_484_n 0.0598638f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_121 N_VPB_c_89_n N_A_816_1221#_c_484_n 0.0277375f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_122 N_VPB_M1008_b N_A_816_1221#_c_486_n 0.0359239f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_123 N_VPB_M1008_b N_A_816_1221#_c_466_n 0.0108404f $X=6.335 $Y=2.465 $X2=5.52
+ $Y2=8.14
cc_124 N_VPB_M1008_b N_A_816_1221#_c_469_n 0.0226421f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_VPB_c_100_p N_A_816_1221#_c_469_n 0.0158392f $X=10.8 $Y=4.07 $X2=0
+ $Y2=0
cc_126 N_VPB_c_89_n N_A_816_1221#_c_469_n 0.00101808f $X=10.8 $Y=4.07 $X2=0
+ $Y2=0
cc_127 N_VPB_M1008_b N_A_816_1221#_c_491_n 0.0140344f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_128 N_VPB_c_89_n N_A_816_1221#_c_491_n 0.00102452f $X=10.8 $Y=4.07 $X2=0
+ $Y2=0
cc_129 N_VPB_M1008_b N_A_816_1221#_c_493_n 7.08293e-19 $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_130 N_VPB_M1008_b N_A_1406_429#_c_571_n 0.0879205f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_131 N_VPB_M1008_b N_A_1406_429#_c_572_n 0.126927f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_132 N_VPB_M1008_b N_A_1406_429#_c_582_n 0.065776f $X=6.335 $Y=2.465 $X2=0.24
+ $Y2=0
cc_133 N_VPB_c_100_p N_A_1406_429#_c_582_n 0.0386846f $X=10.8 $Y=4.07 $X2=0.24
+ $Y2=0
cc_134 N_VPB_c_89_n N_A_1406_429#_c_582_n 0.0111068f $X=10.8 $Y=4.07 $X2=0.24
+ $Y2=0
cc_135 N_VPB_M1008_b N_A_1406_429#_M17_noxref_g 0.114482f $X=6.335 $Y=2.465
+ $X2=0 $Y2=0
cc_136 N_VPB_M1008_b N_A_1406_429#_M1014_g 0.0378065f $X=6.335 $Y=2.465 $X2=10.8
+ $Y2=0
cc_137 N_VPB_M1008_b N_A_1406_429#_c_587_n 0.0221842f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_138 N_VPB_c_100_p N_A_1406_429#_c_587_n 0.015847f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_139 N_VPB_c_89_n N_A_1406_429#_c_587_n 0.00100899f $X=10.8 $Y=4.07 $X2=0
+ $Y2=0
cc_140 N_VPB_M1008_b N_A_1406_429#_c_577_n 0.00203039f $X=6.335 $Y=2.465
+ $X2=5.52 $Y2=0.06
cc_141 N_VPB_M1008_b N_A_1406_429#_c_578_n 0.00832153f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_VPB_M1008_b N_A_1406_429#_c_579_n 3.1372e-19 $X=6.335 $Y=2.465 $X2=5.52
+ $Y2=8.08
cc_143 N_VPB_M1008_b N_VPWR_c_670_n 0.00511699f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_144 N_VPB_c_89_n N_VPWR_c_670_n 0.0033293f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_145 N_VPB_M1008_b N_VPWR_c_672_n 0.00888593f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_146 N_VPB_c_100_p N_VPWR_c_672_n 0.0130681f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_147 N_VPB_c_89_n N_VPWR_c_672_n 0.00251628f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_148 N_VPB_M1008_b N_VPWR_c_675_n 0.00453345f $X=6.335 $Y=2.465 $X2=10.8
+ $Y2=8.14
cc_149 N_VPB_c_100_p N_VPWR_c_675_n 0.0272989f $X=10.8 $Y=4.07 $X2=10.8 $Y2=8.14
cc_150 N_VPB_c_89_n N_VPWR_c_675_n 0.00212134f $X=10.8 $Y=4.07 $X2=10.8 $Y2=8.14
cc_151 N_VPB_X19_noxref_D1 N_VPWR_c_668_n 0.0565882f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_152 N_VPB_M1008_b N_VPWR_c_668_n 0.0536814f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_153 N_VPB_c_88_n N_VPWR_c_668_n 0.00613319f $X=0.24 $Y=4.07 $X2=0 $Y2=0
cc_154 N_VPB_c_100_p N_VPWR_c_668_n 0.0186198f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_155 N_VPB_c_89_n N_VPWR_c_668_n 1.16209f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_156 N_VPB_M1008_b N_VPWR_c_683_n 0.0194246f $X=6.335 $Y=2.465 $X2=5.52
+ $Y2=0.06
cc_157 N_VPB_c_100_p N_VPWR_c_683_n 0.0235561f $X=10.8 $Y=4.07 $X2=5.52 $Y2=0.06
cc_158 N_VPB_c_89_n N_VPWR_c_683_n 0.00207094f $X=10.8 $Y=4.07 $X2=5.52 $Y2=0.06
cc_159 N_VPB_X19_noxref_D1 N_VPWR_c_669_n 0.0336658f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_160 N_VPB_M1008_b N_VPWR_c_669_n 0.0365696f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_161 N_VPB_c_88_n N_VPWR_c_669_n 0.00613319f $X=0.24 $Y=4.07 $X2=0 $Y2=0
cc_162 N_VPB_c_100_p N_VPWR_c_669_n 0.0171788f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_163 N_VPB_c_89_n N_VPWR_c_669_n 1.15492f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_164 N_VPB_M1008_b X 0.0077824f $X=6.335 $Y=2.465 $X2=-0.33 $Y2=-0.265
cc_165 N_VPB_M1008_b N_X_c_758_n 0.0518911f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_166 N_VPB_c_100_p N_X_c_758_n 0.0158392f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_167 N_VPB_c_89_n N_X_c_758_n 0.00101808f $X=10.8 $Y=4.07 $X2=0 $Y2=0
cc_168 N_VPB_M1008_b X 0.00990693f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_169 N_LVPWR_M1005_b N_A_c_226_n 0.0176162f $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_170 N_LVPWR_M1005_b N_A_M1005_g 0.0225938f $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_171 N_LVPWR_c_178_p N_A_M1005_g 0.00135859f $X=3.57 $Y=2.33 $X2=0 $Y2=0
cc_172 LVPWR N_A_M1005_g 0.0109749f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_173 N_LVPWR_c_175_n N_A_M1005_g 0.00417272f $X=3.93 $Y=3.19 $X2=0 $Y2=0
cc_174 N_LVPWR_M1005_b N_A_c_228_n 6.60476e-19 $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_175 N_LVPWR_M1005_b N_A_c_230_n 0.00547003f $X=2.8 $Y=2.015 $X2=0.24 $Y2=0
cc_176 LVPWR N_A_573_897#_M1005_s 5.28909e-19 $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_177 N_LVPWR_M1005_b N_A_573_897#_M1017_g 0.0221724f $X=2.8 $Y=2.015 $X2=0.24
+ $Y2=0
cc_178 N_LVPWR_c_178_p N_A_573_897#_M1017_g 0.00208937f $X=3.57 $Y=2.33 $X2=0.24
+ $Y2=0
cc_179 LVPWR N_A_573_897#_M1017_g 0.00767826f $X=0.07 $Y=3.02 $X2=0.24 $Y2=0
cc_180 N_LVPWR_c_175_n N_A_573_897#_M1017_g 0.0112605f $X=3.93 $Y=3.19 $X2=0.24
+ $Y2=0
cc_181 N_LVPWR_M1005_b N_A_573_897#_c_263_n 0.00262762f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_182 N_LVPWR_c_178_p N_A_573_897#_c_263_n 0.00156473f $X=3.57 $Y=2.33 $X2=0
+ $Y2=0
cc_183 N_LVPWR_M1005_b N_A_573_897#_c_264_n 0.0500919f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_184 N_LVPWR_c_178_p N_A_573_897#_c_264_n 8.98083e-19 $X=3.57 $Y=2.33 $X2=0
+ $Y2=0
cc_185 LVPWR N_A_573_897#_c_264_n 0.0236806f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_186 N_LVPWR_c_175_n N_A_573_897#_c_264_n 0.0814701f $X=3.93 $Y=3.19 $X2=0
+ $Y2=0
cc_187 N_LVPWR_M1005_b N_A_573_897#_c_281_n 0.0232362f $X=2.8 $Y=2.015 $X2=5.52
+ $Y2=0.06
cc_188 N_LVPWR_c_178_p N_A_573_897#_c_281_n 0.00429663f $X=3.57 $Y=2.33 $X2=5.52
+ $Y2=0.06
cc_189 N_LVPWR_c_178_p N_A_573_897#_c_267_n 0.0229916f $X=3.57 $Y=2.33 $X2=5.52
+ $Y2=8.08
cc_190 N_LVPWR_M1005_b N_A_573_897#_c_268_n 0.0124783f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_191 N_LVPWR_M1005_b N_A_573_897#_c_285_n 0.016229f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_192 LVPWR N_A_573_897#_c_285_n 0.0263553f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_193 LVPWR N_A_772_151#_M1017_d 0.00288751f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_194 N_LVPWR_M1005_b N_A_772_151#_c_344_n 0.00801775f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_195 N_LVPWR_c_178_p N_A_772_151#_c_344_n 0.00252726f $X=3.57 $Y=2.33 $X2=0
+ $Y2=0
cc_196 LVPWR N_A_772_151#_c_344_n 0.0235018f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_197 LVPWR N_A_772_151#_c_352_n 0.0320105f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_198 N_LVPWR_M1005_b N_A_772_151#_c_353_n 0.016687f $X=2.8 $Y=2.015 $X2=10.8
+ $Y2=8.14
cc_199 LVPWR N_A_772_151#_c_353_n 0.0115771f $X=0.07 $Y=3.02 $X2=10.8 $Y2=8.14
cc_200 N_LVPWR_c_175_n N_A_772_151#_c_353_n 0.0160139f $X=3.93 $Y=3.19 $X2=10.8
+ $Y2=8.14
cc_201 LVPWR N_A_772_151#_c_346_n 0.0405719f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_202 LVPWR N_A_1400_777#_M15_noxref_d 0.0030514f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_203 LVPWR N_A_1400_777#_c_394_n 0.0713199f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_204 LVPWR N_A_1400_777#_c_400_n 0.00789846f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_205 LVPWR N_A_1400_777#_c_401_n 0.0940362f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_206 LVPWR N_A_816_1221#_M13_noxref_s 0.00604067f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_207 LVPWR N_A_816_1221#_M15_noxref_g 0.00917664f $X=0.07 $Y=3.02 $X2=0.24
+ $Y2=8.14
cc_208 LVPWR N_A_816_1221#_c_484_n 0.0393386f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_209 LVPWR N_A_1406_429#_c_572_n 0.0108188f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_210 LVPWR N_A_1406_429#_M17_noxref_g 0.0151226f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_211 LVPWR N_VPWR_M17_noxref_d 0.00297482f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_212 LVPWR N_VPWR_c_672_n 0.0428658f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_213 N_LVPWR_M1005_b N_VPWR_c_668_n 0.00618401f $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_214 N_LVPWR_c_175_n N_VPWR_c_668_n 0.0268368f $X=3.93 $Y=3.19 $X2=0 $Y2=0
cc_215 LVPWR N_VPWR_c_683_n 0.0674099f $X=0.07 $Y=3.02 $X2=5.52 $Y2=0.06
cc_216 N_LVPWR_M1005_b N_VPWR_c_669_n 0.00793792f $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_217 LVPWR N_VPWR_c_669_n 1.13227f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_218 N_LVPWR_c_175_n N_VPWR_c_669_n 0.0680381f $X=3.93 $Y=3.19 $X2=0 $Y2=0
cc_219 N_A_c_227_n N_A_573_897#_c_261_n 0.014409f $X=3.355 $Y=1.705 $X2=0
+ $Y2=8.025
cc_220 N_A_M1005_g N_A_573_897#_M1017_g 0.019196f $X=3.355 $Y=2.615 $X2=0.24
+ $Y2=0
cc_221 N_A_c_228_n N_A_573_897#_c_263_n 0.0226068f $X=3.355 $Y=1.87 $X2=0 $Y2=0
cc_222 N_A_M1005_g N_A_573_897#_c_264_n 0.00201071f $X=3.355 $Y=2.615 $X2=0
+ $Y2=0
cc_223 N_A_c_226_n N_A_573_897#_c_266_n 0.00930167f $X=3.28 $Y=1.87 $X2=0 $Y2=0
cc_224 N_A_c_227_n N_A_573_897#_c_266_n 0.00615095f $X=3.355 $Y=1.705 $X2=0
+ $Y2=0
cc_225 A N_A_573_897#_c_266_n 0.0165667f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_226 N_A_c_230_n N_A_573_897#_c_266_n 0.00155799f $X=2.66 $Y=1.695 $X2=0 $Y2=0
cc_227 N_A_c_226_n N_A_573_897#_c_281_n 0.00930167f $X=3.28 $Y=1.87 $X2=5.52
+ $Y2=0.06
cc_228 N_A_M1005_g N_A_573_897#_c_281_n 0.00805052f $X=3.355 $Y=2.615 $X2=5.52
+ $Y2=0.06
cc_229 A N_A_573_897#_c_281_n 0.015787f $X=2.555 $Y=1.58 $X2=5.52 $Y2=0.06
cc_230 N_A_c_230_n N_A_573_897#_c_281_n 0.00146896f $X=2.66 $Y=1.695 $X2=5.52
+ $Y2=0.06
cc_231 N_A_c_226_n N_A_573_897#_c_267_n 0.00131023f $X=3.28 $Y=1.87 $X2=5.52
+ $Y2=8.08
cc_232 N_A_c_228_n N_A_573_897#_c_267_n 0.0196537f $X=3.355 $Y=1.87 $X2=5.52
+ $Y2=8.08
cc_233 N_A_c_226_n N_A_573_897#_c_301_n 0.0104509f $X=3.28 $Y=1.87 $X2=0 $Y2=0
cc_234 A N_A_573_897#_c_301_n 0.0198664f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_235 N_A_M1005_g N_VPWR_c_669_n 3.17298e-19 $X=3.355 $Y=2.615 $X2=0 $Y2=0
cc_236 N_A_c_227_n N_VGND_c_771_n 0.00386936f $X=3.355 $Y=1.705 $X2=0 $Y2=0
cc_237 N_A_c_227_n N_VGND_c_780_n 0.00555051f $X=3.355 $Y=1.705 $X2=10.8
+ $Y2=8.14
cc_238 N_A_c_227_n N_VGND_c_788_n 0.00523016f $X=3.355 $Y=1.705 $X2=0 $Y2=0
cc_239 N_A_573_897#_c_261_n N_A_772_151#_c_342_n 0.00286882f $X=3.785 $Y=1.705
+ $X2=0 $Y2=0
cc_240 N_A_573_897#_c_261_n N_A_772_151#_c_343_n 0.00280304f $X=3.785 $Y=1.705
+ $X2=0 $Y2=0
cc_241 N_A_573_897#_M1017_g N_A_772_151#_c_343_n 0.00253691f $X=3.785 $Y=2.615
+ $X2=0 $Y2=0
cc_242 N_A_573_897#_c_267_n N_A_772_151#_c_343_n 0.020811f $X=4.145 $Y=1.87
+ $X2=0 $Y2=0
cc_243 N_A_573_897#_c_268_n N_A_772_151#_c_343_n 0.00542196f $X=4.145 $Y=1.87
+ $X2=0 $Y2=0
cc_244 N_A_573_897#_M1017_g N_A_772_151#_c_344_n 0.00123902f $X=3.785 $Y=2.615
+ $X2=0 $Y2=0
cc_245 N_A_573_897#_c_267_n N_A_772_151#_c_344_n 0.0353505f $X=4.145 $Y=1.87
+ $X2=0 $Y2=0
cc_246 N_A_573_897#_c_268_n N_A_772_151#_c_344_n 0.0105631f $X=4.145 $Y=1.87
+ $X2=0 $Y2=0
cc_247 N_A_573_897#_c_267_n N_A_772_151#_c_345_n 0.0316368f $X=4.145 $Y=1.87
+ $X2=0 $Y2=0
cc_248 N_A_573_897#_c_268_n N_A_772_151#_c_345_n 0.0102771f $X=4.145 $Y=1.87
+ $X2=0 $Y2=0
cc_249 N_A_573_897#_c_260_n N_A_816_1221#_c_497_n 0.0401197f $X=3.83 $Y=5.995
+ $X2=0 $Y2=0
cc_250 N_A_573_897#_c_262_n N_A_816_1221#_c_497_n 0.0401197f $X=4.61 $Y=5.995
+ $X2=0 $Y2=0
cc_251 N_A_573_897#_c_262_n N_A_816_1221#_c_464_n 0.059011f $X=4.61 $Y=5.995
+ $X2=0 $Y2=0
cc_252 N_A_573_897#_c_262_n N_A_816_1221#_c_465_n 0.0346695f $X=4.61 $Y=5.995
+ $X2=5.52 $Y2=0.057
cc_253 N_A_573_897#_c_264_n N_VPWR_c_668_n 0.0547753f $X=3.03 $Y=4.65 $X2=0
+ $Y2=0
cc_254 N_A_573_897#_c_265_n N_VPWR_c_668_n 0.00922839f $X=3.03 $Y=4.65 $X2=0
+ $Y2=0
cc_255 N_A_573_897#_c_264_n N_VPWR_c_669_n 0.0361756f $X=3.03 $Y=4.65 $X2=0
+ $Y2=0
cc_256 N_A_573_897#_c_285_n N_VPWR_c_669_n 3.87848e-19 $X=3.075 $Y=3.055 $X2=0
+ $Y2=0
cc_257 N_A_573_897#_c_261_n N_VGND_c_771_n 0.00386936f $X=3.785 $Y=1.705 $X2=0
+ $Y2=0
cc_258 N_A_573_897#_c_263_n N_VGND_c_771_n 0.00139629f $X=3.75 $Y=1.87 $X2=0
+ $Y2=0
cc_259 N_A_573_897#_c_266_n N_VGND_c_771_n 0.001542f $X=3.14 $Y=0.9 $X2=0 $Y2=0
cc_260 N_A_573_897#_c_267_n N_VGND_c_771_n 0.0179406f $X=4.145 $Y=1.87 $X2=0
+ $Y2=0
cc_261 N_A_573_897#_c_260_n N_VGND_c_772_n 0.0146836f $X=3.83 $Y=5.995 $X2=10.8
+ $Y2=0
cc_262 N_A_573_897#_c_262_n N_VGND_c_772_n 0.0181045f $X=4.61 $Y=5.995 $X2=10.8
+ $Y2=0
cc_263 N_A_573_897#_c_260_n N_VGND_c_774_n 0.0034209f $X=3.83 $Y=5.995 $X2=0
+ $Y2=0
cc_264 N_A_573_897#_c_266_n N_VGND_c_780_n 0.0123012f $X=3.14 $Y=0.9 $X2=10.8
+ $Y2=8.14
cc_265 N_A_573_897#_c_259_n N_VGND_c_782_n 0.0176616f $X=3.195 $Y=5.83 $X2=5.52
+ $Y2=0.057
cc_266 N_A_573_897#_c_260_n N_VGND_c_782_n 0.0635146f $X=3.83 $Y=5.995 $X2=5.52
+ $Y2=0.057
cc_267 N_A_573_897#_c_262_n N_VGND_c_782_n 0.00129485f $X=4.61 $Y=5.995 $X2=5.52
+ $Y2=0.057
cc_268 N_A_573_897#_c_264_n N_VGND_c_782_n 8.6599e-19 $X=3.03 $Y=4.65 $X2=5.52
+ $Y2=0.057
cc_269 N_A_573_897#_c_261_n N_VGND_c_783_n 0.00555051f $X=3.785 $Y=1.705 $X2=0
+ $Y2=0
cc_270 N_A_573_897#_c_260_n N_VGND_c_785_n 0.00129485f $X=3.83 $Y=5.995 $X2=0
+ $Y2=0
cc_271 N_A_573_897#_c_262_n N_VGND_c_785_n 0.0582646f $X=4.61 $Y=5.995 $X2=0
+ $Y2=0
cc_272 N_A_573_897#_c_261_n N_VGND_c_788_n 0.00523016f $X=3.785 $Y=1.705 $X2=0
+ $Y2=0
cc_273 N_A_573_897#_c_266_n N_VGND_c_788_n 0.0105954f $X=3.14 $Y=0.9 $X2=0 $Y2=0
cc_274 N_A_573_897#_c_260_n N_VGND_c_792_n 0.0157032f $X=3.83 $Y=5.995 $X2=0
+ $Y2=0
cc_275 N_A_573_897#_c_262_n N_VGND_c_792_n 0.0157032f $X=4.61 $Y=5.995 $X2=0
+ $Y2=0
cc_276 N_A_772_151#_c_341_n N_A_816_1221#_c_484_n 0.00523594f $X=6.515 $Y=2.145
+ $X2=0 $Y2=0
cc_277 N_A_772_151#_c_341_n N_A_1406_429#_c_572_n 0.019016f $X=6.515 $Y=2.145
+ $X2=0 $Y2=0
cc_278 N_A_772_151#_c_342_n N_VGND_c_771_n 0.00154986f $X=4 $Y=0.9 $X2=0 $Y2=0
cc_279 N_A_772_151#_c_340_n N_VGND_c_776_n 0.0146836f $X=5.735 $Y=2.145 $X2=0
+ $Y2=0
cc_280 N_A_772_151#_c_341_n N_VGND_c_776_n 0.0181045f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_281 N_A_772_151#_c_340_n N_VGND_c_778_n 0.0034209f $X=5.735 $Y=2.145 $X2=0
+ $Y2=0
cc_282 N_A_772_151#_c_342_n N_VGND_c_783_n 0.0120367f $X=4 $Y=0.9 $X2=0 $Y2=0
cc_283 N_A_772_151#_c_340_n N_VGND_c_786_n 0.0582646f $X=5.735 $Y=2.145 $X2=0
+ $Y2=0
cc_284 N_A_772_151#_c_341_n N_VGND_c_786_n 0.00129485f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_285 N_A_772_151#_c_343_n N_VGND_c_786_n 0.027388f $X=4.645 $Y=2.145 $X2=0
+ $Y2=0
cc_286 N_A_772_151#_c_352_n N_VGND_c_786_n 0.0457912f $X=5.625 $Y=2.31 $X2=0
+ $Y2=0
cc_287 N_A_772_151#_c_345_n N_VGND_c_786_n 0.0237705f $X=4.645 $Y=1.41 $X2=0
+ $Y2=0
cc_288 N_A_772_151#_c_346_n N_VGND_c_786_n 0.00991638f $X=5.485 $Y=2.31 $X2=0
+ $Y2=0
cc_289 N_A_772_151#_c_340_n N_VGND_c_787_n 0.00129485f $X=5.735 $Y=2.145 $X2=0
+ $Y2=0
cc_290 N_A_772_151#_c_341_n N_VGND_c_787_n 0.0582646f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_291 N_A_772_151#_c_340_n N_VGND_c_788_n 0.0157032f $X=5.735 $Y=2.145 $X2=0
+ $Y2=0
cc_292 N_A_772_151#_c_341_n N_VGND_c_788_n 0.0157032f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_293 N_A_772_151#_c_342_n N_VGND_c_788_n 0.0112977f $X=4 $Y=0.9 $X2=0 $Y2=0
cc_294 N_A_772_151#_c_340_n N_A_1197_107#_c_874_n 0.0401197f $X=5.735 $Y=2.145
+ $X2=0 $Y2=8.025
cc_295 N_A_772_151#_c_341_n N_A_1197_107#_c_874_n 0.0401197f $X=6.515 $Y=2.145
+ $X2=0 $Y2=8.025
cc_296 N_A_772_151#_c_341_n N_A_1197_107#_c_867_n 0.0402565f $X=6.515 $Y=2.145
+ $X2=0.24 $Y2=0
cc_297 N_A_772_151#_c_341_n N_A_1197_107#_c_877_n 0.0255423f $X=6.515 $Y=2.145
+ $X2=0.24 $Y2=0
cc_298 N_A_772_151#_c_352_n N_A_1197_107#_c_877_n 0.0151525f $X=5.625 $Y=2.31
+ $X2=0.24 $Y2=0
cc_299 N_A_1400_777#_c_397_n N_A_816_1221#_M15_noxref_g 0.00249821f $X=7.6
+ $Y=4.05 $X2=0.24 $Y2=8.14
cc_300 N_A_1400_777#_c_401_n N_A_816_1221#_M15_noxref_g 0.100961f $X=8.465
+ $Y=2.495 $X2=0.24 $Y2=8.14
cc_301 N_A_1400_777#_c_394_n N_A_816_1221#_c_484_n 0.092172f $X=7.6 $Y=4.05
+ $X2=0 $Y2=0
cc_302 N_A_1400_777#_c_397_n N_A_816_1221#_c_484_n 0.0157312f $X=7.6 $Y=4.05
+ $X2=0 $Y2=0
cc_303 N_A_1400_777#_M1008_g N_A_816_1221#_c_486_n 0.0226969f $X=7.25 $Y=5.175
+ $X2=0 $Y2=0
cc_304 N_A_1400_777#_M1008_g N_A_816_1221#_c_466_n 0.00407172f $X=7.25 $Y=5.175
+ $X2=5.52 $Y2=8.14
cc_305 N_A_1400_777#_c_390_n N_A_816_1221#_c_466_n 0.0160763f $X=8.075 $Y=6.055
+ $X2=5.52 $Y2=8.14
cc_306 N_A_1400_777#_c_390_n N_A_816_1221#_c_467_n 0.0799786f $X=8.075 $Y=6.055
+ $X2=0 $Y2=0
cc_307 N_A_1400_777#_c_390_n N_A_816_1221#_c_468_n 0.00272945f $X=8.075 $Y=6.055
+ $X2=0 $Y2=0
cc_308 N_A_1400_777#_c_390_n N_A_816_1221#_c_469_n 0.0160763f $X=8.075 $Y=6.055
+ $X2=0 $Y2=0
cc_309 N_A_1400_777#_M1009_g N_A_816_1221#_c_469_n 0.0414133f $X=8.075 $Y=5.175
+ $X2=0 $Y2=0
cc_310 N_A_1400_777#_M1008_g N_A_816_1221#_c_491_n 0.0067799f $X=7.25 $Y=5.175
+ $X2=0 $Y2=0
cc_311 N_A_1400_777#_M1008_g N_A_816_1221#_c_493_n 0.0111918f $X=7.25 $Y=5.175
+ $X2=0 $Y2=0
cc_312 N_A_1400_777#_c_390_n N_A_816_1221#_c_470_n 0.00162697f $X=8.075 $Y=6.055
+ $X2=0 $Y2=0
cc_313 N_A_1400_777#_c_390_n N_A_816_1221#_c_471_n 0.00654091f $X=8.075 $Y=6.055
+ $X2=0 $Y2=0
cc_314 N_A_1400_777#_c_404_n N_A_1406_429#_c_569_n 0.0566308f $X=8.465 $Y=0.68
+ $X2=0 $Y2=0
cc_315 N_A_1400_777#_c_404_n N_A_1406_429#_c_570_n 0.0589667f $X=8.465 $Y=0.68
+ $X2=0 $Y2=0
cc_316 N_A_1400_777#_c_394_n N_A_1406_429#_c_572_n 0.0741581f $X=7.6 $Y=4.05
+ $X2=0 $Y2=0
cc_317 N_A_1400_777#_c_397_n N_A_1406_429#_c_572_n 0.0202601f $X=7.6 $Y=4.05
+ $X2=0 $Y2=0
cc_318 N_A_1400_777#_c_400_n N_A_1406_429#_c_572_n 0.0264615f $X=8.17 $Y=2.6
+ $X2=0 $Y2=0
cc_319 N_A_1400_777#_c_429_p N_A_1406_429#_c_572_n 0.0321807f $X=7.765 $Y=2.6
+ $X2=0 $Y2=0
cc_320 N_A_1400_777#_c_401_n N_A_1406_429#_c_572_n 0.0345162f $X=8.465 $Y=2.495
+ $X2=0 $Y2=0
cc_321 N_A_1400_777#_c_404_n N_A_1406_429#_c_572_n 0.0581717f $X=8.465 $Y=0.68
+ $X2=0 $Y2=0
cc_322 N_A_1400_777#_c_401_n N_A_1406_429#_M17_noxref_g 0.0217522f $X=8.465
+ $Y=2.495 $X2=0 $Y2=0
cc_323 N_A_1400_777#_M1009_g N_A_1406_429#_c_587_n 0.00417504f $X=8.075 $Y=5.175
+ $X2=0 $Y2=0
cc_324 N_A_1400_777#_c_390_n N_A_1406_429#_c_579_n 3.0034e-19 $X=8.075 $Y=6.055
+ $X2=5.52 $Y2=8.08
cc_325 N_A_1400_777#_M1008_g N_VPWR_c_670_n 0.0513745f $X=7.25 $Y=5.175 $X2=0
+ $Y2=0
cc_326 N_A_1400_777#_c_390_n N_VPWR_c_670_n 0.00406276f $X=8.075 $Y=6.055 $X2=0
+ $Y2=0
cc_327 N_A_1400_777#_M1009_g N_VPWR_c_670_n 0.0591544f $X=8.075 $Y=5.175 $X2=0
+ $Y2=0
cc_328 N_A_1400_777#_c_394_n N_VPWR_c_670_n 0.0229228f $X=7.6 $Y=4.05 $X2=0
+ $Y2=0
cc_329 N_A_1400_777#_c_397_n N_VPWR_c_670_n 0.00320086f $X=7.6 $Y=4.05 $X2=0
+ $Y2=0
cc_330 N_A_1400_777#_c_394_n N_VPWR_c_672_n 0.0559598f $X=7.6 $Y=4.05 $X2=0
+ $Y2=0
cc_331 N_A_1400_777#_c_397_n N_VPWR_c_672_n 0.00878144f $X=7.6 $Y=4.05 $X2=0
+ $Y2=0
cc_332 N_A_1400_777#_c_400_n N_VPWR_c_672_n 0.0138302f $X=8.17 $Y=2.6 $X2=0
+ $Y2=0
cc_333 N_A_1400_777#_c_401_n N_VPWR_c_672_n 0.0495989f $X=8.465 $Y=2.495 $X2=0
+ $Y2=0
cc_334 N_A_1400_777#_M1008_g N_VPWR_c_668_n 0.0199766f $X=7.25 $Y=5.175 $X2=0
+ $Y2=0
cc_335 N_A_1400_777#_M1009_g N_VPWR_c_668_n 0.0172597f $X=8.075 $Y=5.175 $X2=0
+ $Y2=0
cc_336 N_A_1400_777#_c_394_n N_VPWR_c_668_n 0.011691f $X=7.6 $Y=4.05 $X2=0 $Y2=0
cc_337 N_A_1400_777#_c_397_n N_VPWR_c_668_n 0.0110402f $X=7.6 $Y=4.05 $X2=0
+ $Y2=0
cc_338 N_A_1400_777#_c_401_n N_VPWR_c_683_n 0.0325388f $X=8.465 $Y=2.495
+ $X2=5.52 $Y2=0.06
cc_339 N_A_1400_777#_c_394_n N_VPWR_c_669_n 0.0567963f $X=7.6 $Y=4.05 $X2=0
+ $Y2=0
cc_340 N_A_1400_777#_c_397_n N_VPWR_c_669_n 0.00562867f $X=7.6 $Y=4.05 $X2=0
+ $Y2=0
cc_341 N_A_1400_777#_c_401_n N_VPWR_c_669_n 0.032272f $X=8.465 $Y=2.495 $X2=0
+ $Y2=0
cc_342 N_A_1400_777#_c_404_n N_VGND_c_788_n 0.0423355f $X=8.465 $Y=0.68 $X2=0
+ $Y2=0
cc_343 N_A_1400_777#_c_400_n N_A_1197_107#_c_867_n 0.00653533f $X=8.17 $Y=2.6
+ $X2=0.24 $Y2=0
cc_344 N_A_1400_777#_c_429_p N_A_1197_107#_c_867_n 0.0532075f $X=7.765 $Y=2.6
+ $X2=0.24 $Y2=0
cc_345 N_A_1400_777#_c_404_n N_A_1197_107#_c_867_n 0.00902002f $X=8.465 $Y=0.68
+ $X2=0.24 $Y2=0
cc_346 N_A_1400_777#_c_404_n N_A_1197_107#_c_868_n 0.0728339f $X=8.465 $Y=0.68
+ $X2=0 $Y2=0
cc_347 N_A_1400_777#_c_404_n N_A_1197_107#_c_869_n 0.0382279f $X=8.465 $Y=0.68
+ $X2=0 $Y2=0
cc_348 N_A_1400_777#_c_401_n N_A_1197_107#_c_873_n 0.0156266f $X=8.465 $Y=2.495
+ $X2=0.24 $Y2=8.14
cc_349 N_A_1400_777#_c_404_n N_A_1197_107#_c_873_n 0.0686214f $X=8.465 $Y=0.68
+ $X2=0.24 $Y2=8.14
cc_350 N_A_816_1221#_M15_noxref_g N_A_1406_429#_c_572_n 0.0837846f $X=8.97
+ $Y=3.025 $X2=0 $Y2=0
cc_351 N_A_816_1221#_c_484_n N_A_1406_429#_c_572_n 0.013688f $X=6.81 $Y=2.96
+ $X2=0 $Y2=0
cc_352 N_A_816_1221#_c_472_n N_A_1406_429#_c_582_n 0.00501669f $X=9.55 $Y=4.535
+ $X2=0.24 $Y2=0
cc_353 N_A_816_1221#_c_479_n N_A_1406_429#_c_582_n 0.0194762f $X=9.55 $Y=4.285
+ $X2=0.24 $Y2=0
cc_354 N_A_816_1221#_M15_noxref_g N_A_1406_429#_M17_noxref_g 0.0334585f $X=8.97
+ $Y=3.025 $X2=0 $Y2=0
cc_355 N_A_816_1221#_c_472_n N_A_1406_429#_M1014_g 0.0112759f $X=9.55 $Y=4.535
+ $X2=10.8 $Y2=0
cc_356 N_A_816_1221#_c_461_n N_A_1406_429#_M1014_g 0.00733127f $X=9.51 $Y=6.285
+ $X2=10.8 $Y2=0
cc_357 N_A_816_1221#_c_462_n N_A_1406_429#_M1007_g 0.0215296f $X=9.55 $Y=6.975
+ $X2=0 $Y2=0
cc_358 N_A_816_1221#_c_472_n N_A_1406_429#_c_587_n 0.00282356f $X=9.55 $Y=4.535
+ $X2=0 $Y2=0
cc_359 N_A_816_1221#_M1013_g N_A_1406_429#_c_587_n 0.0296294f $X=9.55 $Y=5.175
+ $X2=0 $Y2=0
cc_360 N_A_816_1221#_c_461_n N_A_1406_429#_c_587_n 0.0105971f $X=9.51 $Y=6.285
+ $X2=0 $Y2=0
cc_361 N_A_816_1221#_c_482_n N_A_1406_429#_c_587_n 0.0110834f $X=9.55 $Y=6.055
+ $X2=0 $Y2=0
cc_362 N_A_816_1221#_c_469_n N_A_1406_429#_c_587_n 0.0848056f $X=8.465 $Y=4.57
+ $X2=0 $Y2=0
cc_363 N_A_816_1221#_c_460_n N_A_1406_429#_c_575_n 0.00780381f $X=9.3 $Y=6.45
+ $X2=5.52 $Y2=0
cc_364 N_A_816_1221#_c_462_n N_A_1406_429#_c_575_n 0.0361306f $X=9.55 $Y=6.975
+ $X2=5.52 $Y2=0
cc_365 N_A_816_1221#_c_470_n N_A_1406_429#_c_575_n 0.0299745f $X=8.7 $Y=6.45
+ $X2=5.52 $Y2=0
cc_366 N_A_816_1221#_c_471_n N_A_1406_429#_c_575_n 0.00313758f $X=8.7 $Y=6.45
+ $X2=5.52 $Y2=0
cc_367 N_A_816_1221#_c_461_n N_A_1406_429#_c_577_n 0.0206482f $X=9.51 $Y=6.285
+ $X2=5.52 $Y2=0.06
cc_368 N_A_816_1221#_c_462_n N_A_1406_429#_c_577_n 0.0315255f $X=9.55 $Y=6.975
+ $X2=5.52 $Y2=0.06
cc_369 N_A_816_1221#_c_482_n N_A_1406_429#_c_577_n 0.00111228f $X=9.55 $Y=6.055
+ $X2=5.52 $Y2=0.06
cc_370 N_A_816_1221#_c_461_n N_A_1406_429#_c_578_n 0.0215844f $X=9.51 $Y=6.285
+ $X2=0 $Y2=0
cc_371 N_A_816_1221#_c_460_n N_A_1406_429#_c_579_n 0.0192396f $X=9.3 $Y=6.45
+ $X2=5.52 $Y2=8.08
cc_372 N_A_816_1221#_c_462_n N_A_1406_429#_c_579_n 6.3561e-19 $X=9.55 $Y=6.975
+ $X2=5.52 $Y2=8.08
cc_373 N_A_816_1221#_c_469_n N_A_1406_429#_c_579_n 0.00309819f $X=8.465 $Y=4.57
+ $X2=5.52 $Y2=8.08
cc_374 N_A_816_1221#_c_470_n N_A_1406_429#_c_579_n 0.0218197f $X=8.7 $Y=6.45
+ $X2=5.52 $Y2=8.08
cc_375 N_A_816_1221#_c_467_n N_VPWR_c_670_n 0.0283836f $X=8.3 $Y=6.45 $X2=0
+ $Y2=0
cc_376 N_A_816_1221#_c_469_n N_VPWR_c_670_n 0.0682339f $X=8.465 $Y=4.57 $X2=0
+ $Y2=0
cc_377 N_A_816_1221#_c_491_n N_VPWR_c_670_n 0.0488156f $X=6.86 $Y=4.57 $X2=0
+ $Y2=0
cc_378 N_A_816_1221#_c_493_n N_VPWR_c_670_n 0.0126f $X=6.86 $Y=5.78 $X2=0 $Y2=0
cc_379 N_A_816_1221#_M15_noxref_g N_VPWR_c_672_n 0.0398607f $X=8.97 $Y=3.025
+ $X2=0 $Y2=0
cc_380 N_A_816_1221#_c_472_n N_VPWR_c_675_n 0.00410736f $X=9.55 $Y=4.535
+ $X2=10.8 $Y2=8.14
cc_381 N_A_816_1221#_M1013_g N_VPWR_c_675_n 0.040127f $X=9.55 $Y=5.175 $X2=10.8
+ $Y2=8.14
cc_382 N_A_816_1221#_c_482_n N_VPWR_c_675_n 0.00618186f $X=9.55 $Y=6.055
+ $X2=10.8 $Y2=8.14
cc_383 N_A_816_1221#_c_472_n N_VPWR_c_668_n 0.00547212f $X=9.55 $Y=4.535 $X2=0
+ $Y2=0
cc_384 N_A_816_1221#_M1013_g N_VPWR_c_668_n 0.017691f $X=9.55 $Y=5.175 $X2=0
+ $Y2=0
cc_385 N_A_816_1221#_c_484_n N_VPWR_c_668_n 0.0127452f $X=6.81 $Y=2.96 $X2=0
+ $Y2=0
cc_386 N_A_816_1221#_c_469_n N_VPWR_c_668_n 0.0415768f $X=8.465 $Y=4.57 $X2=0
+ $Y2=0
cc_387 N_A_816_1221#_c_491_n N_VPWR_c_668_n 0.0577545f $X=6.86 $Y=4.57 $X2=0
+ $Y2=0
cc_388 N_A_816_1221#_M15_noxref_g N_VPWR_c_683_n 0.00205779f $X=8.97 $Y=3.025
+ $X2=5.52 $Y2=0.06
cc_389 N_A_816_1221#_M13_noxref_s N_VPWR_c_669_n 4.93918e-19 $X=6.665 $Y=2.815
+ $X2=0 $Y2=0
cc_390 N_A_816_1221#_M15_noxref_g N_VPWR_c_669_n 0.0241983f $X=8.97 $Y=3.025
+ $X2=0 $Y2=0
cc_391 N_A_816_1221#_c_484_n N_VPWR_c_669_n 0.0395191f $X=6.81 $Y=2.96 $X2=0
+ $Y2=0
cc_392 N_A_816_1221#_c_497_n N_VGND_c_772_n 0.0211458f $X=4.22 $Y=6.25 $X2=10.8
+ $Y2=0
cc_393 N_A_816_1221#_c_497_n N_VGND_c_782_n 0.0648349f $X=4.22 $Y=6.25 $X2=5.52
+ $Y2=0.057
cc_394 N_A_816_1221#_c_497_n N_VGND_c_785_n 0.0648349f $X=4.22 $Y=6.25 $X2=0
+ $Y2=0
cc_395 N_A_816_1221#_c_464_n N_VGND_c_785_n 0.0476157f $X=6.695 $Y=5.83 $X2=0
+ $Y2=0
cc_396 N_A_816_1221#_c_462_n N_VGND_c_790_n 0.0340179f $X=9.55 $Y=6.975 $X2=0
+ $Y2=0
cc_397 N_A_816_1221#_c_462_n N_VGND_c_792_n 0.0241606f $X=9.55 $Y=6.975 $X2=0
+ $Y2=0
cc_398 N_A_816_1221#_c_497_n N_VGND_c_792_n 0.0240827f $X=4.22 $Y=6.25 $X2=0
+ $Y2=0
cc_399 N_A_816_1221#_c_470_n N_VGND_c_792_n 0.00990816f $X=8.7 $Y=6.45 $X2=0
+ $Y2=0
cc_400 N_A_816_1221#_c_471_n N_VGND_c_792_n 0.00128885f $X=8.7 $Y=6.45 $X2=0
+ $Y2=0
cc_401 N_A_816_1221#_c_484_n N_A_1197_107#_c_867_n 0.0129567f $X=6.81 $Y=2.96
+ $X2=0.24 $Y2=0
cc_402 N_A_1406_429#_c_572_n N_VPWR_c_672_n 0.0207994f $X=9.105 $Y=2.31 $X2=0
+ $Y2=0
cc_403 N_A_1406_429#_c_582_n N_VPWR_c_675_n 0.00326676f $X=10.16 $Y=3.905
+ $X2=10.8 $Y2=8.14
cc_404 N_A_1406_429#_M1014_g N_VPWR_c_675_n 0.0571855f $X=10.375 $Y=5.175
+ $X2=10.8 $Y2=8.14
cc_405 N_A_1406_429#_c_587_n N_VPWR_c_675_n 0.0606729f $X=9.16 $Y=4.57 $X2=10.8
+ $Y2=8.14
cc_406 N_A_1406_429#_c_577_n N_VPWR_c_675_n 0.0338611f $X=10.435 $Y=6.39
+ $X2=10.8 $Y2=8.14
cc_407 N_A_1406_429#_c_578_n N_VPWR_c_675_n 0.00426906f $X=10.435 $Y=6.39
+ $X2=10.8 $Y2=8.14
cc_408 N_A_1406_429#_c_582_n N_VPWR_c_668_n 0.00510566f $X=10.16 $Y=3.905 $X2=0
+ $Y2=0
cc_409 N_A_1406_429#_M1014_g N_VPWR_c_668_n 0.0174718f $X=10.375 $Y=5.175 $X2=0
+ $Y2=0
cc_410 N_A_1406_429#_c_587_n N_VPWR_c_668_n 0.0419805f $X=9.16 $Y=4.57 $X2=0
+ $Y2=0
cc_411 N_A_1406_429#_c_582_n N_VPWR_c_683_n 0.00251001f $X=10.16 $Y=3.905
+ $X2=5.52 $Y2=0.06
cc_412 N_A_1406_429#_M17_noxref_g N_VPWR_c_683_n 0.0728548f $X=10.16 $Y=3.025
+ $X2=5.52 $Y2=0.06
cc_413 N_A_1406_429#_c_572_n N_VPWR_c_669_n 0.00214842f $X=9.105 $Y=2.31 $X2=0
+ $Y2=0
cc_414 N_A_1406_429#_c_582_n N_VPWR_c_669_n 0.00188968f $X=10.16 $Y=3.905 $X2=0
+ $Y2=0
cc_415 N_A_1406_429#_M17_noxref_g N_VPWR_c_669_n 0.0110143f $X=10.16 $Y=3.025
+ $X2=0 $Y2=0
cc_416 N_A_1406_429#_M1014_g X 0.00967557f $X=10.375 $Y=5.175 $X2=-0.33
+ $Y2=-0.265
cc_417 N_A_1406_429#_M1007_g X 0.0271496f $X=10.375 $Y=7.23 $X2=0 $Y2=0
cc_418 N_A_1406_429#_M1014_g N_X_c_758_n 0.0322003f $X=10.375 $Y=5.175 $X2=0
+ $Y2=0
cc_419 N_A_1406_429#_M1014_g X 0.0254153f $X=10.375 $Y=5.175 $X2=0 $Y2=0
cc_420 N_A_1406_429#_c_577_n X 0.0268756f $X=10.435 $Y=6.39 $X2=0 $Y2=0
cc_421 N_A_1406_429#_c_569_n N_VGND_c_787_n 0.00364283f $X=8.075 $Y=2.145 $X2=0
+ $Y2=0
cc_422 N_A_1406_429#_c_572_n N_VGND_c_787_n 0.00460353f $X=9.105 $Y=2.31 $X2=0
+ $Y2=0
cc_423 N_A_1406_429#_c_569_n N_VGND_c_788_n 0.0157093f $X=8.075 $Y=2.145 $X2=0
+ $Y2=0
cc_424 N_A_1406_429#_c_570_n N_VGND_c_788_n 0.0157093f $X=8.855 $Y=2.145 $X2=0
+ $Y2=0
cc_425 N_A_1406_429#_M1007_g N_VGND_c_790_n 0.0387435f $X=10.375 $Y=7.23 $X2=0
+ $Y2=0
cc_426 N_A_1406_429#_c_575_n N_VGND_c_790_n 0.0317368f $X=9.16 $Y=7 $X2=0 $Y2=0
cc_427 N_A_1406_429#_c_577_n N_VGND_c_790_n 0.0338611f $X=10.435 $Y=6.39 $X2=0
+ $Y2=0
cc_428 N_A_1406_429#_c_578_n N_VGND_c_790_n 0.00426906f $X=10.435 $Y=6.39 $X2=0
+ $Y2=0
cc_429 N_A_1406_429#_M1007_g N_VGND_c_792_n 0.0208706f $X=10.375 $Y=7.23 $X2=0
+ $Y2=0
cc_430 N_A_1406_429#_c_575_n N_VGND_c_792_n 0.0338942f $X=9.16 $Y=7 $X2=0 $Y2=0
cc_431 N_A_1406_429#_c_572_n N_A_1197_107#_c_867_n 0.0531829f $X=9.105 $Y=2.31
+ $X2=0.24 $Y2=0
cc_432 N_A_1406_429#_c_569_n N_A_1197_107#_c_868_n 0.0433707f $X=8.075 $Y=2.145
+ $X2=0 $Y2=0
cc_433 N_A_1406_429#_c_569_n N_A_1197_107#_c_869_n 0.0181468f $X=8.075 $Y=2.145
+ $X2=0 $Y2=0
cc_434 N_A_1406_429#_c_570_n N_A_1197_107#_c_869_n 0.019032f $X=8.855 $Y=2.145
+ $X2=0 $Y2=0
cc_435 N_A_1406_429#_c_569_n N_A_1197_107#_c_871_n 8.85221e-19 $X=8.075 $Y=2.145
+ $X2=0 $Y2=0
cc_436 N_A_1406_429#_c_570_n N_A_1197_107#_c_873_n 0.0400673f $X=8.855 $Y=2.145
+ $X2=0.24 $Y2=8.14
cc_437 N_A_1406_429#_c_571_n N_A_1197_107#_c_873_n 0.00920651f $X=9.91 $Y=2.31
+ $X2=0.24 $Y2=8.14
cc_438 N_VPWR_c_675_n N_X_c_758_n 0.0682113f $X=9.985 $Y=4.57 $X2=0 $Y2=0
cc_439 N_VPWR_c_668_n N_X_c_758_n 0.0434272f $X=10.165 $Y=4.58 $X2=0 $Y2=0
cc_440 X N_VGND_c_790_n 0.0356028f $X=10.715 $Y=6.76 $X2=0 $Y2=0
cc_441 X N_VGND_c_792_n 0.0326456f $X=10.715 $Y=6.76 $X2=0 $Y2=0
cc_442 N_VGND_c_776_n N_A_1197_107#_c_874_n 0.0211458f $X=6.61 $Y=0.34 $X2=0
+ $Y2=8.025
cc_443 N_VGND_c_786_n N_A_1197_107#_c_874_n 0.0648349f $X=5.525 $Y=0.51 $X2=0
+ $Y2=8.025
cc_444 N_VGND_c_787_n N_A_1197_107#_c_874_n 0.0648349f $X=7.085 $Y=0.51 $X2=0
+ $Y2=8.025
cc_445 N_VGND_c_788_n N_A_1197_107#_c_874_n 0.0240827f $X=7.085 $Y=0.51 $X2=0
+ $Y2=8.025
cc_446 N_VGND_c_787_n N_A_1197_107#_c_867_n 0.0448636f $X=7.085 $Y=0.51 $X2=0.24
+ $Y2=0
cc_447 N_VGND_c_787_n N_A_1197_107#_c_868_n 0.0836091f $X=7.085 $Y=0.51 $X2=0
+ $Y2=0
cc_448 N_VGND_c_788_n N_A_1197_107#_c_868_n 0.0346286f $X=7.085 $Y=0.51 $X2=0
+ $Y2=0
cc_449 N_VGND_c_788_n N_A_1197_107#_c_869_n 0.0537714f $X=7.085 $Y=0.51 $X2=0
+ $Y2=0
cc_450 N_VGND_c_776_n N_A_1197_107#_c_871_n 0.00674464f $X=6.61 $Y=0.34 $X2=0
+ $Y2=0
cc_451 N_VGND_c_788_n N_A_1197_107#_c_871_n 0.00925923f $X=7.085 $Y=0.51 $X2=0
+ $Y2=0
cc_452 N_VGND_c_788_n N_A_1197_107#_c_873_n 0.0381848f $X=7.085 $Y=0.51 $X2=0.24
+ $Y2=8.14
