* File: sky130_fd_sc_hvl__buf_32.spice
* Created: Wed Sep  2 09:04:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__buf_32.pex.spice"
.subckt sky130_fd_sc_hvl__buf_32  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_M1008_g N_A_183_141#_M1008_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1012 N_VGND_M1012_d N_A_M1012_g N_A_183_141#_M1008_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250001
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1027 N_VGND_M1012_d N_A_M1027_g N_A_183_141#_M1027_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250002
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1028 N_VGND_M1028_d N_A_M1028_g N_A_183_141#_M1027_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250002
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1032 N_VGND_M1028_d N_A_M1032_g N_A_183_141#_M1032_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250003
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1043 N_VGND_M1043_d N_A_M1043_g N_A_183_141#_M1032_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250004
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1051 N_VGND_M1043_d N_A_M1051_g N_A_183_141#_M1051_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250005
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1069 N_VGND_M1069_d N_A_M1069_g N_A_183_141#_M1051_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250005
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1074 N_VGND_M1069_d N_A_M1074_g N_A_183_141#_M1074_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250006
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1081 N_VGND_M1081_d N_A_M1081_g N_A_183_141#_M1074_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.195 AS=0.105 PD=1.27 PS=1.03 NRD=18.2286 NRS=0 M=1 R=1.5 SA=250007
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1002 N_X_M1002_d N_A_183_141#_M1002_g N_VGND_M1081_d N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.195 PD=1.03 PS=1.27 NRD=0 NRS=18.2286 M=1 R=1.5 SA=250008
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1003 N_X_M1002_d N_A_183_141#_M1003_g N_VGND_M1003_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250009
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1005 N_X_M1005_d N_A_183_141#_M1005_g N_VGND_M1003_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250010
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1007 N_X_M1005_d N_A_183_141#_M1007_g N_VGND_M1007_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250010
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1009 N_X_M1009_d N_A_183_141#_M1009_g N_VGND_M1007_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250011
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1010 N_X_M1009_d N_A_183_141#_M1010_g N_VGND_M1010_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250012
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1014 N_X_M1014_d N_A_183_141#_M1014_g N_VGND_M1010_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250013
+ SB=250020 A=0.375 P=2.5 MULT=1
MM1015 N_X_M1014_d N_A_183_141#_M1015_g N_VGND_M1015_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250014
+ SB=250019 A=0.375 P=2.5 MULT=1
MM1025 N_X_M1025_d N_A_183_141#_M1025_g N_VGND_M1015_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250014
+ SB=250018 A=0.375 P=2.5 MULT=1
MM1031 N_X_M1025_d N_A_183_141#_M1031_g N_VGND_M1031_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250015
+ SB=250017 A=0.375 P=2.5 MULT=1
MM1038 N_X_M1038_d N_A_183_141#_M1038_g N_VGND_M1031_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250016
+ SB=250016 A=0.375 P=2.5 MULT=1
MM1040 N_X_M1038_d N_A_183_141#_M1040_g N_VGND_M1040_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250017
+ SB=250016 A=0.375 P=2.5 MULT=1
MM1044 N_X_M1044_d N_A_183_141#_M1044_g N_VGND_M1040_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250017
+ SB=250015 A=0.375 P=2.5 MULT=1
MM1047 N_X_M1044_d N_A_183_141#_M1047_g N_VGND_M1047_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250018
+ SB=250014 A=0.375 P=2.5 MULT=1
MM1048 N_X_M1048_d N_A_183_141#_M1048_g N_VGND_M1047_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250019
+ SB=250013 A=0.375 P=2.5 MULT=1
MM1052 N_X_M1048_d N_A_183_141#_M1052_g N_VGND_M1052_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250012 A=0.375 P=2.5 MULT=1
MM1053 N_X_M1053_d N_A_183_141#_M1053_g N_VGND_M1052_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250012 A=0.375 P=2.5 MULT=1
MM1056 N_X_M1053_d N_A_183_141#_M1056_g N_VGND_M1056_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250011 A=0.375 P=2.5 MULT=1
MM1057 N_X_M1057_d N_A_183_141#_M1057_g N_VGND_M1056_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250010 A=0.375 P=2.5 MULT=1
MM1058 N_X_M1057_d N_A_183_141#_M1058_g N_VGND_M1058_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250009 A=0.375 P=2.5 MULT=1
MM1061 N_X_M1061_d N_A_183_141#_M1061_g N_VGND_M1058_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250009 A=0.375 P=2.5 MULT=1
MM1062 N_X_M1061_d N_A_183_141#_M1062_g N_VGND_M1062_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250008 A=0.375 P=2.5 MULT=1
MM1067 N_X_M1067_d N_A_183_141#_M1067_g N_VGND_M1062_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250007 A=0.375 P=2.5 MULT=1
MM1068 N_X_M1067_d N_A_183_141#_M1068_g N_VGND_M1068_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250006 A=0.375 P=2.5 MULT=1
MM1071 N_X_M1071_d N_A_183_141#_M1071_g N_VGND_M1068_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250005 A=0.375 P=2.5 MULT=1
MM1072 N_X_M1071_d N_A_183_141#_M1072_g N_VGND_M1072_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250005 A=0.375 P=2.5 MULT=1
MM1076 N_X_M1076_d N_A_183_141#_M1076_g N_VGND_M1072_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250004 A=0.375 P=2.5 MULT=1
MM1077 N_X_M1076_d N_A_183_141#_M1077_g N_VGND_M1077_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250003 A=0.375 P=2.5 MULT=1
MM1078 N_X_M1078_d N_A_183_141#_M1078_g N_VGND_M1077_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1079 N_X_M1078_d N_A_183_141#_M1079_g N_VGND_M1079_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1082 N_X_M1082_d N_A_183_141#_M1082_g N_VGND_M1079_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1083 N_X_M1082_d N_A_183_141#_M1083_g N_VGND_M1083_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250020
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_183_141#_M1000_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250020 A=0.75 P=4 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_183_141#_M1000_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001 SB=250020
+ A=0.75 P=4 MULT=1
MM1006 N_VPWR_M1001_d N_A_M1006_g N_A_183_141#_M1006_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002 SB=250020
+ A=0.75 P=4 MULT=1
MM1016 N_VPWR_M1016_d N_A_M1016_g N_A_183_141#_M1006_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002 SB=250020
+ A=0.75 P=4 MULT=1
MM1019 N_VPWR_M1016_d N_A_M1019_g N_A_183_141#_M1019_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250003 SB=250020
+ A=0.75 P=4 MULT=1
MM1035 N_VPWR_M1035_d N_A_M1035_g N_A_183_141#_M1019_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250004 SB=250020
+ A=0.75 P=4 MULT=1
MM1039 N_VPWR_M1035_d N_A_M1039_g N_A_183_141#_M1039_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250005 SB=250020
+ A=0.75 P=4 MULT=1
MM1049 N_VPWR_M1049_d N_A_M1049_g N_A_183_141#_M1039_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250005 SB=250020
+ A=0.75 P=4 MULT=1
MM1064 N_VPWR_M1049_d N_A_M1064_g N_A_183_141#_M1064_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250006 SB=250020
+ A=0.75 P=4 MULT=1
MM1070 N_VPWR_M1070_d N_A_M1070_g N_A_183_141#_M1064_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.39 AS=0.21 PD=2.02 PS=1.78 NRD=15.2609 NRS=0 M=1 R=3 SA=250007
+ SB=250020 A=0.75 P=4 MULT=1
MM1004 N_VPWR_M1070_d N_A_183_141#_M1004_g N_X_M1004_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.39 AS=0.21 PD=2.02 PS=1.78 NRD=15.2609 NRS=0 M=1 R=3 SA=250008
+ SB=250020 A=0.75 P=4 MULT=1
MM1011 N_VPWR_M1011_d N_A_183_141#_M1011_g N_X_M1004_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250009 SB=250020
+ A=0.75 P=4 MULT=1
MM1013 N_VPWR_M1011_d N_A_183_141#_M1013_g N_X_M1013_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250010 SB=250020
+ A=0.75 P=4 MULT=1
MM1017 N_VPWR_M1017_d N_A_183_141#_M1017_g N_X_M1013_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250010 SB=250020
+ A=0.75 P=4 MULT=1
MM1018 N_VPWR_M1017_d N_A_183_141#_M1018_g N_X_M1018_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250011 SB=250020
+ A=0.75 P=4 MULT=1
MM1020 N_VPWR_M1020_d N_A_183_141#_M1020_g N_X_M1018_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250012 SB=250020
+ A=0.75 P=4 MULT=1
MM1021 N_VPWR_M1020_d N_A_183_141#_M1021_g N_X_M1021_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250013 SB=250020
+ A=0.75 P=4 MULT=1
MM1022 N_VPWR_M1022_d N_A_183_141#_M1022_g N_X_M1021_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250014 SB=250019
+ A=0.75 P=4 MULT=1
MM1023 N_VPWR_M1022_d N_A_183_141#_M1023_g N_X_M1023_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250014 SB=250018
+ A=0.75 P=4 MULT=1
MM1024 N_VPWR_M1024_d N_A_183_141#_M1024_g N_X_M1023_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250015 SB=250017
+ A=0.75 P=4 MULT=1
MM1026 N_VPWR_M1024_d N_A_183_141#_M1026_g N_X_M1026_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250016 SB=250016
+ A=0.75 P=4 MULT=1
MM1029 N_VPWR_M1029_d N_A_183_141#_M1029_g N_X_M1026_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250017 SB=250016
+ A=0.75 P=4 MULT=1
MM1030 N_VPWR_M1029_d N_A_183_141#_M1030_g N_X_M1030_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250017 SB=250015
+ A=0.75 P=4 MULT=1
MM1033 N_VPWR_M1033_d N_A_183_141#_M1033_g N_X_M1030_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250018 SB=250014
+ A=0.75 P=4 MULT=1
MM1034 N_VPWR_M1033_d N_A_183_141#_M1034_g N_X_M1034_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250019 SB=250013
+ A=0.75 P=4 MULT=1
MM1036 N_VPWR_M1036_d N_A_183_141#_M1036_g N_X_M1034_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250012
+ A=0.75 P=4 MULT=1
MM1037 N_VPWR_M1036_d N_A_183_141#_M1037_g N_X_M1037_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250012
+ A=0.75 P=4 MULT=1
MM1041 N_VPWR_M1041_d N_A_183_141#_M1041_g N_X_M1037_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250011
+ A=0.75 P=4 MULT=1
MM1042 N_VPWR_M1041_d N_A_183_141#_M1042_g N_X_M1042_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250010
+ A=0.75 P=4 MULT=1
MM1045 N_VPWR_M1045_d N_A_183_141#_M1045_g N_X_M1042_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250009
+ A=0.75 P=4 MULT=1
MM1046 N_VPWR_M1045_d N_A_183_141#_M1046_g N_X_M1046_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250009
+ A=0.75 P=4 MULT=1
MM1050 N_VPWR_M1050_d N_A_183_141#_M1050_g N_X_M1046_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250008
+ A=0.75 P=4 MULT=1
MM1054 N_VPWR_M1050_d N_A_183_141#_M1054_g N_X_M1054_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250007
+ A=0.75 P=4 MULT=1
MM1055 N_VPWR_M1055_d N_A_183_141#_M1055_g N_X_M1054_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250006
+ A=0.75 P=4 MULT=1
MM1059 N_VPWR_M1055_d N_A_183_141#_M1059_g N_X_M1059_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250005
+ A=0.75 P=4 MULT=1
MM1060 N_VPWR_M1060_d N_A_183_141#_M1060_g N_X_M1059_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250005
+ A=0.75 P=4 MULT=1
MM1063 N_VPWR_M1060_d N_A_183_141#_M1063_g N_X_M1063_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250004
+ A=0.75 P=4 MULT=1
MM1065 N_VPWR_M1065_d N_A_183_141#_M1065_g N_X_M1063_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250003
+ A=0.75 P=4 MULT=1
MM1066 N_VPWR_M1065_d N_A_183_141#_M1066_g N_X_M1066_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250002
+ A=0.75 P=4 MULT=1
MM1073 N_VPWR_M1073_d N_A_183_141#_M1073_g N_X_M1066_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250002
+ A=0.75 P=4 MULT=1
MM1075 N_VPWR_M1073_d N_A_183_141#_M1075_g N_X_M1075_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020 SB=250001
+ A=0.75 P=4 MULT=1
MM1080 N_VPWR_M1080_d N_A_183_141#_M1080_g N_X_M1075_s N_VPB_M1000_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250020
+ SB=250000 A=0.75 P=4 MULT=1
DX84_noxref N_VNB_M1008_b N_VPB_M1000_b NWDIODE A=89.076 P=73.72
*
.include "sky130_fd_sc_hvl__buf_32.pxi.spice"
*
.ends
*
*
