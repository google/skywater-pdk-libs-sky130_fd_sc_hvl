* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1 A SLEEP_B LVPWR VGND VNB VPB VPWR X
*.PININFO A:I SLEEP_B:I LVPWR:I VGND:I VNB:I VPB:I VPWR:I X:O
MM8 X t1 VPB phv m=1 w=0.75 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MM3 t1 t2 VPB phv m=1 w=0.42 l=2.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MI7 isolate_ahv SLEEP_B VPB phv m=1 w=1.5 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 t4 t3 LVPWR phighvt m=1 w=1.12 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 t3 A LVPWR phighvt m=1 w=1.12 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MM4 t2 t1 VPB phv m=1 w=0.42 l=2.0 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MM9 t2 isolate_ahv VNB nhv m=1 w=1.0 l=0.8 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI34 t4 t3 VNB nshort m=1 w=0.74 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MM7 X t1 VNB nhv m=1 w=0.75 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MI16 t2 t3 VNB nhv m=2 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MI15 t1 t4 VNB nhv m=2 w=1.0 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MMIN1 t3 A VNB nshort m=1 w=0.74 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI6 isolate_ahv SLEEP_B VNB nhv m=1 w=0.75 l=0.5 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI23 net54 SLEEP_B VNB nhv m=2 w=5.0 l=0.6 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1
