* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_1528_579# a_1570_457# a_1124_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 a_425_107# SCE a_567_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X2 VGND a_2518_445# a_2789_147# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_2365_445# a_2789_147# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 VGND CLK a_1570_457# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_30_515# SCE VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 a_567_107# a_30_515# a_723_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 VPWR a_2789_147# a_3531_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X8 a_2518_445# a_1570_457# a_2747_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_268_659# a_30_515# a_567_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X10 VPWR CLK a_1570_457# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X11 a_567_107# a_1570_457# a_1124_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X12 VGND SCD a_425_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 a_567_107# D a_581_659# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X14 VGND a_1067_107# a_1454_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 VGND a_3531_107# Q_N VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X16 a_268_659# SCD VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X17 a_1067_107# a_1726_453# a_2518_445# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X18 a_1067_107# a_1124_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X19 a_1124_81# a_1726_453# a_567_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 VPWR a_3531_107# Q_N VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X21 a_1726_453# a_1570_457# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X22 a_723_107# D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X23 Q a_2789_147# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X24 a_1124_81# a_1726_453# a_1454_173# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X25 a_30_515# SCE VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X26 a_1067_107# a_1124_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X27 a_2747_173# a_2789_147# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X28 VGND a_2789_147# a_3531_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X29 VPWR a_2518_445# a_2789_147# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X30 Q a_2789_147# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X31 a_2365_445# a_1726_453# a_2518_445# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X32 a_1726_453# a_1570_457# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X33 VPWR a_1067_107# a_1528_579# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X34 VPWR SCE a_581_659# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X35 a_2518_445# a_1570_457# a_1067_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
.ends
