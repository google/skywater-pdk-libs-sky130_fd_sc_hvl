# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__dfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.80000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.850000 0.810000 4.165000 2.105000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.340000 0.515000 16.690000 3.755000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.045000 0.665000 14.425000 1.495000 ;
        RECT 14.045000 1.495000 14.380000 1.780000 ;
        RECT 14.130000 1.780000 14.380000 3.755000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  2.980000 1.505000  3.665000 2.120000 ;
        RECT  3.495000 0.460000  6.625000 0.630000 ;
        RECT  3.495000 0.630000  3.665000 1.505000 ;
        RECT  6.455000 0.630000  6.625000 1.125000 ;
        RECT  6.455000 1.125000  8.515000 1.295000 ;
        RECT  7.165000 1.825000  8.515000 1.995000 ;
        RECT  8.345000 0.265000 11.075000 0.435000 ;
        RECT  8.345000 0.435000  8.515000 1.125000 ;
        RECT  8.345000 1.295000  8.515000 1.825000 ;
        RECT 10.905000 0.435000 11.075000 0.960000 ;
        RECT 10.905000 0.960000 11.840000 1.130000 ;
        RECT 11.510000 1.130000 11.840000 1.350000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.595000 1.175000 0.925000 1.720000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 16.800000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 16.800000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 16.800000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 16.800000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 17.130000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 16.800000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.800000 0.085000 ;
      RECT  0.000000  3.985000 16.800000 4.155000 ;
      RECT  0.165000  0.495000  0.495000 0.995000 ;
      RECT  0.165000  0.995000  0.415000 2.275000 ;
      RECT  0.165000  2.275000  1.835000 2.445000 ;
      RECT  0.165000  2.445000  0.415000 3.455000 ;
      RECT  0.595000  2.625000  1.485000 3.705000 ;
      RECT  0.675000  0.365000  1.625000 0.995000 ;
      RECT  1.505000  1.900000  1.835000 2.275000 ;
      RECT  1.665000  2.445000  1.835000 3.635000 ;
      RECT  1.665000  3.635000  3.205000 3.805000 ;
      RECT  1.805000  0.495000  2.185000 0.995000 ;
      RECT  2.015000  0.995000  2.185000 1.550000 ;
      RECT  2.015000  1.550000  2.275000 3.455000 ;
      RECT  2.365000  0.365000  3.315000 1.325000 ;
      RECT  2.525000  2.300000  4.515000 2.470000 ;
      RECT  2.525000  2.470000  2.855000 3.420000 ;
      RECT  3.035000  2.650000  3.905000 2.820000 ;
      RECT  3.035000  2.820000  3.205000 3.635000 ;
      RECT  3.385000  3.000000  3.555000 3.705000 ;
      RECT  3.735000  2.820000  3.905000 3.600000 ;
      RECT  3.735000  3.600000  5.565000 3.770000 ;
      RECT  4.085000  3.000000  4.515000 3.420000 ;
      RECT  4.345000  0.825000  4.655000 1.325000 ;
      RECT  4.345000  1.325000  4.515000 2.300000 ;
      RECT  4.345000  2.470000  4.515000 3.000000 ;
      RECT  4.695000  1.505000  5.925000 1.780000 ;
      RECT  4.695000  1.780000  4.865000 2.820000 ;
      RECT  4.865000  3.000000  5.215000 3.420000 ;
      RECT  5.045000  2.200000  6.275000 2.370000 ;
      RECT  5.045000  2.370000  5.215000 3.000000 ;
      RECT  5.270000  0.825000  5.600000 1.155000 ;
      RECT  5.270000  1.155000  6.275000 1.325000 ;
      RECT  5.395000  2.550000  5.650000 2.875000 ;
      RECT  5.395000  2.875000  7.035000 3.045000 ;
      RECT  5.395000  3.045000  5.565000 3.600000 ;
      RECT  5.595000  1.780000  5.925000 2.020000 ;
      RECT  5.745000  3.225000  6.685000 3.705000 ;
      RECT  6.105000  1.325000  6.275000 1.475000 ;
      RECT  6.105000  1.475000  8.165000 1.645000 ;
      RECT  6.105000  1.645000  6.275000 2.200000 ;
      RECT  6.105000  2.370000  6.275000 2.525000 ;
      RECT  6.105000  2.525000  7.385000 2.695000 ;
      RECT  6.455000  1.825000  6.785000 2.175000 ;
      RECT  6.455000  2.175000  9.025000 2.345000 ;
      RECT  6.865000  3.045000  7.035000 3.635000 ;
      RECT  6.865000  3.635000  7.735000 3.805000 ;
      RECT  7.215000  0.365000  8.165000 0.945000 ;
      RECT  7.215000  2.695000  7.385000 3.455000 ;
      RECT  7.565000  2.700000  9.375000 2.870000 ;
      RECT  7.565000  2.870000  7.735000 3.635000 ;
      RECT  7.915000  3.050000  8.865000 3.705000 ;
      RECT  8.695000  0.615000  9.025000 2.175000 ;
      RECT  8.695000  2.345000  9.025000 2.520000 ;
      RECT  9.205000  1.230000 10.375000 1.400000 ;
      RECT  9.205000  1.400000  9.375000 2.700000 ;
      RECT  9.555000  2.270000 10.410000 2.440000 ;
      RECT  9.555000  2.440000  9.805000 3.350000 ;
      RECT  9.580000  0.615000 10.725000 0.785000 ;
      RECT  9.580000  0.785000  9.910000 0.995000 ;
      RECT  9.725000  1.580000 10.060000 2.090000 ;
      RECT 10.090000  1.070000 10.375000 1.230000 ;
      RECT 10.240000  2.000000 12.530000 2.170000 ;
      RECT 10.240000  2.170000 10.410000 2.270000 ;
      RECT 10.555000  0.785000 10.725000 2.000000 ;
      RECT 10.590000  2.350000 11.540000 3.705000 ;
      RECT 10.930000  1.310000 11.260000 1.530000 ;
      RECT 10.930000  1.530000 12.880000 1.700000 ;
      RECT 10.930000  1.700000 11.260000 1.820000 ;
      RECT 11.255000  0.365000 12.205000 0.780000 ;
      RECT 11.965000  2.350000 12.880000 2.520000 ;
      RECT 11.965000  2.520000 12.295000 2.770000 ;
      RECT 12.200000  1.880000 12.530000 2.000000 ;
      RECT 12.710000  0.515000 13.075000 0.975000 ;
      RECT 12.710000  0.975000 12.880000 1.530000 ;
      RECT 12.710000  1.700000 12.880000 2.350000 ;
      RECT 13.060000  2.175000 13.950000 3.755000 ;
      RECT 13.255000  0.365000 13.845000 1.495000 ;
      RECT 14.665000  0.825000 15.015000 1.505000 ;
      RECT 14.665000  1.505000 16.160000 1.835000 ;
      RECT 14.665000  1.835000 14.995000 3.005000 ;
      RECT 15.175000  2.175000 16.125000 3.755000 ;
      RECT 15.195000  0.365000 16.145000 1.325000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.595000  3.505000  0.765000 3.675000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.705000  0.395000  0.875000 0.565000 ;
      RECT  0.955000  3.505000  1.125000 3.675000 ;
      RECT  1.065000  0.395000  1.235000 0.565000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.315000  3.505000  1.485000 3.675000 ;
      RECT  1.425000  0.395000  1.595000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  1.580000  2.245000 1.750000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.395000  0.395000  2.565000 0.565000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.755000  0.395000  2.925000 0.565000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.115000  0.395000  3.285000 0.565000 ;
      RECT  3.385000  3.505000  3.555000 3.675000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.580000  5.125000 1.750000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.770000  3.505000  5.940000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.130000  3.505000  6.300000 3.675000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.490000  3.505000  6.660000 3.675000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.245000  0.395000  7.415000 0.565000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.605000  0.395000  7.775000 0.565000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  7.945000  3.505000  8.115000 3.675000 ;
      RECT  7.965000  0.395000  8.135000 0.565000 ;
      RECT  8.305000  3.505000  8.475000 3.675000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.665000  3.505000  8.835000 3.675000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  1.580000  9.925000 1.750000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.620000  3.505000 10.790000 3.675000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.980000  3.505000 11.150000 3.675000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.285000  0.395000 11.455000 0.565000 ;
      RECT 11.340000  3.505000 11.510000 3.675000 ;
      RECT 11.645000  0.395000 11.815000 0.565000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.005000  0.395000 12.175000 0.565000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 13.060000  3.505000 13.230000 3.675000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.285000  0.395000 13.455000 0.565000 ;
      RECT 13.420000  3.505000 13.590000 3.675000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.645000  0.395000 13.815000 0.565000 ;
      RECT 13.780000  3.505000 13.950000 3.675000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.205000  3.505000 15.375000 3.675000 ;
      RECT 15.225000  0.395000 15.395000 0.565000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.565000  3.505000 15.735000 3.675000 ;
      RECT 15.585000  0.395000 15.755000 0.565000 ;
      RECT 15.925000  3.505000 16.095000 3.675000 ;
      RECT 15.945000  0.395000 16.115000 0.565000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
    LAYER met1 ;
      RECT 2.015000 1.550000 2.305000 1.595000 ;
      RECT 2.015000 1.595000 9.985000 1.735000 ;
      RECT 2.015000 1.735000 2.305000 1.780000 ;
      RECT 4.895000 1.550000 5.185000 1.595000 ;
      RECT 4.895000 1.735000 5.185000 1.780000 ;
      RECT 9.695000 1.550000 9.985000 1.595000 ;
      RECT 9.695000 1.735000 9.985000 1.780000 ;
  END
END sky130_fd_sc_hvl__dfrbp_1
END LIBRARY
