* File: sky130_fd_sc_hvl__einvn_1.spice
* Created: Fri Aug 28 09:35:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__einvn_1.pex.spice"
.subckt sky130_fd_sc_hvl__einvn_1  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_TE_B_M1001_g N_A_30_173#_M1001_s N_VNB_M1001_b NHV L=0.5
+ W=0.42 AD=0.190131 AS=0.1113 PD=1.09128 PS=1.37 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1002 A_437_107# N_A_30_173#_M1002_g N_VGND_M1001_d N_VNB_M1001_b NHV L=0.5
+ W=0.75 AD=0.07875 AS=0.339519 PD=0.96 PS=1.94872 NRD=7.5924 NRS=0 M=1 R=1.5
+ SA=250001 SB=250001 A=0.375 P=2.5 MULT=1
MM1003 N_Z_M1003_d N_A_M1003_g A_437_107# N_VNB_M1001_b NHV L=0.5 W=0.75
+ AD=0.21375 AS=0.07875 PD=2.07 PS=0.96 NRD=0 NRS=7.5924 M=1 R=1.5 SA=250002
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_TE_B_M1005_g N_A_30_173#_M1005_s N_VPB_M1005_b PHV L=0.5
+ W=0.75 AD=0.221933 AS=0.21375 PD=1.37 PS=2.07 NRD=57.2809 NRS=0 M=1 R=1.5
+ SA=250000 SB=250002 A=0.375 P=2.5 MULT=1
MM1004 A_413_443# N_TE_B_M1004_g N_VPWR_M1005_d N_VPB_M1005_b PHV L=0.5 W=1.5
+ AD=0.2475 AS=0.443867 PD=1.83 PS=2.74 NRD=14.0003 NRS=6.3603 M=1 R=3 SA=250001
+ SB=250001 A=0.75 P=4 MULT=1
MM1000 N_Z_M1000_d N_A_M1000_g A_413_443# N_VPB_M1005_b PHV L=0.5 W=1.5
+ AD=0.4275 AS=0.2475 PD=3.57 PS=1.83 NRD=0 NRS=14.0003 M=1 R=3 SA=250001
+ SB=250000 A=0.75 P=4 MULT=1
DX6_noxref N_VNB_M1001_b N_VPB_M1005_b NWDIODE A=10.452 P=13.24
*
.include "sky130_fd_sc_hvl__einvn_1.pxi.spice"
*
.ends
*
*
