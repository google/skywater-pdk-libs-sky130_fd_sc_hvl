* File: sky130_fd_sc_hvl__buf_16.pex.spice
* Created: Fri Aug 28 09:32:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__BUF_16%VNB 5 7 17 26
r89 17 26 5.23549 $w=2.3e-07 $l=8.16e-06 $layer=MET1_cond $X=17.52 $Y=0 $X2=9.36
+ $Y2=0
r90 7 26 0.30797 $w=2.3e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r91 7 11 5.54346 $w=2.3e-07 $l=8.64e-06 $layer=MET1_cond $X=8.88 $Y=0 $X2=0.24
+ $Y2=0
r92 5 17 0.502703 $w=1.7e-07 $l=3.145e-06 $layer=mcon $count=18 $X=17.52 $Y=0
+ $X2=17.52 $Y2=0
r93 5 11 0.502703 $w=1.7e-07 $l=3.145e-06 $layer=mcon $count=18 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_16%VPB 4 6 14 15 23
r137 15 23 5.23549 $w=2.3e-07 $l=8.16e-06 $layer=MET1_cond $X=17.52 $Y=4.07
+ $X2=9.36 $Y2=4.07
r138 14 15 0.502703 $w=1.7e-07 $l=3.145e-06 $layer=mcon $count=18 $X=17.52
+ $Y=4.07 $X2=17.52 $Y2=4.07
r139 9 14 1127.36 $w=1.68e-07 $l=1.728e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=17.52 $Y2=4.07
r140 9 10 0.502703 $w=1.7e-07 $l=3.145e-06 $layer=mcon $count=18 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r141 6 23 0.30797 $w=2.3e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=4.07
+ $X2=9.36 $Y2=4.07
r142 6 10 5.54346 $w=2.3e-07 $l=8.64e-06 $layer=MET1_cond $X=8.88 $Y=4.07
+ $X2=0.24 $Y2=4.07
r143 4 14 9.83784 $w=1.7e-07 $l=1.75624e-05 $layer=licon1_NTAP_notbjt $count=18
+ $X=0 $Y=3.985 $X2=17.52 $Y2=4.07
r144 4 9 9.83784 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=18
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_16%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34
+ 36 38 41 43 44 45 46 47 48 49 68 69
c132 68 0 1.42377e-19 $X=4.465 $Y=1.73
c133 13 0 3.19988e-20 $X=1.445 $Y=2.965
r134 67 69 10.7006 $w=5e-07 $l=1e-07 $layer=POLY_cond $X=4.465 $Y=1.815
+ $X2=4.565 $Y2=1.815
r135 67 68 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6 $X=4.465
+ $Y=1.73 $X2=4.465 $Y2=1.73
r136 65 67 72.764 $w=5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.785 $Y=1.815
+ $X2=4.465 $Y2=1.815
r137 64 65 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.005 $Y=1.815
+ $X2=3.785 $Y2=1.815
r138 63 64 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.225 $Y=1.815
+ $X2=3.005 $Y2=1.815
r139 62 63 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.445 $Y=1.815
+ $X2=2.225 $Y2=1.815
r140 61 62 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.665 $Y=1.815
+ $X2=1.445 $Y2=1.815
r141 58 61 29.9617 $w=5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.385 $Y=1.815
+ $X2=0.665 $Y2=1.815
r142 58 59 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6 $X=0.385
+ $Y=1.73 $X2=0.385 $Y2=1.73
r143 49 68 42.4197 $w=2.33e-07 $l=8.65e-07 $layer=LI1_cond $X=3.6 $Y=1.697
+ $X2=4.465 $Y2=1.697
r144 48 49 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.697
+ $X2=3.6 $Y2=1.697
r145 47 48 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.697
+ $X2=3.12 $Y2=1.697
r146 46 47 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.697
+ $X2=2.64 $Y2=1.697
r147 45 46 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.697
+ $X2=2.16 $Y2=1.697
r148 44 45 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.697
+ $X2=1.68 $Y2=1.697
r149 43 44 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.697
+ $X2=1.2 $Y2=1.697
r150 43 59 16.4284 $w=2.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.72 $Y=1.697
+ $X2=0.385 $Y2=1.697
r151 39 69 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.565 $Y=2.065
+ $X2=4.565 $Y2=1.815
r152 39 41 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=4.565 $Y=2.065
+ $X2=4.565 $Y2=2.965
r153 36 69 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.565 $Y=1.565
+ $X2=4.565 $Y2=1.815
r154 36 38 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.565 $Y=1.565
+ $X2=4.565 $Y2=1.08
r155 32 65 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.785 $Y=2.065
+ $X2=3.785 $Y2=1.815
r156 32 34 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=3.785 $Y=2.065
+ $X2=3.785 $Y2=2.965
r157 29 65 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.785 $Y=1.565
+ $X2=3.785 $Y2=1.815
r158 29 31 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.785 $Y=1.565
+ $X2=3.785 $Y2=1.08
r159 25 64 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.005 $Y=2.065
+ $X2=3.005 $Y2=1.815
r160 25 27 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=3.005 $Y=2.065
+ $X2=3.005 $Y2=2.965
r161 22 64 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.005 $Y=1.565
+ $X2=3.005 $Y2=1.815
r162 22 24 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.005 $Y=1.565
+ $X2=3.005 $Y2=1.08
r163 18 63 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.225 $Y=2.065
+ $X2=2.225 $Y2=1.815
r164 18 20 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=2.225 $Y=2.065
+ $X2=2.225 $Y2=2.965
r165 15 63 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.225 $Y=1.565
+ $X2=2.225 $Y2=1.815
r166 15 17 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.225 $Y=1.565
+ $X2=2.225 $Y2=1.08
r167 11 62 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.445 $Y=2.065
+ $X2=1.445 $Y2=1.815
r168 11 13 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=1.445 $Y=2.065
+ $X2=1.445 $Y2=2.965
r169 8 62 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.445 $Y=1.565
+ $X2=1.445 $Y2=1.815
r170 8 10 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.445 $Y=1.565
+ $X2=1.445 $Y2=1.08
r171 4 61 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.665 $Y=2.065
+ $X2=0.665 $Y2=1.815
r172 4 6 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=0.665 $Y=2.065 $X2=0.665
+ $Y2=2.965
r173 1 61 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.665 $Y=1.565
+ $X2=0.665 $Y2=1.815
r174 1 3 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.665 $Y=1.565
+ $X2=0.665 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_16%A_183_141# 1 2 3 4 5 6 19 21 24 26 28 31 33
+ 35 38 40 42 45 47 49 52 54 56 59 61 63 66 68 70 73 75 77 80 82 84 87 89 91 94
+ 96 98 101 103 105 108 110 112 115 117 119 122 124 126 129 133 137 141 142 143
+ 144 147 151 155 157 161 167 169 171 173 174 175 176 181 182 183 184 187 188
+ 189 190 191 194 195 196 197 198 201 202 203 204 205 208 209 210 211 212 215
+ 216 217 218 219 222 223 224 226 228 229 231 232
c482 124 0 1.42377e-19 $X=17.045 $Y=1.565
r483 231 232 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.245 $Y=1.665
+ $X2=5.245 $Y2=1.665
r484 229 268 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=16.025
+ $Y=1.73 $X2=16.025 $Y2=1.73
r485 228 229 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.035 $Y=1.665
+ $X2=16.035 $Y2=1.665
r486 226 228 0.250226 $w=2.3e-07 $l=3.9e-07 $layer=MET1_cond $X=15.645 $Y=1.665
+ $X2=16.035 $Y2=1.665
r487 223 226 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=15.53 $Y=1.665
+ $X2=15.645 $Y2=1.665
r488 223 224 0.876223 $w=1.7e-07 $l=9.1e-07 $layer=MET1_cond $X=15.53 $Y=1.665
+ $X2=14.62 $Y2=1.665
r489 222 263 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.465
+ $Y=1.73 $X2=14.465 $Y2=1.73
r490 221 222 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.475 $Y=1.665
+ $X2=14.475 $Y2=1.665
r491 219 221 0.250226 $w=2.3e-07 $l=3.9e-07 $layer=MET1_cond $X=14.085 $Y=1.665
+ $X2=14.475 $Y2=1.665
r492 218 224 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=14.505
+ $Y=1.665 $X2=14.62 $Y2=1.665
r493 218 221 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=14.505 $Y=1.665
+ $X2=14.475 $Y2=1.665
r494 216 219 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=13.97 $Y=1.665
+ $X2=14.085 $Y2=1.665
r495 216 217 0.876223 $w=1.7e-07 $l=9.1e-07 $layer=MET1_cond $X=13.97 $Y=1.665
+ $X2=13.06 $Y2=1.665
r496 215 258 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.905
+ $Y=1.73 $X2=12.905 $Y2=1.73
r497 214 215 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.915 $Y=1.665
+ $X2=12.915 $Y2=1.665
r498 212 214 0.250226 $w=2.3e-07 $l=3.9e-07 $layer=MET1_cond $X=12.525 $Y=1.665
+ $X2=12.915 $Y2=1.665
r499 211 217 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=12.945
+ $Y=1.665 $X2=13.06 $Y2=1.665
r500 211 214 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=12.945 $Y=1.665
+ $X2=12.915 $Y2=1.665
r501 209 212 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=12.41 $Y=1.665
+ $X2=12.525 $Y2=1.665
r502 209 210 0.876223 $w=1.7e-07 $l=9.1e-07 $layer=MET1_cond $X=12.41 $Y=1.665
+ $X2=11.5 $Y2=1.665
r503 208 253 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.345
+ $Y=1.73 $X2=11.345 $Y2=1.73
r504 207 208 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.355 $Y=1.665
+ $X2=11.355 $Y2=1.665
r505 205 207 0.250226 $w=2.3e-07 $l=3.9e-07 $layer=MET1_cond $X=10.965 $Y=1.665
+ $X2=11.355 $Y2=1.665
r506 204 210 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=11.385
+ $Y=1.665 $X2=11.5 $Y2=1.665
r507 204 207 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=11.385 $Y=1.665
+ $X2=11.355 $Y2=1.665
r508 202 205 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=10.85 $Y=1.665
+ $X2=10.965 $Y2=1.665
r509 202 203 0.876223 $w=1.7e-07 $l=9.1e-07 $layer=MET1_cond $X=10.85 $Y=1.665
+ $X2=9.94 $Y2=1.665
r510 201 248 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.785
+ $Y=1.73 $X2=9.785 $Y2=1.73
r511 200 201 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.795 $Y=1.665
+ $X2=9.795 $Y2=1.665
r512 198 200 0.250226 $w=2.3e-07 $l=3.9e-07 $layer=MET1_cond $X=9.405 $Y=1.665
+ $X2=9.795 $Y2=1.665
r513 197 203 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=9.825 $Y=1.665
+ $X2=9.94 $Y2=1.665
r514 197 200 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=9.825 $Y=1.665
+ $X2=9.795 $Y2=1.665
r515 195 198 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=9.29 $Y=1.665
+ $X2=9.405 $Y2=1.665
r516 195 196 0.876223 $w=1.7e-07 $l=9.1e-07 $layer=MET1_cond $X=9.29 $Y=1.665
+ $X2=8.38 $Y2=1.665
r517 194 243 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.225
+ $Y=1.73 $X2=8.225 $Y2=1.73
r518 193 194 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.235 $Y=1.665
+ $X2=8.235 $Y2=1.665
r519 191 193 0.250226 $w=2.3e-07 $l=3.9e-07 $layer=MET1_cond $X=7.845 $Y=1.665
+ $X2=8.235 $Y2=1.665
r520 190 196 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=8.265 $Y=1.665
+ $X2=8.38 $Y2=1.665
r521 190 193 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=8.265 $Y=1.665
+ $X2=8.235 $Y2=1.665
r522 188 191 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=7.73 $Y=1.665
+ $X2=7.845 $Y2=1.665
r523 188 189 0.876223 $w=1.7e-07 $l=9.1e-07 $layer=MET1_cond $X=7.73 $Y=1.665
+ $X2=6.82 $Y2=1.665
r524 187 238 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.665
+ $Y=1.73 $X2=6.665 $Y2=1.73
r525 186 187 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.675 $Y=1.665
+ $X2=6.675 $Y2=1.665
r526 184 186 0.250226 $w=2.3e-07 $l=3.9e-07 $layer=MET1_cond $X=6.285 $Y=1.665
+ $X2=6.675 $Y2=1.665
r527 183 189 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=6.705 $Y=1.665
+ $X2=6.82 $Y2=1.665
r528 183 186 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=6.705 $Y=1.665
+ $X2=6.675 $Y2=1.665
r529 182 231 0.0841272 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=5.36 $Y=1.665
+ $X2=5.245 $Y2=1.665
r530 181 184 0.0789558 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=6.17 $Y=1.665
+ $X2=6.285 $Y2=1.665
r531 181 182 0.779935 $w=1.7e-07 $l=8.1e-07 $layer=MET1_cond $X=6.17 $Y=1.665
+ $X2=5.36 $Y2=1.665
r532 178 232 6.959 $w=5.48e-07 $l=3.2e-07 $layer=LI1_cond $X=5.075 $Y=1.985
+ $X2=5.075 $Y2=1.665
r533 177 232 5.54545 $w=5.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.075 $Y=1.41
+ $X2=5.075 $Y2=1.665
r534 172 175 6.19399 $w=2.8e-07 $l=1.75e-07 $layer=LI1_cond $X=4.29 $Y=2.125
+ $X2=4.115 $Y2=2.125
r535 171 178 7.79946 $w=2.8e-07 $l=3.37824e-07 $layer=LI1_cond $X=4.8 $Y=2.125
+ $X2=5.075 $Y2=1.985
r536 171 172 20.9909 $w=2.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.8 $Y=2.125
+ $X2=4.29 $Y2=2.125
r537 170 176 5.75112 $w=2.15e-07 $l=1.23e-07 $layer=LI1_cond $X=4.27 $Y=1.302
+ $X2=4.147 $Y2=1.302
r538 169 177 8.67418 $w=2.15e-07 $l=3.24538e-07 $layer=LI1_cond $X=4.8 $Y=1.302
+ $X2=5.075 $Y2=1.41
r539 169 170 28.4091 $w=2.13e-07 $l=5.3e-07 $layer=LI1_cond $X=4.8 $Y=1.302
+ $X2=4.27 $Y2=1.302
r540 165 176 0.876697 $w=2.45e-07 $l=1.07e-07 $layer=LI1_cond $X=4.147 $Y=1.195
+ $X2=4.147 $Y2=1.302
r541 165 167 14.1115 $w=2.43e-07 $l=3e-07 $layer=LI1_cond $X=4.147 $Y=1.195
+ $X2=4.147 $Y2=0.895
r542 161 163 41.1587 $w=3.48e-07 $l=1.25e-06 $layer=LI1_cond $X=4.115 $Y=2.34
+ $X2=4.115 $Y2=3.59
r543 159 175 0.552779 $w=3.5e-07 $l=1.4e-07 $layer=LI1_cond $X=4.115 $Y=2.265
+ $X2=4.115 $Y2=2.125
r544 159 161 2.46952 $w=3.48e-07 $l=7.5e-08 $layer=LI1_cond $X=4.115 $Y=2.265
+ $X2=4.115 $Y2=2.34
r545 158 173 8.20698 $w=2.15e-07 $l=1.95e-07 $layer=LI1_cond $X=2.79 $Y=1.302
+ $X2=2.595 $Y2=1.302
r546 157 176 5.75112 $w=2.15e-07 $l=1.22e-07 $layer=LI1_cond $X=4.025 $Y=1.302
+ $X2=4.147 $Y2=1.302
r547 157 158 66.1985 $w=2.13e-07 $l=1.235e-06 $layer=LI1_cond $X=4.025 $Y=1.302
+ $X2=2.79 $Y2=1.302
r548 156 174 5.6179 $w=2.8e-07 $l=1.55e-07 $layer=LI1_cond $X=2.71 $Y=2.125
+ $X2=2.555 $Y2=2.125
r549 155 175 6.19399 $w=2.8e-07 $l=1.75e-07 $layer=LI1_cond $X=3.94 $Y=2.125
+ $X2=4.115 $Y2=2.125
r550 155 156 50.6252 $w=2.78e-07 $l=1.23e-06 $layer=LI1_cond $X=3.94 $Y=2.125
+ $X2=2.71 $Y2=2.125
r551 151 153 46.4695 $w=3.08e-07 $l=1.25e-06 $layer=LI1_cond $X=2.555 $Y=2.34
+ $X2=2.555 $Y2=3.59
r552 149 174 0.978733 $w=3.1e-07 $l=1.4e-07 $layer=LI1_cond $X=2.555 $Y=2.265
+ $X2=2.555 $Y2=2.125
r553 149 151 2.78817 $w=3.08e-07 $l=7.5e-08 $layer=LI1_cond $X=2.555 $Y=2.265
+ $X2=2.555 $Y2=2.34
r554 145 173 0.684683 $w=3.9e-07 $l=1.07e-07 $layer=LI1_cond $X=2.595 $Y=1.195
+ $X2=2.595 $Y2=1.302
r555 145 147 8.86495 $w=3.88e-07 $l=3e-07 $layer=LI1_cond $X=2.595 $Y=1.195
+ $X2=2.595 $Y2=0.895
r556 143 173 8.20698 $w=2.15e-07 $l=1.95e-07 $layer=LI1_cond $X=2.4 $Y=1.302
+ $X2=2.595 $Y2=1.302
r557 143 144 65.9305 $w=2.13e-07 $l=1.23e-06 $layer=LI1_cond $X=2.4 $Y=1.302
+ $X2=1.17 $Y2=1.302
r558 141 174 5.6179 $w=2.8e-07 $l=1.55e-07 $layer=LI1_cond $X=2.4 $Y=2.125
+ $X2=2.555 $Y2=2.125
r559 141 142 51.0368 $w=2.78e-07 $l=1.24e-06 $layer=LI1_cond $X=2.4 $Y=2.125
+ $X2=1.16 $Y2=2.125
r560 137 139 46.4695 $w=3.08e-07 $l=1.25e-06 $layer=LI1_cond $X=1.005 $Y=2.34
+ $X2=1.005 $Y2=3.59
r561 135 142 6.83944 $w=2.8e-07 $l=2.13834e-07 $layer=LI1_cond $X=1.005 $Y=2.265
+ $X2=1.16 $Y2=2.125
r562 135 137 2.78817 $w=3.08e-07 $l=7.5e-08 $layer=LI1_cond $X=1.005 $Y=2.265
+ $X2=1.005 $Y2=2.34
r563 131 144 7.36541 $w=2.15e-07 $l=2.25233e-07 $layer=LI1_cond $X=0.992
+ $Y=1.195 $X2=1.17 $Y2=1.302
r564 131 133 8.92738 $w=3.53e-07 $l=2.75e-07 $layer=LI1_cond $X=0.992 $Y=1.195
+ $X2=0.992 $Y2=0.92
r565 124 129 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=17.045 $Y=2.005
+ $X2=17.045 $Y2=2.965
r566 124 126 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=17.045 $Y=1.565
+ $X2=17.045 $Y2=1.08
r567 117 124 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=16.265 $Y=1.785
+ $X2=17.045 $Y2=1.785
r568 117 268 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=16.265 $Y=1.785
+ $X2=16.025 $Y2=1.785
r569 117 122 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=16.265 $Y=2.005
+ $X2=16.265 $Y2=2.965
r570 117 119 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=16.265 $Y=1.565
+ $X2=16.265 $Y2=1.08
r571 110 268 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=15.485 $Y=1.785
+ $X2=16.025 $Y2=1.785
r572 110 115 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=15.485 $Y=2.005
+ $X2=15.485 $Y2=2.965
r573 110 112 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=15.485 $Y=1.565
+ $X2=15.485 $Y2=1.08
r574 103 110 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=14.705 $Y=1.785
+ $X2=15.485 $Y2=1.785
r575 103 263 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=14.705 $Y=1.785
+ $X2=14.465 $Y2=1.785
r576 103 108 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=14.705 $Y=2.005
+ $X2=14.705 $Y2=2.965
r577 103 105 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=14.705 $Y=1.565
+ $X2=14.705 $Y2=1.08
r578 96 263 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=13.925 $Y=1.785
+ $X2=14.465 $Y2=1.785
r579 96 101 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=13.925 $Y=2.005
+ $X2=13.925 $Y2=2.965
r580 96 98 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=13.925 $Y=1.565
+ $X2=13.925 $Y2=1.08
r581 89 96 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=13.145 $Y=1.785
+ $X2=13.925 $Y2=1.785
r582 89 258 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=13.145 $Y=1.785
+ $X2=12.905 $Y2=1.785
r583 89 94 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=13.145 $Y=2.005
+ $X2=13.145 $Y2=2.965
r584 89 91 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=13.145 $Y=1.565
+ $X2=13.145 $Y2=1.08
r585 82 258 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=12.365 $Y=1.785
+ $X2=12.905 $Y2=1.785
r586 82 87 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=12.365 $Y=2.005
+ $X2=12.365 $Y2=2.965
r587 82 84 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=12.365 $Y=1.565
+ $X2=12.365 $Y2=1.08
r588 75 82 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=11.585 $Y=1.785
+ $X2=12.365 $Y2=1.785
r589 75 253 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=11.585 $Y=1.785
+ $X2=11.345 $Y2=1.785
r590 75 80 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=11.585 $Y=2.005
+ $X2=11.585 $Y2=2.965
r591 75 77 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.585 $Y=1.565
+ $X2=11.585 $Y2=1.08
r592 68 253 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=10.805 $Y=1.785
+ $X2=11.345 $Y2=1.785
r593 68 73 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=10.805 $Y=2.005
+ $X2=10.805 $Y2=2.965
r594 68 70 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=10.805 $Y=1.565
+ $X2=10.805 $Y2=1.08
r595 61 68 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=10.025 $Y=1.785
+ $X2=10.805 $Y2=1.785
r596 61 248 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=10.025 $Y=1.785
+ $X2=9.785 $Y2=1.785
r597 61 66 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=10.025 $Y=2.005
+ $X2=10.025 $Y2=2.965
r598 61 63 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=10.025 $Y=1.565
+ $X2=10.025 $Y2=1.08
r599 54 248 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=9.245 $Y=1.785
+ $X2=9.785 $Y2=1.785
r600 54 59 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=9.245 $Y=2.005
+ $X2=9.245 $Y2=2.965
r601 54 56 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.245 $Y=1.565
+ $X2=9.245 $Y2=1.08
r602 47 54 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=8.465 $Y=1.785
+ $X2=9.245 $Y2=1.785
r603 47 243 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=8.465 $Y=1.785
+ $X2=8.225 $Y2=1.785
r604 47 52 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=8.465 $Y=2.005
+ $X2=8.465 $Y2=2.965
r605 47 49 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=8.465 $Y=1.565
+ $X2=8.465 $Y2=1.08
r606 40 243 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=7.685 $Y=1.785
+ $X2=8.225 $Y2=1.785
r607 40 45 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=7.685 $Y=2.005
+ $X2=7.685 $Y2=2.965
r608 40 42 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.685 $Y=1.565
+ $X2=7.685 $Y2=1.08
r609 33 40 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=6.905 $Y=1.785
+ $X2=7.685 $Y2=1.785
r610 33 238 30.3357 $w=4.4e-07 $l=2.4e-07 $layer=POLY_cond $X=6.905 $Y=1.785
+ $X2=6.665 $Y2=1.785
r611 33 38 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=6.905 $Y=2.005
+ $X2=6.905 $Y2=2.965
r612 33 35 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.905 $Y=1.565
+ $X2=6.905 $Y2=1.08
r613 26 238 68.2552 $w=4.4e-07 $l=5.4e-07 $layer=POLY_cond $X=6.125 $Y=1.785
+ $X2=6.665 $Y2=1.785
r614 26 31 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=6.125 $Y=2.005
+ $X2=6.125 $Y2=2.965
r615 26 28 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.125 $Y=1.565
+ $X2=6.125 $Y2=1.08
r616 19 26 98.5909 $w=4.4e-07 $l=7.8e-07 $layer=POLY_cond $X=5.345 $Y=1.785
+ $X2=6.125 $Y2=1.785
r617 19 24 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=5.345 $Y=2.005
+ $X2=5.345 $Y2=2.965
r618 19 21 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=5.345 $Y=1.565
+ $X2=5.345 $Y2=1.08
r619 6 163 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=4.035
+ $Y=2.215 $X2=4.175 $Y2=3.59
r620 6 161 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.035
+ $Y=2.215 $X2=4.175 $Y2=2.34
r621 5 153 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.475
+ $Y=2.215 $X2=2.615 $Y2=3.59
r622 5 151 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.475
+ $Y=2.215 $X2=2.615 $Y2=2.34
r623 4 139 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=0.915
+ $Y=2.215 $X2=1.055 $Y2=3.59
r624 4 137 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.915
+ $Y=2.215 $X2=1.055 $Y2=2.34
r625 3 167 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=4.035
+ $Y=0.705 $X2=4.175 $Y2=0.895
r626 2 147 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=2.475
+ $Y=0.705 $X2=2.615 $Y2=0.895
r627 1 133 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=0.915
+ $Y=0.705 $X2=1.055 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 37 40 49 60
+ 71 82 93 104 115 126 137 148 159 163
c205 40 0 3.19988e-20 $X=0.275 $Y=2.36
r206 162 163 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.515 $Y=3.56
+ $X2=17.515 $Y2=3.56
r207 159 162 27.081 $w=5.28e-07 $l=1.2e-06 $layer=LI1_cond $X=17.335 $Y=2.36
+ $X2=17.335 $Y2=3.56
r208 154 163 0.491399 $w=3.7e-07 $l=1.28e-06 $layer=MET1_cond $X=16.235 $Y=3.63
+ $X2=17.515 $Y2=3.63
r209 152 154 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=15.515 $Y=3.63
+ $X2=16.235 $Y2=3.63
r210 151 156 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=15.875 $Y=3.56
+ $X2=15.875 $Y2=3.59
r211 151 154 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.235 $Y=3.56
+ $X2=16.235 $Y2=3.56
r212 151 152 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.515 $Y=3.56
+ $X2=15.515 $Y2=3.56
r213 148 151 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=15.875 $Y=2.34
+ $X2=15.875 $Y2=3.56
r214 143 152 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=14.675 $Y=3.63
+ $X2=15.515 $Y2=3.63
r215 141 143 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=13.955 $Y=3.63
+ $X2=14.675 $Y2=3.63
r216 140 145 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=14.315 $Y=3.56
+ $X2=14.315 $Y2=3.59
r217 140 143 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.675 $Y=3.56
+ $X2=14.675 $Y2=3.56
r218 140 141 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.955 $Y=3.56
+ $X2=13.955 $Y2=3.56
r219 137 140 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=14.315 $Y=2.34
+ $X2=14.315 $Y2=3.56
r220 132 141 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=13.115 $Y=3.63
+ $X2=13.955 $Y2=3.63
r221 130 132 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=12.395 $Y=3.63
+ $X2=13.115 $Y2=3.63
r222 129 134 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=12.755 $Y=3.56
+ $X2=12.755 $Y2=3.59
r223 129 132 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.115 $Y=3.56
+ $X2=13.115 $Y2=3.56
r224 129 130 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.395 $Y=3.56
+ $X2=12.395 $Y2=3.56
r225 126 129 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=12.755 $Y=2.34
+ $X2=12.755 $Y2=3.56
r226 121 130 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=11.555 $Y=3.63
+ $X2=12.395 $Y2=3.63
r227 119 121 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.835 $Y=3.63
+ $X2=11.555 $Y2=3.63
r228 118 123 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=11.195 $Y=3.56
+ $X2=11.195 $Y2=3.59
r229 118 121 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.555 $Y=3.56
+ $X2=11.555 $Y2=3.56
r230 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.835 $Y=3.56
+ $X2=10.835 $Y2=3.56
r231 115 118 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=11.195 $Y=2.34
+ $X2=11.195 $Y2=3.56
r232 110 119 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=9.995 $Y=3.63
+ $X2=10.835 $Y2=3.63
r233 108 110 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=9.275 $Y=3.63
+ $X2=9.995 $Y2=3.63
r234 107 112 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=9.635 $Y=3.56
+ $X2=9.635 $Y2=3.59
r235 107 110 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.995 $Y=3.56
+ $X2=9.995 $Y2=3.56
r236 107 108 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.275 $Y=3.56
+ $X2=9.275 $Y2=3.56
r237 104 107 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=9.635 $Y=2.34
+ $X2=9.635 $Y2=3.56
r238 97 99 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.715 $Y=3.63
+ $X2=8.435 $Y2=3.63
r239 96 101 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=8.075 $Y=3.56
+ $X2=8.075 $Y2=3.59
r240 96 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.435 $Y=3.56
+ $X2=8.435 $Y2=3.56
r241 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.715 $Y=3.56
+ $X2=7.715 $Y2=3.56
r242 93 96 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=8.075 $Y=2.34
+ $X2=8.075 $Y2=3.56
r243 88 97 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=6.875 $Y=3.63
+ $X2=7.715 $Y2=3.63
r244 86 88 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=6.155 $Y=3.63
+ $X2=6.875 $Y2=3.63
r245 85 90 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=6.515 $Y=3.56
+ $X2=6.515 $Y2=3.59
r246 85 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.875 $Y=3.56
+ $X2=6.875 $Y2=3.56
r247 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.155 $Y=3.56
+ $X2=6.155 $Y2=3.56
r248 82 85 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=6.515 $Y=2.34
+ $X2=6.515 $Y2=3.56
r249 77 86 0.341676 $w=3.7e-07 $l=8.9e-07 $layer=MET1_cond $X=5.265 $Y=3.63
+ $X2=6.155 $Y2=3.63
r250 75 77 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=4.545 $Y=3.63
+ $X2=5.265 $Y2=3.63
r251 74 79 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=4.905 $Y=3.56
+ $X2=4.905 $Y2=3.57
r252 74 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.265 $Y=3.56
+ $X2=5.265 $Y2=3.56
r253 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.545 $Y=3.56
+ $X2=4.545 $Y2=3.56
r254 71 74 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=4.905 $Y=2.55
+ $X2=4.905 $Y2=3.56
r255 66 75 0.330159 $w=3.7e-07 $l=8.6e-07 $layer=MET1_cond $X=3.685 $Y=3.63
+ $X2=4.545 $Y2=3.63
r256 64 66 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.965 $Y=3.63
+ $X2=3.685 $Y2=3.63
r257 63 68 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=3.325 $Y=3.56
+ $X2=3.325 $Y2=3.57
r258 63 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.685 $Y=3.56
+ $X2=3.685 $Y2=3.56
r259 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.965 $Y=3.56
+ $X2=2.965 $Y2=3.56
r260 60 63 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=3.325 $Y=2.55
+ $X2=3.325 $Y2=3.56
r261 55 64 0.314802 $w=3.7e-07 $l=8.2e-07 $layer=MET1_cond $X=2.145 $Y=3.63
+ $X2=2.965 $Y2=3.63
r262 53 55 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.425 $Y=3.63
+ $X2=2.145 $Y2=3.63
r263 52 57 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=1.785 $Y=3.56
+ $X2=1.785 $Y2=3.57
r264 52 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.145 $Y=3.56
+ $X2=2.145 $Y2=3.56
r265 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.425 $Y=3.56
+ $X2=1.425 $Y2=3.56
r266 49 52 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=1.785 $Y=2.55
+ $X2=1.785 $Y2=3.56
r267 44 53 0.318641 $w=3.7e-07 $l=8.3e-07 $layer=MET1_cond $X=0.595 $Y=3.63
+ $X2=1.425 $Y2=3.63
r268 43 46 0.209838 $w=5.68e-07 $l=1e-08 $layer=LI1_cond $X=0.395 $Y=3.56
+ $X2=0.395 $Y2=3.57
r269 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.595 $Y=3.56
+ $X2=0.595 $Y2=3.56
r270 40 43 25.1806 $w=5.68e-07 $l=1.2e-06 $layer=LI1_cond $X=0.395 $Y=2.36
+ $X2=0.395 $Y2=3.56
r271 37 108 0.151643 $w=3.7e-07 $l=3.95e-07 $layer=MET1_cond $X=8.88 $Y=3.63
+ $X2=9.275 $Y2=3.63
r272 37 99 0.170838 $w=3.7e-07 $l=4.45e-07 $layer=MET1_cond $X=8.88 $Y=3.63
+ $X2=8.435 $Y2=3.63
r273 12 162 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=17.295
+ $Y=2.215 $X2=17.435 $Y2=3.57
r274 12 159 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=17.295
+ $Y=2.215 $X2=17.435 $Y2=2.36
r275 11 156 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=15.735
+ $Y=2.215 $X2=15.875 $Y2=3.59
r276 11 148 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=15.735
+ $Y=2.215 $X2=15.875 $Y2=2.34
r277 10 145 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=14.175
+ $Y=2.215 $X2=14.315 $Y2=3.59
r278 10 137 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=14.175
+ $Y=2.215 $X2=14.315 $Y2=2.34
r279 9 134 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=12.615
+ $Y=2.215 $X2=12.755 $Y2=3.59
r280 9 126 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=12.615
+ $Y=2.215 $X2=12.755 $Y2=2.34
r281 8 123 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=11.055
+ $Y=2.215 $X2=11.195 $Y2=3.59
r282 8 115 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=11.055
+ $Y=2.215 $X2=11.195 $Y2=2.34
r283 7 112 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=9.495
+ $Y=2.215 $X2=9.635 $Y2=3.59
r284 7 104 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=9.495
+ $Y=2.215 $X2=9.635 $Y2=2.34
r285 6 101 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=7.935
+ $Y=2.215 $X2=8.075 $Y2=3.59
r286 6 93 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=7.935
+ $Y=2.215 $X2=8.075 $Y2=2.34
r287 5 90 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=6.375
+ $Y=2.215 $X2=6.515 $Y2=3.59
r288 5 82 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=6.375
+ $Y=2.215 $X2=6.515 $Y2=2.34
r289 4 79 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=2.215 $X2=4.955 $Y2=3.57
r290 4 71 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=2.215 $X2=4.955 $Y2=2.55
r291 3 68 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=3.255
+ $Y=2.215 $X2=3.395 $Y2=3.57
r292 3 60 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=3.255
+ $Y=2.215 $X2=3.395 $Y2=2.55
r293 2 57 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=2.215 $X2=1.835 $Y2=3.57
r294 2 49 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=2.215 $X2=1.835 $Y2=2.55
r295 1 46 300 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.215 $X2=0.275 $Y2=3.57
r296 1 40 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.215 $X2=0.275 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 49
+ 66 76 86 96 106 116 126 136 145 146 148 149 151 152 154 155 158 159 160 162
+ 163 165 166
r208 154 158 0.539214 $w=1.7e-07 $l=5.6e-07 $layer=MET1_cond $X=11.83 $Y=2.405
+ $X2=11.27 $Y2=2.405
r209 139 143 35.1355 $w=4.08e-07 $l=1.25e-06 $layer=LI1_cond $X=16.695 $Y=2.34
+ $X2=16.695 $Y2=3.59
r210 136 139 38.9301 $w=4.08e-07 $l=1.385e-06 $layer=LI1_cond $X=16.695 $Y=0.955
+ $X2=16.695 $Y2=2.34
r211 129 133 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=15.095 $Y=2.34
+ $X2=15.095 $Y2=3.59
r212 126 129 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=15.095 $Y=0.955
+ $X2=15.095 $Y2=2.34
r213 119 123 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=13.535 $Y=2.34
+ $X2=13.535 $Y2=3.59
r214 116 119 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=13.535 $Y=0.955
+ $X2=13.535 $Y2=2.34
r215 109 113 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=11.975 $Y=2.34
+ $X2=11.975 $Y2=3.59
r216 106 109 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=11.975 $Y=0.955
+ $X2=11.975 $Y2=2.34
r217 99 103 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=10.415 $Y=2.34
+ $X2=10.415 $Y2=3.59
r218 96 99 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=10.415 $Y=0.955
+ $X2=10.415 $Y2=2.34
r219 89 93 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=8.855 $Y=2.34
+ $X2=8.855 $Y2=3.59
r220 86 89 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=8.855 $Y=0.955
+ $X2=8.855 $Y2=2.34
r221 79 83 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=7.295 $Y=2.34
+ $X2=7.295 $Y2=3.59
r222 76 79 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=7.295 $Y=0.955
+ $X2=7.295 $Y2=2.34
r223 69 73 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=5.735 $Y=2.34
+ $X2=5.735 $Y2=3.59
r224 66 69 48.3677 $w=3.28e-07 $l=1.385e-06 $layer=LI1_cond $X=5.735 $Y=0.955
+ $X2=5.735 $Y2=2.34
r225 49 165 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=16.655 $Y=2.405
+ $X2=16.51 $Y2=2.405
r226 49 166 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.095 $Y=2.405
+ $X2=15.24 $Y2=2.405
r227 49 162 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.095 $Y=2.405
+ $X2=14.95 $Y2=2.405
r228 49 163 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.535 $Y=2.405
+ $X2=13.68 $Y2=2.405
r229 49 159 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.535 $Y=2.405
+ $X2=13.39 $Y2=2.405
r230 49 160 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.975 $Y=2.405
+ $X2=12.12 $Y2=2.405
r231 49 154 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.975 $Y=2.405
+ $X2=11.83 $Y2=2.405
r232 49 155 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.415 $Y=2.405
+ $X2=10.56 $Y2=2.405
r233 49 151 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.415 $Y=2.405
+ $X2=10.27 $Y2=2.405
r234 49 152 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.855 $Y=2.405
+ $X2=9 $Y2=2.405
r235 49 148 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.855 $Y=2.405
+ $X2=8.71 $Y2=2.405
r236 49 149 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.295 $Y=2.405
+ $X2=7.44 $Y2=2.405
r237 49 145 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.295 $Y=2.405
+ $X2=7.15 $Y2=2.405
r238 49 146 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.735 $Y=2.405
+ $X2=5.88 $Y2=2.405
r239 49 165 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=15.875 $Y=2.405
+ $X2=16.51 $Y2=2.405
r240 49 166 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=15.875 $Y=2.405
+ $X2=15.24 $Y2=2.405
r241 49 162 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=14.315 $Y=2.405
+ $X2=14.95 $Y2=2.405
r242 49 163 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=14.315 $Y=2.405
+ $X2=13.68 $Y2=2.405
r243 49 159 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=12.755 $Y=2.405
+ $X2=13.39 $Y2=2.405
r244 49 160 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=12.755 $Y=2.405
+ $X2=12.12 $Y2=2.405
r245 49 158 0.0722162 $w=1.7e-07 $l=7.5e-08 $layer=MET1_cond $X=11.195 $Y=2.405
+ $X2=11.27 $Y2=2.405
r246 49 155 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=11.195 $Y=2.405
+ $X2=10.56 $Y2=2.405
r247 49 151 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=9.635 $Y=2.405
+ $X2=10.27 $Y2=2.405
r248 49 152 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=9.635 $Y=2.405
+ $X2=9 $Y2=2.405
r249 49 148 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=8.075 $Y=2.405
+ $X2=8.71 $Y2=2.405
r250 49 149 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=8.075 $Y=2.405
+ $X2=7.44 $Y2=2.405
r251 49 145 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=6.515 $Y=2.405
+ $X2=7.15 $Y2=2.405
r252 49 146 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=6.515 $Y=2.405
+ $X2=5.88 $Y2=2.405
r253 49 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.655 $Y=2.405
+ $X2=16.655 $Y2=2.405
r254 49 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.095 $Y=2.405
+ $X2=15.095 $Y2=2.405
r255 49 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.535 $Y=2.405
+ $X2=13.535 $Y2=2.405
r256 49 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.975 $Y=2.405
+ $X2=11.975 $Y2=2.405
r257 49 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.415 $Y=2.405
+ $X2=10.415 $Y2=2.405
r258 49 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.855 $Y=2.405
+ $X2=8.855 $Y2=2.405
r259 49 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.295 $Y=2.405
+ $X2=7.295 $Y2=2.405
r260 49 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.735 $Y=2.405
+ $X2=5.735 $Y2=2.405
r261 16 143 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=16.515
+ $Y=2.215 $X2=16.655 $Y2=3.59
r262 16 139 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=16.515
+ $Y=2.215 $X2=16.655 $Y2=2.34
r263 15 133 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=14.955
+ $Y=2.215 $X2=15.095 $Y2=3.59
r264 15 129 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=14.955
+ $Y=2.215 $X2=15.095 $Y2=2.34
r265 14 123 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=13.395
+ $Y=2.215 $X2=13.535 $Y2=3.59
r266 14 119 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=13.395
+ $Y=2.215 $X2=13.535 $Y2=2.34
r267 13 113 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=11.835
+ $Y=2.215 $X2=11.975 $Y2=3.59
r268 13 109 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=11.835
+ $Y=2.215 $X2=11.975 $Y2=2.34
r269 12 103 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=10.275
+ $Y=2.215 $X2=10.415 $Y2=3.59
r270 12 99 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=10.275
+ $Y=2.215 $X2=10.415 $Y2=2.34
r271 11 93 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=8.715
+ $Y=2.215 $X2=8.855 $Y2=3.59
r272 11 89 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=8.715
+ $Y=2.215 $X2=8.855 $Y2=2.34
r273 10 83 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=7.155
+ $Y=2.215 $X2=7.295 $Y2=3.59
r274 10 79 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=7.155
+ $Y=2.215 $X2=7.295 $Y2=2.34
r275 9 73 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=5.595
+ $Y=2.215 $X2=5.735 $Y2=3.59
r276 9 69 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=5.595
+ $Y=2.215 $X2=5.735 $Y2=2.34
r277 8 136 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=16.515
+ $Y=0.705 $X2=16.655 $Y2=0.955
r278 7 126 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=14.955
+ $Y=0.705 $X2=15.095 $Y2=0.955
r279 6 116 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=13.395
+ $Y=0.705 $X2=13.535 $Y2=0.955
r280 5 106 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=11.835
+ $Y=0.705 $X2=11.975 $Y2=0.955
r281 4 96 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=10.275
+ $Y=0.705 $X2=10.415 $Y2=0.955
r282 3 86 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=8.715
+ $Y=0.705 $X2=8.855 $Y2=0.955
r283 2 76 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=7.155
+ $Y=0.705 $X2=7.295 $Y2=0.955
r284 1 66 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=5.595
+ $Y=0.705 $X2=5.735 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 37 40 47 56
+ 65 74 83 92 101 110 119 128 137 138
r171 137 141 10.0425 $w=5.28e-07 $l=4.45e-07 $layer=LI1_cond $X=17.335 $Y=0.51
+ $X2=17.335 $Y2=0.955
r172 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.515 $Y=0.51
+ $X2=17.515 $Y2=0.51
r173 132 138 0.491399 $w=3.7e-07 $l=1.28e-06 $layer=MET1_cond $X=16.235 $Y=0.44
+ $X2=17.515 $Y2=0.44
r174 129 132 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=15.515 $Y=0.44
+ $X2=16.235 $Y2=0.44
r175 128 134 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=15.875 $Y=0.51
+ $X2=15.875 $Y2=0.92
r176 128 132 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.235 $Y=0.51
+ $X2=16.235 $Y2=0.51
r177 128 129 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.515 $Y=0.51
+ $X2=15.515 $Y2=0.51
r178 123 129 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=14.675 $Y=0.44
+ $X2=15.515 $Y2=0.44
r179 120 123 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=13.955 $Y=0.44
+ $X2=14.675 $Y2=0.44
r180 119 125 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=14.315 $Y=0.51
+ $X2=14.315 $Y2=0.92
r181 119 123 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.675 $Y=0.51
+ $X2=14.675 $Y2=0.51
r182 119 120 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.955 $Y=0.51
+ $X2=13.955 $Y2=0.51
r183 114 120 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=13.115 $Y=0.44
+ $X2=13.955 $Y2=0.44
r184 111 114 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=12.395 $Y=0.44
+ $X2=13.115 $Y2=0.44
r185 110 116 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=12.755 $Y=0.51
+ $X2=12.755 $Y2=0.92
r186 110 114 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.115 $Y=0.51
+ $X2=13.115 $Y2=0.51
r187 110 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.395 $Y=0.51
+ $X2=12.395 $Y2=0.51
r188 105 111 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=11.555 $Y=0.44
+ $X2=12.395 $Y2=0.44
r189 102 105 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.835 $Y=0.44
+ $X2=11.555 $Y2=0.44
r190 101 107 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=11.195 $Y=0.51
+ $X2=11.195 $Y2=0.92
r191 101 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.555 $Y=0.51
+ $X2=11.555 $Y2=0.51
r192 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.835 $Y=0.51
+ $X2=10.835 $Y2=0.51
r193 96 102 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=9.995 $Y=0.44
+ $X2=10.835 $Y2=0.44
r194 93 96 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=9.275 $Y=0.44
+ $X2=9.995 $Y2=0.44
r195 92 98 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=9.635 $Y=0.51
+ $X2=9.635 $Y2=0.92
r196 92 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.995 $Y=0.51
+ $X2=9.995 $Y2=0.51
r197 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.275 $Y=0.51
+ $X2=9.275 $Y2=0.51
r198 84 87 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.715 $Y=0.44
+ $X2=8.435 $Y2=0.44
r199 83 89 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=8.075 $Y=0.51
+ $X2=8.075 $Y2=0.92
r200 83 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.435 $Y=0.51
+ $X2=8.435 $Y2=0.51
r201 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.715 $Y=0.51
+ $X2=7.715 $Y2=0.51
r202 78 84 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=6.875 $Y=0.44
+ $X2=7.715 $Y2=0.44
r203 75 78 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=6.155 $Y=0.44
+ $X2=6.875 $Y2=0.44
r204 74 80 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=6.515 $Y=0.51
+ $X2=6.515 $Y2=0.92
r205 74 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.875 $Y=0.51
+ $X2=6.875 $Y2=0.51
r206 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.155 $Y=0.51
+ $X2=6.155 $Y2=0.51
r207 69 75 0.349354 $w=3.7e-07 $l=9.1e-07 $layer=MET1_cond $X=5.245 $Y=0.44
+ $X2=6.155 $Y2=0.44
r208 66 69 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=4.525 $Y=0.44
+ $X2=5.245 $Y2=0.44
r209 65 71 5.62022 $w=8.88e-07 $l=4.1e-07 $layer=LI1_cond $X=4.885 $Y=0.51
+ $X2=4.885 $Y2=0.92
r210 65 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.245 $Y=0.51
+ $X2=5.245 $Y2=0.51
r211 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.525 $Y=0.51
+ $X2=4.525 $Y2=0.51
r212 60 66 0.291768 $w=3.7e-07 $l=7.6e-07 $layer=MET1_cond $X=3.765 $Y=0.44
+ $X2=4.525 $Y2=0.44
r213 57 60 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.045 $Y=0.44
+ $X2=3.765 $Y2=0.44
r214 56 62 5.86145 $w=8.93e-07 $l=4.3e-07 $layer=LI1_cond $X=3.407 $Y=0.51
+ $X2=3.407 $Y2=0.94
r215 56 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.765 $Y=0.51
+ $X2=3.765 $Y2=0.51
r216 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.045 $Y=0.51
+ $X2=3.045 $Y2=0.51
r217 51 57 0.345515 $w=3.7e-07 $l=9e-07 $layer=MET1_cond $X=2.145 $Y=0.44
+ $X2=3.045 $Y2=0.44
r218 48 51 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.425 $Y=0.44
+ $X2=2.145 $Y2=0.44
r219 47 53 5.89438 $w=8.88e-07 $l=4.3e-07 $layer=LI1_cond $X=1.785 $Y=0.51
+ $X2=1.785 $Y2=0.94
r220 47 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.145 $Y=0.51
+ $X2=2.145 $Y2=0.51
r221 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.425 $Y=0.51
+ $X2=1.425 $Y2=0.51
r222 41 48 0.332078 $w=3.7e-07 $l=8.65e-07 $layer=MET1_cond $X=0.56 $Y=0.44
+ $X2=1.425 $Y2=0.44
r223 40 44 9.61334 $w=5.33e-07 $l=4.3e-07 $layer=LI1_cond $X=0.377 $Y=0.51
+ $X2=0.377 $Y2=0.94
r224 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.56 $Y=0.51
+ $X2=0.56 $Y2=0.51
r225 37 93 0.151643 $w=3.7e-07 $l=3.95e-07 $layer=MET1_cond $X=8.88 $Y=0.44
+ $X2=9.275 $Y2=0.44
r226 37 87 0.170838 $w=3.7e-07 $l=4.45e-07 $layer=MET1_cond $X=8.88 $Y=0.44
+ $X2=8.435 $Y2=0.44
r227 12 141 91 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=2 $X=17.295
+ $Y=0.705 $X2=17.435 $Y2=0.955
r228 11 134 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=15.735
+ $Y=0.705 $X2=15.875 $Y2=0.92
r229 10 125 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=14.175
+ $Y=0.705 $X2=14.315 $Y2=0.92
r230 9 116 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=12.615
+ $Y=0.705 $X2=12.755 $Y2=0.92
r231 8 107 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=11.055
+ $Y=0.705 $X2=11.195 $Y2=0.92
r232 7 98 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=9.495
+ $Y=0.705 $X2=9.635 $Y2=0.92
r233 6 89 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=7.935
+ $Y=0.705 $X2=8.075 $Y2=0.92
r234 5 80 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=6.375
+ $Y=0.705 $X2=6.515 $Y2=0.92
r235 4 71 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=4.815
+ $Y=0.705 $X2=4.955 $Y2=0.92
r236 3 62 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.255
+ $Y=0.705 $X2=3.395 $Y2=0.94
r237 2 53 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.705 $X2=1.835 $Y2=0.94
r238 1 44 91 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.705 $X2=0.275 $Y2=0.94
.ends

