* NGSPICE file created from sky130_fd_sc_hvl__mux2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__mux2_1 A0 A1 S VGND VNB VPB VPWR X
M1000 a_671_491# A1 a_94_81# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1001 a_373_107# S VGND VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=3.7755e+11p ps=3.69e+06u
M1002 VPWR a_94_81# X VPB phv w=1.5e+06u l=500000u
+  ad=5.913e+11p pd=5.19e+06u as=4.275e+11p ps=3.57e+06u
M1003 VGND a_713_81# a_671_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1004 a_373_491# S VPWR VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1005 VPWR a_713_81# a_671_491# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_94_81# A1 a_373_107# VNB nhv w=420000u l=500000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1007 a_94_81# A0 a_373_491# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_713_81# S VGND VNB nhv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1009 VGND a_94_81# X VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=2.1375e+11p ps=2.07e+06u
M1010 a_713_81# S VPWR VPB phv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1011 a_671_107# A0 a_94_81# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends

