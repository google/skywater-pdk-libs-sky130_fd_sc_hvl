* File: sky130_fd_sc_hvl__sdlxtp_1.pex.spice
* Created: Wed Sep  2 09:10:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%VNB 5 7 11 25
r92 7 25 1.08507e-05 $w=1.152e-05 $l=1e-09 $layer=MET1_cond $X=5.76 $Y=0.057
+ $X2=5.76 $Y2=0.058
r93 7 11 0.00061849 $w=1.152e-05 $l=5.7e-08 $layer=MET1_cond $X=5.76 $Y=0.057
+ $X2=5.76 $Y2=0
r94 5 11 0.775 $w=1.7e-07 $l=2.04e-06 $layer=mcon $count=12 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r95 5 11 0.775 $w=1.7e-07 $l=2.04e-06 $layer=mcon $count=12 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%VPB 4 6 14 21
r114 10 21 0.00061849 $w=1.152e-05 $l=5.7e-08 $layer=MET1_cond $X=5.76 $Y=4.07
+ $X2=5.76 $Y2=4.013
r115 10 14 0.775 $w=1.7e-07 $l=2.04e-06 $layer=mcon $count=12 $X=11.28 $Y=4.07
+ $X2=11.28 $Y2=4.07
r116 9 14 720.257 $w=1.68e-07 $l=1.104e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=11.28 $Y2=4.07
r117 9 10 0.775 $w=1.7e-07 $l=2.04e-06 $layer=mcon $count=12 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r118 6 21 1.08507e-05 $w=1.152e-05 $l=1e-09 $layer=MET1_cond $X=5.76 $Y=4.012
+ $X2=5.76 $Y2=4.013
r119 4 14 15.1667 $w=1.7e-07 $l=1.13224e-05 $layer=licon1_NTAP_notbjt $count=12
+ $X=0 $Y=3.985 $X2=11.28 $Y2=4.07
r120 4 9 15.1667 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=12
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%SCE 3 6 8 10 13 17 18 21 25 26 28 29 30 34
+ 36 43 58
c78 26 0 3.90348e-19 $X=2.82 $Y=1.53
r79 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.34
+ $Y=2.61 $X2=1.34 $Y2=2.61
r80 40 43 73.8649 $w=3.85e-07 $l=5.9e-07 $layer=POLY_cond $X=0.75 $Y=2.625
+ $X2=1.34 $Y2=2.625
r81 37 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=2.61 $X2=0.75 $Y2=2.61
r82 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=2.27 $X2=0.75 $Y2=2.27
r83 34 40 8.13766 $w=3.85e-07 $l=6.5e-08 $layer=POLY_cond $X=0.685 $Y=2.625
+ $X2=0.75 $Y2=2.625
r84 34 36 16.5859 $w=5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.685 $Y=2.425
+ $X2=0.685 $Y2=2.27
r85 30 58 11.859 $w=9.38e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=2.305
+ $X2=1.795 $Y2=2.305
r86 30 44 4.41277 $w=9.38e-07 $l=3.4e-07 $layer=LI1_cond $X=1.68 $Y=2.305
+ $X2=1.34 $Y2=2.305
r87 29 44 1.81702 $w=9.38e-07 $l=1.4e-07 $layer=LI1_cond $X=1.2 $Y=2.305
+ $X2=1.34 $Y2=2.305
r88 29 37 5.84043 $w=9.38e-07 $l=4.5e-07 $layer=LI1_cond $X=1.2 $Y=2.305
+ $X2=0.75 $Y2=2.305
r89 28 37 0.389362 $w=9.38e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=2.305
+ $X2=0.75 $Y2=2.305
r90 26 47 42.7144 $w=5.7e-07 $l=4.45e-07 $layer=POLY_cond $X=2.94 $Y=1.53
+ $X2=2.94 $Y2=1.085
r91 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.82
+ $Y=1.53 $X2=2.82 $Y2=1.53
r92 22 25 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=2.685 $Y=1.57
+ $X2=2.82 $Y2=1.57
r93 20 22 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.685 $Y=1.695
+ $X2=2.685 $Y2=1.57
r94 20 21 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.685 $Y=1.695
+ $X2=2.685 $Y2=1.835
r95 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.6 $Y=1.92
+ $X2=2.685 $Y2=1.835
r96 18 58 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=2.6 $Y=1.92
+ $X2=1.795 $Y2=1.92
r97 17 36 73.299 $w=5e-07 $l=6.85e-07 $layer=POLY_cond $X=0.685 $Y=1.585
+ $X2=0.685 $Y2=2.27
r98 16 17 51.4451 $w=5.2e-07 $l=5e-07 $layer=POLY_cond $X=0.695 $Y=1.085
+ $X2=0.695 $Y2=1.585
r99 13 47 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.975 $Y=0.745
+ $X2=2.975 $Y2=1.085
r100 8 43 27.5429 $w=3.85e-07 $l=2.2e-07 $layer=POLY_cond $X=1.56 $Y=2.625
+ $X2=1.34 $Y2=2.625
r101 8 10 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.56 $Y=2.825 $X2=1.56
+ $Y2=3.31
r102 6 16 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.705 $Y=0.745
+ $X2=0.705 $Y2=1.085
r103 3 34 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.685 $Y=3.145
+ $X2=0.685 $Y2=2.825
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%A_30_587# 1 2 9 13 15 17 23 24 32 33 34 36
+ 43
r84 33 43 132.687 $w=5e-07 $l=1.24e-06 $layer=POLY_cond $X=3.05 $Y=2.07 $X2=3.05
+ $Y2=3.31
r85 32 34 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=3.142 $Y=2.07
+ $X2=3.142 $Y2=1.905
r86 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.115
+ $Y=2.07 $X2=3.115 $Y2=2.07
r87 28 36 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.195 $Y=1.23
+ $X2=2.195 $Y2=0.745
r88 27 29 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=2.13 $Y=1.23 $X2=2.13
+ $Y2=1.26
r89 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.13
+ $Y=1.23 $X2=2.13 $Y2=1.23
r90 24 27 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=2.13 $Y=1.18 $X2=2.13
+ $Y2=1.23
r91 21 34 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.25 $Y=1.265
+ $X2=3.25 $Y2=1.905
r92 18 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=1.18
+ $X2=2.13 $Y2=1.18
r93 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.165 $Y=1.18
+ $X2=3.25 $Y2=1.265
r94 17 18 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.165 $Y=1.18
+ $X2=2.295 $Y2=1.18
r95 16 23 3.44808 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.48 $Y=1.26
+ $X2=0.305 $Y2=1.26
r96 15 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=1.26
+ $X2=2.13 $Y2=1.26
r97 15 16 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=1.965 $Y=1.26
+ $X2=0.48 $Y2=1.26
r98 11 23 3.14896 $w=3e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.255 $Y=1.345
+ $X2=0.305 $Y2=1.26
r99 11 13 82.9759 $w=2.48e-07 $l=1.8e-06 $layer=LI1_cond $X=0.255 $Y=1.345
+ $X2=0.255 $Y2=3.145
r100 7 23 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.305 $Y=1.175
+ $X2=0.305 $Y2=1.26
r101 7 9 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.305 $Y=1.175
+ $X2=0.305 $Y2=0.745
r102 2 13 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.935 $X2=0.295 $Y2=3.145
r103 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.535 $X2=0.315 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%D 3 7 9 10 11 17 18
r41 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.205
+ $Y=2.27 $X2=2.205 $Y2=2.27
r42 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.205 $Y=2.775
+ $X2=2.205 $Y2=3.145
r43 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.205 $Y=2.405
+ $X2=2.205 $Y2=2.775
r44 9 18 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.205 $Y=2.405
+ $X2=2.205 $Y2=2.27
r45 7 17 109.681 $w=5e-07 $l=1.025e-06 $layer=POLY_cond $X=2.27 $Y=3.31 $X2=2.27
+ $Y2=2.285
r46 1 17 114.914 $w=3.02e-07 $l=7.2e-07 $layer=POLY_cond $X=1.485 $Y=2.12
+ $X2=2.205 $Y2=2.12
r47 1 3 129.477 $w=5e-07 $l=1.21e-06 $layer=POLY_cond $X=1.485 $Y=1.955
+ $X2=1.485 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%SCD 3 7 8 9 10 15 21
c41 8 0 1.6729e-19 $X=3.6 $Y=1.665
r42 18 21 100.586 $w=5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.76 $Y=2.37 $X2=3.76
+ $Y2=3.31
r43 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.695
+ $Y=2.37 $X2=3.695 $Y2=2.37
r44 15 18 72.764 $w=5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.76 $Y=1.69 $X2=3.76
+ $Y2=2.37
r45 15 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.695
+ $Y=1.69 $X2=3.695 $Y2=1.69
r46 10 19 1.16915 $w=3.43e-07 $l=3.5e-08 $layer=LI1_cond $X=3.687 $Y=2.405
+ $X2=3.687 $Y2=2.37
r47 9 19 11.1904 $w=3.43e-07 $l=3.35e-07 $layer=LI1_cond $X=3.687 $Y=2.035
+ $X2=3.687 $Y2=2.37
r48 9 16 11.5244 $w=3.43e-07 $l=3.45e-07 $layer=LI1_cond $X=3.687 $Y=2.035
+ $X2=3.687 $Y2=1.69
r49 8 16 0.835104 $w=3.43e-07 $l=2.5e-08 $layer=LI1_cond $X=3.687 $Y=1.665
+ $X2=3.687 $Y2=1.69
r50 7 15 11.2356 $w=5e-07 $l=1.05e-07 $layer=POLY_cond $X=3.76 $Y=1.585 $X2=3.76
+ $Y2=1.69
r51 6 7 46.5243 $w=5.75e-07 $l=5e-07 $layer=POLY_cond $X=3.722 $Y=1.085
+ $X2=3.722 $Y2=1.585
r52 3 6 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.685 $Y=0.745 $X2=3.685
+ $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%GATE 3 7 9 10 11 12 13 20 23
r40 23 25 22.0641 $w=5.7e-07 $l=2.25e-07 $layer=POLY_cond $X=4.505 $Y=1.31
+ $X2=4.505 $Y2=1.085
r41 18 23 5.63189 $w=5.7e-07 $l=6e-08 $layer=POLY_cond $X=4.505 $Y=1.37
+ $X2=4.505 $Y2=1.31
r42 18 20 90.1102 $w=5.7e-07 $l=9.6e-07 $layer=POLY_cond $X=4.505 $Y=1.37
+ $X2=4.505 $Y2=2.33
r43 13 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.52
+ $Y=2.33 $X2=4.52 $Y2=2.33
r44 12 13 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=4.517 $Y=2.035
+ $X2=4.517 $Y2=2.33
r45 11 12 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=4.517 $Y=1.665
+ $X2=4.517 $Y2=2.035
r46 10 11 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=4.517 $Y=1.295
+ $X2=4.517 $Y2=1.665
r47 10 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.52
+ $Y=1.31 $X2=4.52 $Y2=1.31
r48 8 20 19.7116 $w=5.7e-07 $l=2.1e-07 $layer=POLY_cond $X=4.505 $Y=2.54
+ $X2=4.505 $Y2=2.33
r49 8 9 27.696 $w=5.7e-07 $l=2.85e-07 $layer=POLY_cond $X=4.505 $Y=2.54
+ $X2=4.505 $Y2=2.825
r50 7 9 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.54 $Y=3.31 $X2=4.54
+ $Y2=2.825
r51 3 25 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.47 $Y=0.745 $X2=4.47
+ $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%A_1214_107# 1 2 7 9 14 19 21 22 26 28 29
+ 31 32 34 37 38 40
r91 37 38 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=6.33 $Y=0.975
+ $X2=6.33 $Y2=2.585
r92 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.405
+ $Y=2.38 $X2=8.405 $Y2=2.38
r93 32 34 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=8.01 $Y=2.345
+ $X2=8.405 $Y2=2.345
r94 31 32 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.925 $Y=2.215
+ $X2=8.01 $Y2=2.345
r95 30 31 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.925 $Y=1.755
+ $X2=7.925 $Y2=2.215
r96 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.84 $Y=1.67
+ $X2=7.925 $Y2=1.755
r97 28 29 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=7.84 $Y=1.67
+ $X2=7.275 $Y2=1.67
r98 27 40 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.15 $Y=1.25 $X2=7.15
+ $Y2=0.745
r99 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.19
+ $Y=1.25 $X2=7.19 $Y2=1.25
r100 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.19 $Y=1.585
+ $X2=7.275 $Y2=1.67
r101 24 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.19 $Y=1.585
+ $X2=7.19 $Y2=1.25
r102 23 26 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=7.19 $Y=0.435
+ $X2=7.19 $Y2=1.25
r103 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.105 $Y=0.35
+ $X2=7.19 $Y2=0.435
r104 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.105 $Y=0.35
+ $X2=6.415 $Y2=0.35
r105 19 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.41 $Y=2.75
+ $X2=6.41 $Y2=2.585
r106 12 37 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.23 $Y=0.79
+ $X2=6.23 $Y2=0.975
r107 12 14 1.40162 $w=3.68e-07 $l=4.5e-08 $layer=LI1_cond $X=6.23 $Y=0.79
+ $X2=6.23 $Y2=0.745
r108 11 22 8.10976 $w=1.7e-07 $l=2.23495e-07 $layer=LI1_cond $X=6.23 $Y=0.435
+ $X2=6.415 $Y2=0.35
r109 11 14 9.6556 $w=3.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.23 $Y=0.435
+ $X2=6.23 $Y2=0.745
r110 7 35 38.8218 $w=5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.37 $Y=2.775
+ $X2=8.37 $Y2=2.38
r111 7 9 42.8024 $w=5e-07 $l=4e-07 $layer=POLY_cond $X=8.37 $Y=2.775 $X2=8.37
+ $Y2=3.175
r112 2 19 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=6.27
+ $Y=2.625 $X2=6.41 $Y2=2.75
r113 1 14 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.07
+ $Y=0.535 $X2=6.21 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%A_944_107# 1 2 7 9 10 12 14 18 21 24 27 29
+ 34 37 39 42
r111 40 42 63.6685 $w=5e-07 $l=5.95e-07 $layer=POLY_cond $X=5.82 $Y=1.34
+ $X2=5.82 $Y2=0.745
r112 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.755
+ $Y=1.34 $X2=5.755 $Y2=1.34
r113 34 36 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.86 $Y=0.745
+ $X2=4.86 $Y2=0.975
r114 30 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.015 $Y=1.26
+ $X2=4.93 $Y2=1.26
r115 29 39 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=1.26
+ $X2=5.755 $Y2=1.26
r116 29 30 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=5.59 $Y=1.26
+ $X2=5.015 $Y2=1.26
r117 25 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=1.345
+ $X2=4.93 $Y2=1.26
r118 25 27 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=4.93 $Y=1.345
+ $X2=4.93 $Y2=3.175
r119 24 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=1.175
+ $X2=4.93 $Y2=1.26
r120 24 36 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.93 $Y=1.175
+ $X2=4.93 $Y2=0.975
r121 20 40 72.229 $w=5e-07 $l=6.75e-07 $layer=POLY_cond $X=5.82 $Y=2.015
+ $X2=5.82 $Y2=1.34
r122 20 21 20.4101 $w=5e-07 $l=2.95804e-07 $layer=POLY_cond $X=5.82 $Y=2.015
+ $X2=5.92 $Y2=2.265
r123 16 22 64.8397 $w=6.21e-07 $l=9.16941e-07 $layer=POLY_cond $X=7.93 $Y=1.455
+ $X2=7.702 $Y2=2.265
r124 16 18 75.9742 $w=5e-07 $l=7.1e-07 $layer=POLY_cond $X=7.93 $Y=1.455
+ $X2=7.93 $Y2=0.745
r125 12 22 21.3743 $w=6.21e-07 $l=3.45326e-07 $layer=POLY_cond $X=7.475 $Y=2.515
+ $X2=7.702 $Y2=2.265
r126 12 14 88.2799 $w=5e-07 $l=8.25e-07 $layer=POLY_cond $X=7.475 $Y=2.515
+ $X2=7.475 $Y2=3.34
r127 11 21 5.30422 $w=5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.27 $Y=2.265
+ $X2=5.92 $Y2=2.265
r128 10 22 7.93667 $w=5e-07 $l=4.77e-07 $layer=POLY_cond $X=7.225 $Y=2.265
+ $X2=7.702 $Y2=2.265
r129 10 11 102.191 $w=5e-07 $l=9.55e-07 $layer=POLY_cond $X=7.225 $Y=2.265
+ $X2=6.27 $Y2=2.265
r130 7 21 20.4101 $w=5e-07 $l=2.95804e-07 $layer=POLY_cond $X=6.02 $Y=2.515
+ $X2=5.92 $Y2=2.265
r131 7 9 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.02 $Y=2.515 $X2=6.02
+ $Y2=3
r132 2 27 600 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=1 $X=4.79
+ $Y=2.935 $X2=4.93 $Y2=3.175
r133 1 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.72
+ $Y=0.535 $X2=4.86 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%A_1678_81# 1 2 7 9 12 14 18 20 22 25 27 32
+ 37 41
c77 37 0 1.37987e-19 $X=9.58 $Y=1.49
c78 22 0 1.67544e-19 $X=10.38 $Y=1.49
r79 32 35 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=9.55 $Y=2.27
+ $X2=9.55 $Y2=2.425
r80 28 41 27.9441 $w=6.9e-07 $l=3.75e-07 $layer=POLY_cond $X=8.705 $Y=1.41
+ $X2=9.08 $Y2=1.41
r81 28 38 4.84365 $w=6.9e-07 $l=6.5e-08 $layer=POLY_cond $X=8.705 $Y=1.41
+ $X2=8.64 $Y2=1.41
r82 27 30 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=8.705 $Y=1.23
+ $X2=8.705 $Y2=1.49
r83 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.705
+ $Y=1.23 $X2=8.705 $Y2=1.23
r84 24 25 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=10.465 $Y=1.575
+ $X2=10.465 $Y2=2.185
r85 23 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.745 $Y=1.49
+ $X2=9.58 $Y2=1.49
r86 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.38 $Y=1.49
+ $X2=10.465 $Y2=1.575
r87 22 23 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.38 $Y=1.49
+ $X2=9.745 $Y2=1.49
r88 21 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.715 $Y=2.27
+ $X2=9.55 $Y2=2.27
r89 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.38 $Y=2.27
+ $X2=10.465 $Y2=2.185
r90 20 21 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=10.38 $Y=2.27
+ $X2=9.715 $Y2=2.27
r91 16 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.58 $Y=1.405
+ $X2=9.58 $Y2=1.49
r92 16 18 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=9.58 $Y=1.405
+ $X2=9.58 $Y2=1.075
r93 15 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.87 $Y=1.49
+ $X2=8.705 $Y2=1.49
r94 14 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.415 $Y=1.49
+ $X2=9.58 $Y2=1.49
r95 14 15 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=9.415 $Y=1.49
+ $X2=8.87 $Y2=1.49
r96 10 41 10.3696 $w=5e-07 $l=3.45e-07 $layer=POLY_cond $X=9.08 $Y=1.755
+ $X2=9.08 $Y2=1.41
r97 10 12 151.948 $w=5e-07 $l=1.42e-06 $layer=POLY_cond $X=9.08 $Y=1.755
+ $X2=9.08 $Y2=3.175
r98 7 38 10.3696 $w=5e-07 $l=3.45e-07 $layer=POLY_cond $X=8.64 $Y=1.065 $X2=8.64
+ $Y2=1.41
r99 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.64 $Y=1.065 $X2=8.64
+ $Y2=0.745
r100 2 35 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=9.405
+ $Y=2.215 $X2=9.55 $Y2=2.425
r101 1 18 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.455
+ $Y=0.865 $X2=9.58 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%A_1480_107# 1 2 9 13 17 21 25 29 31 33 34
+ 35 38 39 40 42 46 48 50 57
c123 21 0 1.67544e-19 $X=10.845 $Y=0.91
c124 13 0 1.37987e-19 $X=9.97 $Y=1.075
r125 56 57 0.798551 $w=6.7e-07 $l=1e-08 $layer=POLY_cond $X=10.835 $Y=1.75
+ $X2=10.845 $Y2=1.75
r126 52 54 2.39565 $w=6.7e-07 $l=3e-08 $layer=POLY_cond $X=9.94 $Y=1.75 $X2=9.97
+ $Y2=1.75
r127 49 56 63.8841 $w=6.7e-07 $l=8e-07 $layer=POLY_cond $X=10.035 $Y=1.75
+ $X2=10.835 $Y2=1.75
r128 49 54 5.19058 $w=6.7e-07 $l=6.5e-08 $layer=POLY_cond $X=10.035 $Y=1.75
+ $X2=9.97 $Y2=1.75
r129 48 50 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=10.035 $Y=1.88
+ $X2=9.87 $Y2=1.88
r130 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.035
+ $Y=1.88 $X2=10.035 $Y2=1.88
r131 44 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.92 $Y=1.92
+ $X2=8.835 $Y2=1.92
r132 44 50 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=8.92 $Y=1.92
+ $X2=9.87 $Y2=1.92
r133 41 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.835 $Y=2.005
+ $X2=8.835 $Y2=1.92
r134 41 42 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.835 $Y=2.005
+ $X2=8.835 $Y2=2.655
r135 39 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.75 $Y=1.92
+ $X2=8.835 $Y2=1.92
r136 39 40 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.75 $Y=1.92
+ $X2=8.36 $Y2=1.92
r137 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.275 $Y=1.835
+ $X2=8.36 $Y2=1.92
r138 37 38 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.275 $Y=1.245
+ $X2=8.275 $Y2=1.835
r139 36 45 2.50919 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.03 $Y=2.74
+ $X2=7.865 $Y2=2.74
r140 35 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.75 $Y=2.74
+ $X2=8.835 $Y2=2.655
r141 35 36 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=8.75 $Y=2.74
+ $X2=8.03 $Y2=2.74
r142 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.19 $Y=1.16
+ $X2=8.275 $Y2=1.245
r143 33 34 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=8.19 $Y=1.16
+ $X2=7.705 $Y2=1.16
r144 29 45 14.0725 $w=3.3e-07 $l=3.5e-07 $layer=LI1_cond $X=7.865 $Y=3.09
+ $X2=7.865 $Y2=2.74
r145 29 31 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=7.865 $Y=3.09
+ $X2=7.865 $Y2=3.59
r146 23 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.58 $Y=1.075
+ $X2=7.705 $Y2=1.16
r147 23 25 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=7.58 $Y=1.075
+ $X2=7.58 $Y2=0.745
r148 19 57 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.845 $Y=1.415
+ $X2=10.845 $Y2=1.75
r149 19 21 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=10.845 $Y=1.415
+ $X2=10.845 $Y2=0.91
r150 15 56 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.835 $Y=2.085
+ $X2=10.835 $Y2=1.75
r151 15 17 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=10.835 $Y=2.085
+ $X2=10.835 $Y2=2.965
r152 11 54 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.97 $Y=1.415
+ $X2=9.97 $Y2=1.75
r153 11 13 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=9.97 $Y=1.415 $X2=9.97
+ $Y2=1.075
r154 7 52 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.94 $Y=2.085
+ $X2=9.94 $Y2=1.75
r155 7 9 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=9.94 $Y=2.085 $X2=9.94
+ $Y2=2.425
r156 2 31 600 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=1 $X=7.725
+ $Y=2.965 $X2=7.865 $Y2=3.59
r157 2 29 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=7.725
+ $Y=2.965 $X2=7.865 $Y2=3.09
r158 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.4
+ $Y=0.535 $X2=7.54 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%VPWR 1 2 3 4 5 16 19 36 40 47 56 63
r90 60 63 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.01 $Y=3.63
+ $X2=10.73 $Y2=3.63
r91 59 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.73 $Y=3.59
+ $X2=10.73 $Y2=3.59
r92 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.01 $Y=3.59
+ $X2=10.01 $Y2=3.59
r93 56 59 12.4568 $w=9.48e-07 $l=9.7e-07 $layer=LI1_cond $X=10.37 $Y=2.62
+ $X2=10.37 $Y2=3.59
r94 53 60 0.188114 $w=3.7e-07 $l=4.9e-07 $layer=MET1_cond $X=9.52 $Y=3.63
+ $X2=10.01 $Y2=3.63
r95 51 53 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.8 $Y=3.63
+ $X2=9.52 $Y2=3.63
r96 50 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.52 $Y=3.59
+ $X2=9.52 $Y2=3.59
r97 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.8 $Y=3.59 $X2=8.8
+ $Y2=3.59
r98 47 50 5.32947 $w=9.48e-07 $l=4.15e-07 $layer=LI1_cond $X=9.16 $Y=3.175
+ $X2=9.16 $Y2=3.59
r99 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.63 $Y=3.59
+ $X2=5.63 $Y2=3.59
r100 40 43 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.63 $Y=2.75
+ $X2=5.63 $Y2=3.59
r101 37 44 0.548985 $w=3.7e-07 $l=1.43e-06 $layer=MET1_cond $X=4.2 $Y=3.63
+ $X2=5.63 $Y2=3.63
r102 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.2 $Y=3.59
+ $X2=4.2 $Y2=3.59
r103 34 36 0.854342 $w=6.98e-07 $l=5e-08 $layer=LI1_cond $X=4.15 $Y=3.375
+ $X2=4.2 $Y2=3.375
r104 31 37 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.48 $Y=3.63
+ $X2=4.2 $Y2=3.63
r105 30 34 11.4482 $w=6.98e-07 $l=6.7e-07 $layer=LI1_cond $X=3.48 $Y=3.375
+ $X2=4.15 $Y2=3.375
r106 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.48 $Y=3.59
+ $X2=3.48 $Y2=3.59
r107 27 31 0.800443 $w=3.7e-07 $l=2.085e-06 $layer=MET1_cond $X=1.395 $Y=3.63
+ $X2=3.48 $Y2=3.63
r108 25 27 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.675 $Y=3.63
+ $X2=1.395 $Y2=3.63
r109 24 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.395 $Y=3.59
+ $X2=1.395 $Y2=3.59
r110 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.675 $Y=3.59
+ $X2=0.675 $Y2=3.59
r111 22 24 0.642105 $w=9.48e-07 $l=5e-08 $layer=LI1_cond $X=1.035 $Y=3.54
+ $X2=1.035 $Y2=3.59
r112 19 22 5.90737 $w=9.48e-07 $l=4.6e-07 $layer=LI1_cond $X=1.035 $Y=3.08
+ $X2=1.035 $Y2=3.54
r113 16 51 1.16707 $w=3.7e-07 $l=3.04e-06 $layer=MET1_cond $X=5.76 $Y=3.63
+ $X2=8.8 $Y2=3.63
r114 16 44 0.0499077 $w=3.7e-07 $l=1.3e-07 $layer=MET1_cond $X=5.76 $Y=3.63
+ $X2=5.63 $Y2=3.63
r115 5 59 400 $w=1.7e-07 $l=1.49708e-06 $layer=licon1_PDIFF $count=1 $X=10.19
+ $Y=2.215 $X2=10.445 $Y2=3.59
r116 5 56 400 $w=1.7e-07 $l=5.17011e-07 $layer=licon1_PDIFF $count=1 $X=10.19
+ $Y=2.215 $X2=10.445 $Y2=2.62
r117 4 47 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=9.33
+ $Y=2.965 $X2=9.47 $Y2=3.175
r118 3 40 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=5.485
+ $Y=2.625 $X2=5.63 $Y2=2.75
r119 2 34 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=4.01
+ $Y=2.935 $X2=4.15 $Y2=3.11
r120 1 22 600 $w=1.7e-07 $l=7.12881e-07 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=2.935 $X2=1.17 $Y2=3.54
r121 1 19 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=2.935 $X2=1.17 $Y2=3.08
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%A_489_107# 1 2 3 4 15 17 19 20 22 23 24 26
+ 27 30 31 32 34 35 36 38 39 40 44 46 50 52 56 57
c150 24 0 1.52001e-19 $X=3.685 $Y=1.26
c151 22 0 7.10574e-20 $X=3.6 $Y=1.175
r152 56 57 9.48656 $w=4.93e-07 $l=1.65e-07 $layer=LI1_cond $X=7.002 $Y=3.09
+ $X2=7.002 $Y2=2.925
r153 54 57 127.219 $w=1.68e-07 $l=1.95e-06 $layer=LI1_cond $X=6.84 $Y=0.975
+ $X2=6.84 $Y2=2.925
r154 52 54 10.3829 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.76 $Y=0.755
+ $X2=6.76 $Y2=0.975
r155 46 48 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.745
+ $X2=2.585 $Y2=0.83
r156 43 56 1.98138 $w=4.93e-07 $l=8.2e-08 $layer=LI1_cond $X=7.002 $Y=3.172
+ $X2=7.002 $Y2=3.09
r157 43 44 10.221 $w=4.93e-07 $l=4.23e-07 $layer=LI1_cond $X=7.002 $Y=3.172
+ $X2=7.002 $Y2=3.595
r158 39 44 9.18857 $w=1.7e-07 $l=2.86363e-07 $layer=LI1_cond $X=6.755 $Y=3.68
+ $X2=7.002 $Y2=3.595
r159 39 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.755 $Y=3.68
+ $X2=6.065 $Y2=3.68
r160 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.98 $Y=3.595
+ $X2=6.065 $Y2=3.68
r161 37 38 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=5.98 $Y=2.405
+ $X2=5.98 $Y2=3.595
r162 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.895 $Y=2.32
+ $X2=5.98 $Y2=2.405
r163 35 36 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.895 $Y=2.32
+ $X2=5.365 $Y2=2.32
r164 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.28 $Y=2.405
+ $X2=5.365 $Y2=2.32
r165 33 34 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=5.28 $Y=2.405
+ $X2=5.28 $Y2=3.635
r166 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.195 $Y=3.72
+ $X2=5.28 $Y2=3.635
r167 31 32 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.195 $Y=3.72
+ $X2=4.665 $Y2=3.72
r168 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.58 $Y=3.635
+ $X2=4.665 $Y2=3.72
r169 29 30 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.58 $Y=2.845
+ $X2=4.58 $Y2=3.635
r170 28 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.2 $Y=2.76
+ $X2=4.115 $Y2=2.76
r171 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.495 $Y=2.76
+ $X2=4.58 $Y2=2.845
r172 27 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.495 $Y=2.76
+ $X2=4.2 $Y2=2.76
r173 26 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=2.675
+ $X2=4.115 $Y2=2.76
r174 25 26 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=4.115 $Y=1.345
+ $X2=4.115 $Y2=2.675
r175 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.03 $Y=1.26
+ $X2=4.115 $Y2=1.345
r176 23 24 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.03 $Y=1.26
+ $X2=3.685 $Y2=1.26
r177 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.6 $Y=1.175
+ $X2=3.685 $Y2=1.26
r178 21 22 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.6 $Y=0.915
+ $X2=3.6 $Y2=1.175
r179 19 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.03 $Y=2.76
+ $X2=4.115 $Y2=2.76
r180 19 20 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=4.03 $Y=2.76
+ $X2=2.825 $Y2=2.76
r181 18 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=0.83
+ $X2=2.585 $Y2=0.83
r182 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.515 $Y=0.83
+ $X2=3.6 $Y2=0.915
r183 17 18 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.515 $Y=0.83
+ $X2=2.75 $Y2=0.83
r184 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.7 $Y=2.845
+ $X2=2.825 $Y2=2.76
r185 13 15 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=2.7 $Y=2.845
+ $X2=2.7 $Y2=3.06
r186 4 56 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=6.94
+ $Y=2.965 $X2=7.085 $Y2=3.09
r187 3 15 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.52
+ $Y=2.935 $X2=2.66 $Y2=3.06
r188 2 52 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=6.635
+ $Y=0.535 $X2=6.76 $Y2=0.755
r189 1 46 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.445
+ $Y=0.535 $X2=2.585 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%Q 1 2 7 8 9 10 11 12 13 22
r15 13 40 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=11.23 $Y=3.145
+ $X2=11.23 $Y2=3.59
r16 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=11.23 $Y=2.775
+ $X2=11.23 $Y2=3.145
r17 11 12 14.7445 $w=3.38e-07 $l=4.35e-07 $layer=LI1_cond $X=11.23 $Y=2.34
+ $X2=11.23 $Y2=2.775
r18 10 11 10.3381 $w=3.38e-07 $l=3.05e-07 $layer=LI1_cond $X=11.23 $Y=2.035
+ $X2=11.23 $Y2=2.34
r19 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=11.23 $Y=1.665
+ $X2=11.23 $Y2=2.035
r20 8 9 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=11.23 $Y=1.295
+ $X2=11.23 $Y2=1.665
r21 7 8 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=11.23 $Y=0.925
+ $X2=11.23 $Y2=1.295
r22 7 22 8.30437 $w=3.38e-07 $l=2.45e-07 $layer=LI1_cond $X=11.23 $Y=0.925
+ $X2=11.23 $Y2=0.68
r23 2 40 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=11.085
+ $Y=2.215 $X2=11.225 $Y2=3.59
r24 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=11.085
+ $Y=2.215 $X2=11.225 $Y2=2.34
r25 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.095
+ $Y=0.535 $X2=11.235 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__SDLXTP_1%VGND 1 2 3 4 5 16 19 28 35 48 52 56
r88 58 60 5.90737 $w=9.48e-07 $l=4.6e-07 $layer=LI1_cond $X=10.4 $Y=0.68
+ $X2=10.4 $Y2=1.14
r89 53 56 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.04 $Y=0.44
+ $X2=10.76 $Y2=0.44
r90 52 58 2.56842 $w=9.48e-07 $l=2e-07 $layer=LI1_cond $X=10.4 $Y=0.48 $X2=10.4
+ $Y2=0.68
r91 52 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.76 $Y=0.48
+ $X2=10.76 $Y2=0.48
r92 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.04 $Y=0.48
+ $X2=10.04 $Y2=0.48
r93 49 53 0.368549 $w=3.7e-07 $l=9.6e-07 $layer=MET1_cond $X=9.08 $Y=0.44
+ $X2=10.04 $Y2=0.44
r94 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.08 $Y=0.48
+ $X2=9.08 $Y2=0.48
r95 46 48 1.12838 $w=5.28e-07 $l=5e-08 $layer=LI1_cond $X=9.03 $Y=0.63 $X2=9.08
+ $Y2=0.63
r96 43 49 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.36 $Y=0.44
+ $X2=9.08 $Y2=0.44
r97 42 46 15.1202 $w=5.28e-07 $l=6.7e-07 $layer=LI1_cond $X=8.36 $Y=0.63
+ $X2=9.03 $Y2=0.63
r98 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.36 $Y=0.48
+ $X2=8.36 $Y2=0.48
r99 35 39 5.37222 $w=5.88e-07 $l=2.65e-07 $layer=LI1_cond $X=5.5 $Y=0.48 $X2=5.5
+ $Y2=0.745
r100 28 32 5.37222 $w=5.88e-07 $l=2.65e-07 $layer=LI1_cond $X=4.16 $Y=0.48
+ $X2=4.16 $Y2=0.745
r101 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.34 $Y=0.48
+ $X2=4.34 $Y2=0.48
r102 23 29 1.09221 $w=3.7e-07 $l=2.845e-06 $layer=MET1_cond $X=1.495 $Y=0.44
+ $X2=4.34 $Y2=0.44
r103 20 23 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.775 $Y=0.44
+ $X2=1.495 $Y2=0.44
r104 19 25 3.40316 $w=9.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.135 $Y=0.48
+ $X2=1.135 $Y2=0.745
r105 19 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.495 $Y=0.48
+ $X2=1.495 $Y2=0.48
r106 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.775 $Y=0.48
+ $X2=0.775 $Y2=0.48
r107 16 43 1.02887 $w=3.7e-07 $l=2.68e-06 $layer=MET1_cond $X=5.68 $Y=0.44
+ $X2=8.36 $Y2=0.44
r108 16 29 0.514433 $w=3.7e-07 $l=1.34e-06 $layer=MET1_cond $X=5.68 $Y=0.44
+ $X2=4.34 $Y2=0.44
r109 16 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.68 $Y=0.48
+ $X2=5.68 $Y2=0.48
r110 5 60 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=10.22
+ $Y=0.865 $X2=10.455 $Y2=1.14
r111 5 58 182 $w=1.7e-07 $l=3.14166e-07 $layer=licon1_NDIFF $count=1 $X=10.22
+ $Y=0.865 $X2=10.455 $Y2=0.68
r112 4 46 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.89
+ $Y=0.535 $X2=9.03 $Y2=0.745
r113 3 39 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.285
+ $Y=0.535 $X2=5.43 $Y2=0.745
r114 2 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.535 $X2=4.075 $Y2=0.745
r115 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.955
+ $Y=0.535 $X2=1.095 $Y2=0.745
.ends

