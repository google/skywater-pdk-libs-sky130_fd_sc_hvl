# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__a21o_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__a21o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.805000 1.505000 3.715000 1.835000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.895000 1.505000 4.195000 1.835000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.505000 2.275000 1.750000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.611250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.495000 0.460000 1.325000 ;
        RECT 0.110000 1.325000 0.360000 3.735000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 4.320000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 4.320000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 4.320000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 4.320000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.985000 4.320000 4.155000 ;
      RECT 0.540000  2.280000 1.440000 3.755000 ;
      RECT 0.565000  1.725000 0.895000 1.930000 ;
      RECT 0.565000  1.930000 2.625000 2.100000 ;
      RECT 0.640000  0.365000 2.250000 1.325000 ;
      RECT 1.620000  2.100000 1.870000 3.755000 ;
      RECT 2.320000  2.280000 4.210000 2.450000 ;
      RECT 2.320000  2.450000 2.650000 3.755000 ;
      RECT 2.430000  0.495000 2.680000 1.325000 ;
      RECT 2.455000  1.325000 2.625000 1.930000 ;
      RECT 2.830000  2.630000 3.780000 3.755000 ;
      RECT 2.860000  0.365000 4.170000 1.325000 ;
      RECT 3.960000  2.195000 4.210000 2.280000 ;
      RECT 3.960000  2.450000 4.210000 3.735000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.545000  3.505000 0.715000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.640000  0.395000 0.810000 0.565000 ;
      RECT 0.905000  3.505000 1.075000 3.675000 ;
      RECT 1.000000  0.395000 1.170000 0.565000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.265000  3.505000 1.435000 3.675000 ;
      RECT 1.360000  0.395000 1.530000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.720000  0.395000 1.890000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.080000  0.395000 2.250000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.860000  3.505000 3.030000 3.675000 ;
      RECT 2.890000  0.395000 3.060000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.220000  3.505000 3.390000 3.675000 ;
      RECT 3.250000  0.395000 3.420000 0.565000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.580000  3.505000 3.750000 3.675000 ;
      RECT 3.610000  0.395000 3.780000 0.565000 ;
      RECT 3.970000  0.395000 4.140000 0.565000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
  END
END sky130_fd_sc_hvl__a21o_1
