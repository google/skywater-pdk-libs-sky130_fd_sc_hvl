# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__xnor2_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__xnor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  2.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.580000 2.060000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 1.725000 0.905000 1.930000 ;
        RECT 0.575000 1.930000 3.255000 2.100000 ;
        RECT 1.565000 2.100000 3.255000 2.120000 ;
        RECT 2.925000 1.805000 3.255000 1.930000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.481250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.025000 1.905000 5.155000 2.075000 ;
        RECT 4.025000 2.075000 4.275000 3.755000 ;
        RECT 4.445000 1.545000 5.155000 1.905000 ;
        RECT 4.750000 0.535000 5.155000 1.545000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.610000 0.365000 2.410000 1.050000 ;
        RECT 3.100000 0.365000 3.630000 0.925000 ;
      LAYER mcon ;
        RECT 0.800000 0.395000 0.970000 0.565000 ;
        RECT 1.160000 0.395000 1.330000 0.565000 ;
        RECT 1.520000 0.395000 1.690000 0.565000 ;
        RECT 1.880000 0.395000 2.050000 0.565000 ;
        RECT 2.240000 0.395000 2.410000 0.565000 ;
        RECT 3.100000 0.395000 3.270000 0.565000 ;
        RECT 3.460000 0.395000 3.630000 0.565000 ;
      LAYER met1 ;
        RECT 0.000000 0.255000 5.280000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.115000 5.280000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 5.280000 4.155000 ;
      LAYER mcon ;
        RECT 0.155000 3.985000 0.325000 4.155000 ;
        RECT 0.635000 3.985000 0.805000 4.155000 ;
        RECT 1.115000 3.985000 1.285000 4.155000 ;
        RECT 1.595000 3.985000 1.765000 4.155000 ;
        RECT 2.075000 3.985000 2.245000 4.155000 ;
        RECT 2.555000 3.985000 2.725000 4.155000 ;
        RECT 3.035000 3.985000 3.205000 4.155000 ;
        RECT 3.515000 3.985000 3.685000 4.155000 ;
        RECT 3.995000 3.985000 4.165000 4.155000 ;
        RECT 4.475000 3.985000 4.645000 4.155000 ;
        RECT 4.955000 3.985000 5.125000 4.155000 ;
      LAYER met1 ;
        RECT 0.000000 3.955000 5.280000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.090000 2.630000 0.985000 3.755000 ;
        RECT 1.515000 2.300000 3.845000 3.755000 ;
        RECT 4.465000 2.255000 5.055000 3.755000 ;
      LAYER mcon ;
        RECT 0.095000 3.505000 0.265000 3.675000 ;
        RECT 0.455000 3.505000 0.625000 3.675000 ;
        RECT 0.815000 3.505000 0.985000 3.675000 ;
        RECT 1.515000 3.505000 1.685000 3.675000 ;
        RECT 1.875000 3.505000 2.045000 3.675000 ;
        RECT 2.235000 3.505000 2.405000 3.675000 ;
        RECT 2.595000 3.505000 2.765000 3.675000 ;
        RECT 2.955000 3.505000 3.125000 3.675000 ;
        RECT 3.315000 3.505000 3.485000 3.675000 ;
        RECT 3.675000 3.505000 3.845000 3.675000 ;
        RECT 4.495000 3.505000 4.665000 3.675000 ;
        RECT 4.855000 3.505000 5.025000 3.675000 ;
      LAYER met1 ;
        RECT 0.000000 3.445000 5.280000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.110000 0.495000 0.440000 1.230000 ;
      RECT 0.110000 1.230000 2.410000 1.400000 ;
      RECT 0.110000 1.400000 0.360000 2.280000 ;
      RECT 0.110000 2.280000 1.335000 2.450000 ;
      RECT 1.165000 2.450000 1.335000 3.755000 ;
      RECT 2.240000 1.400000 2.410000 1.455000 ;
      RECT 2.240000 1.455000 3.980000 1.625000 ;
      RECT 2.590000 0.495000 2.920000 1.105000 ;
      RECT 2.590000 1.105000 4.300000 1.285000 ;
      RECT 3.650000 1.625000 3.980000 1.725000 ;
      RECT 3.970000 0.535000 4.300000 1.105000 ;
  END
END sky130_fd_sc_hvl__xnor2_1
