* File: sky130_fd_sc_hvl__xor2_1.pex.spice
* Created: Fri Aug 28 09:40:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__XOR2_1%VNB 5 7 11 25
r31 7 25 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=0.057
+ $X2=2.64 $Y2=0.058
r32 7 11 0.00134943 $w=5.28e-06 $l=5.7e-08 $layer=MET1_cond $X=2.64 $Y=0.057
+ $X2=2.64 $Y2=0
r33 5 11 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r34 5 11 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__XOR2_1%VPB 4 6 14 21
r45 10 21 0.00134943 $w=5.28e-06 $l=5.7e-08 $layer=MET1_cond $X=2.64 $Y=4.07
+ $X2=2.64 $Y2=4.013
r46 10 14 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=4.07
+ $X2=5.04 $Y2=4.07
r47 9 14 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=5.04
+ $Y2=4.07
r48 9 10 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r49 6 21 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=4.012
+ $X2=2.64 $Y2=4.013
r50 4 14 33.0909 $w=1.7e-07 $l=5.08232e-06 $layer=licon1_NTAP_notbjt $count=5
+ $X=0 $Y=3.985 $X2=5.04 $Y2=4.07
r51 4 9 33.0909 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=5
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__XOR2_1%B 1 3 7 9 15 16 17 18 21 25 28
r66 28 31 81.3245 $w=5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.545 $Y=0.91
+ $X2=3.545 $Y2=1.67
r67 18 33 6.90146 $w=2.74e-07 $l=1.55e-07 $layer=LI1_cond $X=3.565 $Y=1.665
+ $X2=3.565 $Y2=1.51
r68 18 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.565
+ $Y=1.67 $X2=3.565 $Y2=1.67
r69 16 33 3.52985 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.415 $Y=1.51
+ $X2=3.565 $Y2=1.51
r70 16 17 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=3.415 $Y=1.51
+ $X2=1.51 $Y2=1.51
r71 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.425 $Y=1.595
+ $X2=1.51 $Y2=1.51
r72 14 15 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.425 $Y=1.595
+ $X2=1.425 $Y2=1.775
r73 12 25 115.031 $w=5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.685 $Y=1.89
+ $X2=0.685 $Y2=2.965
r74 12 21 104.866 $w=5e-07 $l=9.8e-07 $layer=POLY_cond $X=0.685 $Y=1.89
+ $X2=0.685 $Y2=0.91
r75 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.725
+ $Y=1.89 $X2=0.725 $Y2=1.89
r76 9 15 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.34 $Y=1.915
+ $X2=1.425 $Y2=1.775
r77 9 11 25.3126 $w=2.78e-07 $l=6.15e-07 $layer=LI1_cond $X=1.34 $Y=1.915
+ $X2=0.725 $Y2=1.915
r78 7 31 19.7961 $w=5e-07 $l=1.85e-07 $layer=POLY_cond $X=3.545 $Y=1.855
+ $X2=3.545 $Y2=1.67
r79 1 7 89.4433 $w=2.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.185 $Y=1.98
+ $X2=3.545 $Y2=1.98
r80 1 3 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.185 $Y=2.105 $X2=3.185
+ $Y2=2.965
.ends

.subckt PM_SKY130_FD_SC_HVL__XOR2_1%A 1 3 6 8 10 11 13 14 15 16 25
c48 16 0 1.62409e-19 $X=3.12 $Y=2.035
r49 23 25 5.39243 $w=5.81e-07 $l=6.5e-08 $layer=POLY_cond $X=2.34 $Y=1.75
+ $X2=2.405 $Y2=1.75
r50 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.34
+ $Y=1.89 $X2=2.34 $Y2=1.89
r51 21 23 72.5904 $w=5.81e-07 $l=8.75e-07 $layer=POLY_cond $X=1.465 $Y=1.75
+ $X2=2.34 $Y2=1.75
r52 20 21 5.80723 $w=5.81e-07 $l=7e-08 $layer=POLY_cond $X=1.395 $Y=1.75
+ $X2=1.465 $Y2=1.75
r53 15 16 14.7513 $w=3.73e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.962
+ $X2=3.12 $Y2=1.962
r54 15 24 9.21954 $w=3.73e-07 $l=3e-07 $layer=LI1_cond $X=2.64 $Y=1.962 $X2=2.34
+ $Y2=1.962
r55 14 24 5.53173 $w=3.73e-07 $l=1.8e-07 $layer=LI1_cond $X=2.16 $Y=1.962
+ $X2=2.34 $Y2=1.962
r56 11 25 35.673 $w=5.81e-07 $l=5.80991e-07 $layer=POLY_cond $X=2.835 $Y=1.395
+ $X2=2.405 $Y2=1.75
r57 11 13 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.835 $Y=1.395
+ $X2=2.835 $Y2=0.91
r58 8 25 6.38776 $w=5e-07 $l=3.55e-07 $layer=POLY_cond $X=2.405 $Y=2.105
+ $X2=2.405 $Y2=1.75
r59 8 10 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.405 $Y=2.105 $X2=2.405
+ $Y2=2.965
r60 4 21 6.38776 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.465 $Y=1.415
+ $X2=1.465 $Y2=1.75
r61 4 6 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.465 $Y=1.415 $X2=1.465
+ $Y2=0.91
r62 1 20 6.38776 $w=5e-07 $l=3.55e-07 $layer=POLY_cond $X=1.395 $Y=2.105
+ $X2=1.395 $Y2=1.75
r63 1 3 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.395 $Y=2.105 $X2=1.395
+ $Y2=2.965
.ends

.subckt PM_SKY130_FD_SC_HVL__XOR2_1%A_30_443# 1 2 9 11 13 17 20 24 25 26 30 32
+ 35 36 37 42 43
c78 32 0 1.62409e-19 $X=4.55 $Y=2.69
r79 46 48 28.8916 $w=5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.325 $Y=1.855
+ $X2=4.595 $Y2=1.855
r80 43 48 12.8407 $w=5e-07 $l=1.2e-07 $layer=POLY_cond $X=4.715 $Y=1.855
+ $X2=4.595 $Y2=1.855
r81 42 45 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=1.83
+ $X2=4.715 $Y2=1.995
r82 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.715
+ $Y=1.83 $X2=4.715 $Y2=1.83
r83 37 39 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.145 $Y=2.52
+ $X2=3.145 $Y2=2.69
r84 35 45 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.635 $Y=2.605
+ $X2=4.635 $Y2=1.995
r85 33 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.23 $Y=2.69
+ $X2=3.145 $Y2=2.69
r86 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.55 $Y=2.69
+ $X2=4.635 $Y2=2.605
r87 32 33 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=4.55 $Y=2.69
+ $X2=3.23 $Y2=2.69
r88 28 30 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=1.035 $Y=1.425
+ $X2=1.035 $Y2=0.66
r89 27 36 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.38 $Y=2.52
+ $X2=0.255 $Y2=2.52
r90 26 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=2.52
+ $X2=3.145 $Y2=2.52
r91 26 27 174.845 $w=1.68e-07 $l=2.68e-06 $layer=LI1_cond $X=3.06 $Y=2.52
+ $X2=0.38 $Y2=2.52
r92 24 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.91 $Y=1.51
+ $X2=1.035 $Y2=1.425
r93 24 25 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.91 $Y=1.51
+ $X2=0.38 $Y2=1.51
r94 20 22 38.4916 $w=2.48e-07 $l=8.35e-07 $layer=LI1_cond $X=0.255 $Y=2.755
+ $X2=0.255 $Y2=3.59
r95 18 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=2.605
+ $X2=0.255 $Y2=2.52
r96 18 20 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=0.255 $Y=2.605
+ $X2=0.255 $Y2=2.755
r97 15 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=2.435
+ $X2=0.255 $Y2=2.52
r98 15 17 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=0.255 $Y=2.435
+ $X2=0.255 $Y2=2.34
r99 14 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.255 $Y=1.595
+ $X2=0.38 $Y2=1.51
r100 14 17 34.3428 $w=2.48e-07 $l=7.45e-07 $layer=LI1_cond $X=0.255 $Y=1.595
+ $X2=0.255 $Y2=2.34
r101 11 48 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.595 $Y=2.105
+ $X2=4.595 $Y2=1.855
r102 11 13 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.595 $Y=2.105
+ $X2=4.595 $Y2=2.965
r103 7 46 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.325 $Y=1.605
+ $X2=4.325 $Y2=1.855
r104 7 9 74.3691 $w=5e-07 $l=6.95e-07 $layer=POLY_cond $X=4.325 $Y=1.605
+ $X2=4.325 $Y2=0.91
r105 2 22 400 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.215 $X2=0.295 $Y2=3.59
r106 2 20 400 $w=1.7e-07 $l=6.08194e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.215 $X2=0.295 $Y2=2.755
r107 2 17 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.215 $X2=0.295 $Y2=2.34
r108 1 30 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.935
+ $Y=0.535 $X2=1.075 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__XOR2_1%VPWR 1 2 7 10 26 27
r37 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.61 $Y=3.59
+ $X2=4.61 $Y2=3.59
r38 24 26 27.5098 $w=4.48e-07 $l=1.035e-06 $layer=LI1_cond $X=3.575 $Y=3.53
+ $X2=4.61 $Y2=3.53
r39 21 27 0.552824 $w=3.7e-07 $l=1.44e-06 $layer=MET1_cond $X=3.17 $Y=3.63
+ $X2=4.61 $Y2=3.63
r40 20 24 10.7647 $w=4.48e-07 $l=4.05e-07 $layer=LI1_cond $X=3.17 $Y=3.53
+ $X2=3.575 $Y2=3.53
r41 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.17 $Y=3.59
+ $X2=3.17 $Y2=3.59
r42 14 17 0.69103 $w=3.7e-07 $l=1.8e-06 $layer=MET1_cond $X=0.645 $Y=3.63
+ $X2=2.445 $Y2=3.63
r43 13 17 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.445 $Y=3.59
+ $X2=2.445 $Y2=3.59
r44 13 14 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.645 $Y=3.59
+ $X2=0.645 $Y2=3.59
r45 10 13 4.45888 $w=1.968e-06 $l=7.2e-07 $layer=LI1_cond $X=1.545 $Y=2.87
+ $X2=1.545 $Y2=3.59
r46 7 21 0.20347 $w=3.7e-07 $l=5.3e-07 $layer=MET1_cond $X=2.64 $Y=3.63 $X2=3.17
+ $Y2=3.63
r47 7 17 0.0748616 $w=3.7e-07 $l=1.95e-07 $layer=MET1_cond $X=2.64 $Y=3.63
+ $X2=2.445 $Y2=3.63
r48 2 24 600 $w=1.7e-07 $l=1.34318e-06 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=2.215 $X2=3.575 $Y2=3.49
r49 1 13 400 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=2.215 $X2=1.785 $Y2=3.59
r50 1 10 400 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=2.215 $X2=1.785 $Y2=2.87
.ends

.subckt PM_SKY130_FD_SC_HVL__XOR2_1%A_531_443# 1 2 7 9 11 15 19 23
r32 17 23 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=3.125
+ $X2=5.025 $Y2=3.04
r33 17 19 2.30489 $w=2.48e-07 $l=5e-08 $layer=LI1_cond $X=5.025 $Y=3.125
+ $X2=5.025 $Y2=3.175
r34 13 23 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=2.955
+ $X2=5.025 $Y2=3.04
r35 13 15 28.3501 $w=2.48e-07 $l=6.15e-07 $layer=LI1_cond $X=5.025 $Y=2.955
+ $X2=5.025 $Y2=2.34
r36 12 22 3.40825 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.88 $Y=3.04
+ $X2=2.795 $Y2=2.955
r37 11 23 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.9 $Y=3.04
+ $X2=5.025 $Y2=3.04
r38 11 12 131.786 $w=1.68e-07 $l=2.02e-06 $layer=LI1_cond $X=4.9 $Y=3.04
+ $X2=2.88 $Y2=3.04
r39 7 22 3.40825 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.795 $Y=3.125
+ $X2=2.795 $Y2=2.955
r40 7 9 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.795 $Y=3.125
+ $X2=2.795 $Y2=3.59
r41 2 19 300 $w=1.7e-07 $l=1.02762e-06 $layer=licon1_PDIFF $count=2 $X=4.845
+ $Y=2.215 $X2=4.985 $Y2=3.175
r42 2 15 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.845
+ $Y=2.215 $X2=4.985 $Y2=2.34
r43 1 22 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=2.655
+ $Y=2.215 $X2=2.795 $Y2=2.95
r44 1 9 600 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=1 $X=2.655
+ $Y=2.215 $X2=2.795 $Y2=3.59
.ends

.subckt PM_SKY130_FD_SC_HVL__XOR2_1%X 1 2 7 8 9 10 18 33
r21 33 34 1.30711 $w=5.18e-07 $l=3e-08 $layer=LI1_cond $X=4.11 $Y=1.295 $X2=4.11
+ $Y2=1.325
r22 10 29 8.67889 $w=4.03e-07 $l=3.05e-07 $layer=LI1_cond $X=4.167 $Y=2.035
+ $X2=4.167 $Y2=2.34
r23 9 10 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=4.167 $Y=1.665
+ $X2=4.167 $Y2=2.035
r24 8 33 0.644042 $w=5.18e-07 $l=2.8e-08 $layer=LI1_cond $X=4.11 $Y=1.267
+ $X2=4.11 $Y2=1.295
r25 8 16 4.6463 $w=5.18e-07 $l=2.02e-07 $layer=LI1_cond $X=4.11 $Y=1.267
+ $X2=4.11 $Y2=1.065
r26 8 9 8.90654 $w=4.03e-07 $l=3.13e-07 $layer=LI1_cond $X=4.167 $Y=1.352
+ $X2=4.167 $Y2=1.665
r27 8 34 0.768295 $w=4.03e-07 $l=2.7e-08 $layer=LI1_cond $X=4.167 $Y=1.352
+ $X2=4.167 $Y2=1.325
r28 7 16 3.22021 $w=5.18e-07 $l=1.4e-07 $layer=LI1_cond $X=4.11 $Y=0.925
+ $X2=4.11 $Y2=1.065
r29 7 18 6.0954 $w=5.18e-07 $l=2.65e-07 $layer=LI1_cond $X=4.11 $Y=0.925
+ $X2=4.11 $Y2=0.66
r30 2 29 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.06
+ $Y=2.215 $X2=4.205 $Y2=2.34
r31 1 18 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.795
+ $Y=0.535 $X2=3.935 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__XOR2_1%VGND 1 2 3 10 13 26 30 31
r37 30 34 3.64905 $w=5.88e-07 $l=1.8e-07 $layer=LI1_cond $X=4.845 $Y=0.48
+ $X2=4.845 $Y2=0.66
r38 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.025 $Y=0.48
+ $X2=5.025 $Y2=0.48
r39 27 31 0.552824 $w=3.7e-07 $l=1.44e-06 $layer=MET1_cond $X=3.585 $Y=0.44
+ $X2=5.025 $Y2=0.44
r40 26 27 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.585 $Y=0.48
+ $X2=3.585 $Y2=0.48
r41 24 26 23.9841 $w=8.78e-07 $l=1.73e-06 $layer=LI1_cond $X=1.855 $Y=0.805
+ $X2=3.585 $Y2=0.805
r42 20 24 5.96136 $w=8.78e-07 $l=4.3e-07 $layer=LI1_cond $X=1.425 $Y=0.805
+ $X2=1.855 $Y2=0.805
r43 20 21 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.425 $Y=0.48
+ $X2=1.425 $Y2=0.48
r44 14 21 0.330159 $w=3.7e-07 $l=8.6e-07 $layer=MET1_cond $X=0.565 $Y=0.44
+ $X2=1.425 $Y2=0.44
r45 13 17 3.64905 $w=5.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.385 $Y=0.48
+ $X2=0.385 $Y2=0.66
r46 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.565 $Y=0.48
+ $X2=0.565 $Y2=0.48
r47 10 27 0.362791 $w=3.7e-07 $l=9.45e-07 $layer=MET1_cond $X=2.64 $Y=0.44
+ $X2=3.585 $Y2=0.44
r48 10 21 0.466445 $w=3.7e-07 $l=1.215e-06 $layer=MET1_cond $X=2.64 $Y=0.44
+ $X2=1.425 $Y2=0.44
r49 3 34 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.575
+ $Y=0.535 $X2=4.715 $Y2=0.66
r50 2 24 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.715
+ $Y=0.535 $X2=1.855 $Y2=0.66
r51 1 17 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.535 $X2=0.295 $Y2=0.66
.ends

