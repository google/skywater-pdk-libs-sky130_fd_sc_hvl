* File: sky130_fd_sc_hvl__dfxbp_1.pex.spice
* Created: Fri Aug 28 09:34:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%VNB 5 7 11
r99 7 11 0.000511853 $w=1.392e-05 $l=5.7e-08 $layer=MET1_cond $X=6.96 $Y=0.057
+ $X2=6.96 $Y2=0
r100 5 11 0.641379 $w=1.7e-07 $l=2.465e-06 $layer=mcon $count=14 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r101 5 11 0.641379 $w=1.7e-07 $l=2.465e-06 $layer=mcon $count=14 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%VPB 4 6 14
c134 4 0 1.77943e-19 $X=-0.33 $Y=1.885
r135 10 14 0.641379 $w=1.7e-07 $l=2.465e-06 $layer=mcon $count=14 $X=13.68
+ $Y=4.07 $X2=13.68 $Y2=4.07
r136 9 14 876.834 $w=1.68e-07 $l=1.344e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=13.68 $Y2=4.07
r137 9 10 0.641379 $w=1.7e-07 $l=2.465e-06 $layer=mcon $count=14 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r138 6 10 0.000511853 $w=1.392e-05 $l=5.7e-08 $layer=MET1_cond $X=6.96 $Y=4.013
+ $X2=6.96 $Y2=4.07
r139 4 14 12.5517 $w=1.7e-07 $l=1.37224e-05 $layer=licon1_NTAP_notbjt $count=14
+ $X=0 $Y=3.985 $X2=13.68 $Y2=4.07
r140 4 9 12.5517 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=14
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%CLK 3 7 9 10 14
r30 14 17 61.2197 $w=5.2e-07 $l=5.95e-07 $layer=POLY_cond $X=0.675 $Y=1.715
+ $X2=0.675 $Y2=2.31
r31 14 16 19.0347 $w=5.2e-07 $l=1.85e-07 $layer=POLY_cond $X=0.675 $Y=1.715
+ $X2=0.675 $Y2=1.53
r32 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.725 $Y=1.665
+ $X2=0.725 $Y2=2.035
r33 9 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.725
+ $Y=1.715 $X2=0.725 $Y2=1.715
r34 7 17 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.685 $Y=2.815
+ $X2=0.685 $Y2=2.31
r35 3 16 81.3245 $w=5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.665 $Y=0.77 $X2=0.665
+ $Y2=1.53
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%A_30_112# 1 2 9 13 15 17 18 20 23 26 30 32
+ 34 35 37 38 39 41 42 43 45 46 47 50 54 55 59 63 64 67 68 69 71 72 76 77 79 82
+ 84 85 86 90 91 93 97 105
c251 105 0 7.03008e-20 $X=8.08 $Y=1.085
c252 90 0 1.65371e-19 $X=7.26 $Y=2.37
c253 86 0 8.31313e-20 $X=4.92 $Y=2.72
c254 64 0 1.29366e-20 $X=6.395 $Y=2.72
c255 50 0 1.57779e-19 $X=3.965 $Y=1.28
r256 91 97 88.2799 $w=5e-07 $l=8.25e-07 $layer=POLY_cond $X=7.22 $Y=2.37
+ $X2=7.22 $Y2=3.195
r257 90 91 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.26
+ $Y=2.37 $X2=7.26 $Y2=2.37
r258 87 90 3.17915 $w=2.88e-07 $l=8e-08 $layer=LI1_cond $X=7.18 $Y=2.35 $X2=7.26
+ $Y2=2.35
r259 82 101 54.0174 $w=5.2e-07 $l=5.25e-07 $layer=POLY_cond $X=1.455 $Y=1.365
+ $X2=1.455 $Y2=1.89
r260 82 100 26.237 $w=5.2e-07 $l=2.55e-07 $layer=POLY_cond $X=1.455 $Y=1.365
+ $X2=1.455 $Y2=1.11
r261 81 82 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.38
+ $Y=1.365 $X2=1.38 $Y2=1.365
r262 77 105 18.6756 $w=5.3e-07 $l=1.85e-07 $layer=POLY_cond $X=8.08 $Y=1.27
+ $X2=8.08 $Y2=1.085
r263 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.11
+ $Y=1.27 $X2=8.11 $Y2=1.27
r264 74 76 100.945 $w=2.68e-07 $l=2.365e-06 $layer=LI1_cond $X=8.11 $Y=3.635
+ $X2=8.11 $Y2=1.27
r265 73 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.265 $Y=3.72
+ $X2=7.18 $Y2=3.72
r266 72 74 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=7.975 $Y=3.72
+ $X2=8.11 $Y2=3.635
r267 72 73 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.975 $Y=3.72
+ $X2=7.265 $Y2=3.72
r268 71 93 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=3.635
+ $X2=7.18 $Y2=3.72
r269 70 87 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.18 $Y=2.495
+ $X2=7.18 $Y2=2.35
r270 70 71 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=7.18 $Y=2.495
+ $X2=7.18 $Y2=3.635
r271 68 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.095 $Y=3.72
+ $X2=7.18 $Y2=3.72
r272 68 69 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.095 $Y=3.72
+ $X2=6.565 $Y2=3.72
r273 67 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.48 $Y=3.635
+ $X2=6.565 $Y2=3.72
r274 66 67 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=6.48 $Y=2.805
+ $X2=6.48 $Y2=3.635
r275 65 86 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.085 $Y=2.72
+ $X2=4.92 $Y2=2.72
r276 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.395 $Y=2.72
+ $X2=6.48 $Y2=2.805
r277 64 65 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=6.395 $Y=2.72
+ $X2=5.085 $Y2=2.72
r278 62 86 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.92 $Y=2.805
+ $X2=4.92 $Y2=2.72
r279 62 63 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=4.92 $Y=2.805
+ $X2=4.92 $Y2=3.335
r280 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.92
+ $Y=2.37 $X2=4.92 $Y2=2.37
r281 57 86 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.92 $Y=2.635
+ $X2=4.92 $Y2=2.72
r282 57 59 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=4.92 $Y=2.635
+ $X2=4.92 $Y2=2.37
r283 56 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=3.42
+ $X2=4.035 $Y2=3.42
r284 55 63 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.755 $Y=3.42
+ $X2=4.92 $Y2=3.335
r285 55 56 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.755 $Y=3.42
+ $X2=4.12 $Y2=3.42
r286 54 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=3.335
+ $X2=4.035 $Y2=3.42
r287 54 84 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=4.035 $Y=3.335
+ $X2=4.035 $Y2=1.785
r288 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.965
+ $Y=1.28 $X2=3.965 $Y2=1.28
r289 48 84 6.75802 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=4 $Y=1.665 $X2=4
+ $Y2=1.785
r290 48 50 18.4871 $w=2.38e-07 $l=3.85e-07 $layer=LI1_cond $X=4 $Y=1.665 $X2=4
+ $Y2=1.28
r291 46 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=3.42
+ $X2=4.035 $Y2=3.42
r292 46 47 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.95 $Y=3.42 $X2=3.35
+ $Y2=3.42
r293 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.265 $Y=3.335
+ $X2=3.35 $Y2=3.42
r294 44 45 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=3.265 $Y=2.475
+ $X2=3.265 $Y2=3.335
r295 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.18 $Y=2.39
+ $X2=3.265 $Y2=2.475
r296 42 43 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.18 $Y=2.39
+ $X2=2.29 $Y2=2.39
r297 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.205 $Y=2.475
+ $X2=2.29 $Y2=2.39
r298 40 41 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.205 $Y=2.475
+ $X2=2.205 $Y2=3.41
r299 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.12 $Y=3.495
+ $X2=2.205 $Y2=3.41
r300 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.12 $Y=3.495
+ $X2=1.51 $Y2=3.495
r301 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.425 $Y=3.41
+ $X2=1.51 $Y2=3.495
r302 37 83 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=1.425 $Y=3.41
+ $X2=1.425 $Y2=1.87
r303 35 83 7.64045 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.38 $Y=1.705
+ $X2=1.38 $Y2=1.87
r304 34 81 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.38 $Y=1.37 $X2=1.38
+ $Y2=1.285
r305 34 35 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.38 $Y=1.37
+ $X2=1.38 $Y2=1.705
r306 33 79 3.44808 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.44 $Y=1.285
+ $X2=0.275 $Y2=1.285
r307 32 81 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=1.285
+ $X2=1.38 $Y2=1.285
r308 32 33 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.215 $Y=1.285
+ $X2=0.44 $Y2=1.285
r309 28 79 3.14896 $w=3e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.245 $Y=1.37
+ $X2=0.275 $Y2=1.285
r310 28 30 51.0063 $w=2.68e-07 $l=1.195e-06 $layer=LI1_cond $X=0.245 $Y=1.37
+ $X2=0.245 $Y2=2.565
r311 24 79 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.275 $Y=1.2 $X2=0.275
+ $Y2=1.285
r312 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.275 $Y=1.2
+ $X2=0.275 $Y2=0.77
r313 23 105 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.095 $Y=0.765
+ $X2=8.095 $Y2=1.085
r314 18 60 27.4533 $w=5e-07 $l=2.75e-07 $layer=POLY_cond $X=4.855 $Y=2.645
+ $X2=4.855 $Y2=2.37
r315 18 20 25.064 $w=5e-07 $l=2.6e-07 $layer=POLY_cond $X=4.855 $Y=2.645
+ $X2=4.855 $Y2=2.905
r316 15 51 19.0043 $w=5e-07 $l=2.11778e-07 $layer=POLY_cond $X=4.075 $Y=1.085
+ $X2=4.04 $Y2=1.28
r317 15 17 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.075 $Y=1.085
+ $X2=4.075 $Y2=0.765
r318 13 101 98.9805 $w=5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.465 $Y=2.815
+ $X2=1.465 $Y2=1.89
r319 9 100 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.445 $Y=0.77
+ $X2=1.445 $Y2=1.11
r320 2 30 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.44 $X2=0.295 $Y2=2.565
r321 1 26 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.56 $X2=0.275 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%D 3 7 9 12 13 18 19
r43 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.185
+ $Y=1.665 $X2=3.185 $Y2=1.665
r44 13 19 11.239 $w=5.78e-07 $l=5.45e-07 $layer=LI1_cond $X=2.64 $Y=1.835
+ $X2=3.185 $Y2=1.835
r45 11 18 24.8371 $w=5.45e-07 $l=2.53e-07 $layer=POLY_cond $X=3.272 $Y=1.918
+ $X2=3.272 $Y2=1.665
r46 11 12 27.1636 $w=5.45e-07 $l=2.72e-07 $layer=POLY_cond $X=3.272 $Y=1.918
+ $X2=3.272 $Y2=2.19
r47 9 18 28.2731 $w=5.45e-07 $l=2.88e-07 $layer=POLY_cond $X=3.272 $Y=1.377
+ $X2=3.272 $Y2=1.665
r48 9 10 27.1636 $w=5.45e-07 $l=2.72e-07 $layer=POLY_cond $X=3.272 $Y=1.377
+ $X2=3.272 $Y2=1.105
r49 7 12 76.5092 $w=5e-07 $l=7.15e-07 $layer=POLY_cond $X=3.295 $Y=2.905
+ $X2=3.295 $Y2=2.19
r50 3 10 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.295 $Y=0.765 $X2=3.295
+ $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%A_339_112# 1 2 7 9 13 19 21 23 27 31 34 35
+ 36 39 42 43 44 47 49 52 53 55 57 60 62 66
c167 44 0 1.02982e-20 $X=6.485 $Y=0.35
c168 43 0 7.03008e-20 $X=7.175 $Y=0.35
c169 35 0 1.40543e-20 $X=4.81 $Y=0.35
c170 9 0 8.31313e-20 $X=4.075 $Y=2.905
c171 7 0 1.70715e-19 $X=4.075 $Y=2.185
r172 56 62 56.7131 $w=5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.855 $Y=1.295
+ $X2=4.855 $Y2=0.765
r173 55 58 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=4.815 $Y=1.295
+ $X2=4.815 $Y2=1.33
r174 55 57 6.19221 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=4.815 $Y=1.295
+ $X2=4.815 $Y2=1.195
r175 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.815
+ $Y=1.295 $X2=4.815 $Y2=1.295
r176 50 66 63.6685 $w=5e-07 $l=5.95e-07 $layer=POLY_cond $X=7.315 $Y=1.36
+ $X2=7.315 $Y2=0.765
r177 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.31
+ $Y=1.36 $X2=7.31 $Y2=1.36
r178 47 60 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.31 $Y=1.33
+ $X2=7.31 $Y2=1.195
r179 47 49 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=7.31 $Y=1.33 $X2=7.31
+ $Y2=1.36
r180 45 60 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.26 $Y=0.435
+ $X2=7.26 $Y2=1.195
r181 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.175 $Y=0.35
+ $X2=7.26 $Y2=0.435
r182 43 44 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.175 $Y=0.35
+ $X2=6.485 $Y2=0.35
r183 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.4 $Y=0.435
+ $X2=6.485 $Y2=0.35
r184 41 42 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=6.4 $Y=0.435
+ $X2=6.4 $Y2=1.245
r185 40 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.98 $Y=1.33
+ $X2=4.815 $Y2=1.33
r186 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.315 $Y=1.33
+ $X2=6.4 $Y2=1.245
r187 39 40 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=6.315 $Y=1.33
+ $X2=4.98 $Y2=1.33
r188 37 57 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.895 $Y=0.435
+ $X2=4.895 $Y2=1.195
r189 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.81 $Y=0.35
+ $X2=4.895 $Y2=0.435
r190 35 36 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=4.81 $Y=0.35
+ $X2=3.34 $Y2=0.35
r191 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.255 $Y=0.435
+ $X2=3.34 $Y2=0.35
r192 33 34 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.255 $Y=0.435
+ $X2=3.255 $Y2=1.195
r193 32 53 1.54918 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.94 $Y=1.28
+ $X2=1.845 $Y2=1.28
r194 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.17 $Y=1.28
+ $X2=3.255 $Y2=1.195
r195 31 32 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=3.17 $Y=1.28
+ $X2=1.94 $Y2=1.28
r196 29 53 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=1.365
+ $X2=1.845 $Y2=1.28
r197 29 52 60.4163 $w=1.88e-07 $l=1.035e-06 $layer=LI1_cond $X=1.845 $Y=1.365
+ $X2=1.845 $Y2=2.4
r198 25 53 4.92476 $w=1.8e-07 $l=8.9861e-08 $layer=LI1_cond $X=1.835 $Y=1.195
+ $X2=1.845 $Y2=1.28
r199 25 27 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.835 $Y=1.195
+ $X2=1.835 $Y2=0.77
r200 21 52 6.45386 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=2.525
+ $X2=1.815 $Y2=2.4
r201 21 23 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=1.815 $Y=2.525
+ $X2=1.815 $Y2=2.565
r202 19 50 32.6368 $w=5e-07 $l=3.05e-07 $layer=POLY_cond $X=7.315 $Y=1.665
+ $X2=7.315 $Y2=1.36
r203 19 20 68.7313 $w=5.47e-07 $l=1.03937e-06 $layer=POLY_cond $X=7.315 $Y=1.665
+ $X2=8.095 $Y2=2.27
r204 17 56 37.4521 $w=5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.855 $Y=1.645
+ $X2=4.855 $Y2=1.295
r205 11 20 4.97213 $w=5e-07 $l=2.95e-07 $layer=POLY_cond $X=8.095 $Y=2.565
+ $X2=8.095 $Y2=2.27
r206 11 13 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=8.095 $Y=2.565
+ $X2=8.095 $Y2=2.905
r207 7 17 118.975 $w=3.16e-07 $l=9.04986e-07 $layer=POLY_cond $X=4.075 $Y=2.185
+ $X2=4.855 $Y2=1.915
r208 7 9 77.0442 $w=5e-07 $l=7.2e-07 $layer=POLY_cond $X=4.075 $Y=2.185
+ $X2=4.075 $Y2=2.905
r209 2 23 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.715
+ $Y=2.44 $X2=1.855 $Y2=2.565
r210 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.56 $X2=1.835 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%A_1063_85# 1 2 7 11 13 14 17 23 26 28 32
c61 28 0 2.43525e-20 $X=5.565 $Y=0.765
c62 23 0 1.79686e-19 $X=5.765 $Y=2.355
r63 21 32 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.565 $Y=2.355
+ $X2=5.565 $Y2=2.905
r64 21 28 170.139 $w=5e-07 $l=1.59e-06 $layer=POLY_cond $X=5.565 $Y=2.355
+ $X2=5.565 $Y2=0.765
r65 20 23 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.6 $Y=2.355
+ $X2=5.765 $Y2=2.355
r66 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.6
+ $Y=2.355 $X2=5.6 $Y2=2.355
r67 15 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=2.455
+ $X2=6.83 $Y2=2.37
r68 15 17 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.83 $Y=2.455
+ $X2=6.83 $Y2=2.82
r69 14 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=2.285
+ $X2=6.83 $Y2=2.37
r70 13 25 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.83 $Y=1.325
+ $X2=6.83 $Y2=1.16
r71 13 14 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.83 $Y=1.325
+ $X2=6.83 $Y2=2.285
r72 11 25 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=6.83 $Y=0.7 $X2=6.83
+ $Y2=1.16
r73 7 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=2.37 $X2=6.83
+ $Y2=2.37
r74 7 23 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=6.745 $Y=2.37
+ $X2=5.765 $Y2=2.37
r75 2 17 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=6.69
+ $Y=2.695 $X2=6.83 $Y2=2.82
r76 1 25 182 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_NDIFF $count=1 $X=6.69
+ $Y=0.555 $X2=6.83 $Y2=1.16
r77 1 11 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.69
+ $Y=0.555 $X2=6.83 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%A_865_111# 1 2 8 11 13 16 19 21 27 31
c70 27 0 3.45057e-19 $X=6.44 $Y=0.93
c71 8 0 1.77943e-19 $X=4.385 $Y=1.905
r72 22 31 162.114 $w=5e-07 $l=1.515e-06 $layer=POLY_cond $X=6.44 $Y=1.68
+ $X2=6.44 $Y2=3.195
r73 22 27 80.2544 $w=5e-07 $l=7.5e-07 $layer=POLY_cond $X=6.44 $Y=1.68 $X2=6.44
+ $Y2=0.93
r74 21 24 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.375 $Y=1.68
+ $X2=6.375 $Y2=1.99
r75 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.375
+ $Y=1.68 $X2=6.375 $Y2=1.68
r76 16 18 11.0814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.465 $Y=0.775
+ $X2=4.465 $Y2=1.015
r77 14 19 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.55 $Y=1.99
+ $X2=4.425 $Y2=1.99
r78 13 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.21 $Y=1.99
+ $X2=6.375 $Y2=1.99
r79 13 14 108.299 $w=1.68e-07 $l=1.66e-06 $layer=LI1_cond $X=6.21 $Y=1.99
+ $X2=4.55 $Y2=1.99
r80 9 19 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=2.075
+ $X2=4.425 $Y2=1.99
r81 9 11 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=4.425 $Y=2.075
+ $X2=4.425 $Y2=2.905
r82 8 19 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.385 $Y=1.905
+ $X2=4.425 $Y2=1.99
r83 8 18 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=4.385 $Y=1.905
+ $X2=4.385 $Y2=1.015
r84 2 11 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.325
+ $Y=2.695 $X2=4.465 $Y2=2.905
r85 1 16 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=4.325
+ $Y=0.555 $X2=4.465 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%A_1711_85# 1 2 9 13 17 21 23 27 31 33 34 35
+ 38 42 46 51 52 53
c121 33 0 1.42941e-19 $X=10.76 $Y=1.83
r122 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.34
+ $Y=1.81 $X2=10.34 $Y2=1.81
r123 53 55 8.09337 $w=4.07e-07 $l=2.7e-07 $layer=LI1_cond $X=10.07 $Y=1.74
+ $X2=10.34 $Y2=1.74
r124 52 61 50.2236 $w=5.7e-07 $l=5.25e-07 $layer=POLY_cond $X=8.84 $Y=1.655
+ $X2=8.84 $Y2=2.18
r125 52 60 18.3095 $w=5.7e-07 $l=1.85e-07 $layer=POLY_cond $X=8.84 $Y=1.655
+ $X2=8.84 $Y2=1.47
r126 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.94
+ $Y=1.655 $X2=8.94 $Y2=1.655
r127 46 48 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=10.07 $Y=2.84
+ $X2=10.07 $Y2=3.55
r128 44 53 1.96777 $w=3.3e-07 $l=2.35e-07 $layer=LI1_cond $X=10.07 $Y=1.975
+ $X2=10.07 $Y2=1.74
r129 44 46 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=10.07 $Y=1.975
+ $X2=10.07 $Y2=2.84
r130 40 53 1.96777 $w=3.3e-07 $l=2.35e-07 $layer=LI1_cond $X=10.07 $Y=1.505
+ $X2=10.07 $Y2=1.74
r131 40 42 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=10.07 $Y=1.505
+ $X2=10.07 $Y2=0.7
r132 39 51 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.105 $Y=1.59
+ $X2=8.94 $Y2=1.59
r133 38 53 9.18617 $w=4.07e-07 $l=2.2798e-07 $layer=LI1_cond $X=9.905 $Y=1.59
+ $X2=10.07 $Y2=1.74
r134 38 39 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=9.905 $Y=1.59
+ $X2=9.105 $Y2=1.59
r135 33 56 44.0612 $w=5.1e-07 $l=4.2e-07 $layer=POLY_cond $X=10.76 $Y=1.83
+ $X2=10.34 $Y2=1.83
r136 33 34 23.6275 $w=5.1e-07 $l=2.5e-07 $layer=POLY_cond $X=10.76 $Y=1.83
+ $X2=11.01 $Y2=1.83
r137 29 35 20.7486 $w=5e-07 $l=2.59952e-07 $layer=POLY_cond $X=12.36 $Y=1.575
+ $X2=12.35 $Y2=1.83
r138 29 31 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=12.36 $Y=1.575
+ $X2=12.36 $Y2=1.235
r139 25 35 20.7486 $w=5e-07 $l=2.59952e-07 $layer=POLY_cond $X=12.34 $Y=2.085
+ $X2=12.35 $Y2=1.83
r140 25 27 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=12.34 $Y=2.085
+ $X2=12.34 $Y2=2.59
r141 24 34 23.6275 $w=5.1e-07 $l=2.5e-07 $layer=POLY_cond $X=11.26 $Y=1.83
+ $X2=11.01 $Y2=1.83
r142 23 35 5.02287 $w=5.1e-07 $l=2.6e-07 $layer=POLY_cond $X=12.09 $Y=1.83
+ $X2=12.35 $Y2=1.83
r143 23 24 87.0734 $w=5.1e-07 $l=8.3e-07 $layer=POLY_cond $X=12.09 $Y=1.83
+ $X2=11.26 $Y2=1.83
r144 19 34 24.582 $w=5e-07 $l=2.55e-07 $layer=POLY_cond $X=11.01 $Y=2.085
+ $X2=11.01 $Y2=1.83
r145 19 21 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=11.01 $Y=2.085
+ $X2=11.01 $Y2=2.965
r146 15 34 24.582 $w=5e-07 $l=2.55e-07 $layer=POLY_cond $X=11.01 $Y=1.575
+ $X2=11.01 $Y2=1.83
r147 15 17 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=11.01 $Y=1.575
+ $X2=11.01 $Y2=1.07
r148 13 61 77.5793 $w=5e-07 $l=7.25e-07 $layer=POLY_cond $X=8.805 $Y=2.905
+ $X2=8.805 $Y2=2.18
r149 9 60 75.4392 $w=5e-07 $l=7.05e-07 $layer=POLY_cond $X=8.805 $Y=0.765
+ $X2=8.805 $Y2=1.47
r150 2 48 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=9.93
+ $Y=2.695 $X2=10.07 $Y2=3.55
r151 2 46 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.93
+ $Y=2.695 $X2=10.07 $Y2=2.84
r152 1 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.93
+ $Y=0.555 $X2=10.07 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%A_1494_539# 1 2 9 13 17 22 25 26 28 29 30
+ 33 34 37 38 39
c99 33 0 1.42941e-19 $X=9.56 $Y=2.005
r100 38 39 108.299 $w=1.68e-07 $l=1.66e-06 $layer=LI1_cond $X=7.71 $Y=2.675
+ $X2=7.71 $Y2=1.015
r101 37 38 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.62 $Y=2.84
+ $X2=7.62 $Y2=2.675
r102 34 42 54.626 $w=5.55e-07 $l=5.6e-07 $layer=POLY_cond $X=9.652 $Y=2.005
+ $X2=9.652 $Y2=2.565
r103 34 41 18.4754 $w=5.55e-07 $l=1.85e-07 $layer=POLY_cond $X=9.652 $Y=2.005
+ $X2=9.652 $Y2=1.82
r104 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.56
+ $Y=2.005 $X2=9.56 $Y2=2.005
r105 31 33 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=9.56 $Y=2.325
+ $X2=9.56 $Y2=2.005
r106 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.395 $Y=2.41
+ $X2=9.56 $Y2=2.325
r107 29 30 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=9.395 $Y=2.41
+ $X2=8.595 $Y2=2.41
r108 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.51 $Y=2.325
+ $X2=8.595 $Y2=2.41
r109 27 28 106.995 $w=1.68e-07 $l=1.64e-06 $layer=LI1_cond $X=8.51 $Y=0.685
+ $X2=8.51 $Y2=2.325
r110 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.425 $Y=0.6
+ $X2=8.51 $Y2=0.685
r111 25 26 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=8.425 $Y=0.6
+ $X2=7.795 $Y2=0.6
r112 20 39 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=7.667 $Y=0.888
+ $X2=7.667 $Y2=1.015
r113 20 22 5.55884 $w=2.53e-07 $l=1.23e-07 $layer=LI1_cond $X=7.667 $Y=0.888
+ $X2=7.667 $Y2=0.765
r114 19 26 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=7.667 $Y=0.685
+ $X2=7.795 $Y2=0.6
r115 19 22 3.61551 $w=2.53e-07 $l=8e-08 $layer=LI1_cond $X=7.667 $Y=0.685
+ $X2=7.667 $Y2=0.765
r116 15 37 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=7.62 $Y=2.85
+ $X2=7.62 $Y2=2.84
r117 15 17 17.122 $w=3.48e-07 $l=5.2e-07 $layer=LI1_cond $X=7.62 $Y=2.85
+ $X2=7.62 $Y2=3.37
r118 13 42 67.4137 $w=5e-07 $l=6.3e-07 $layer=POLY_cond $X=9.68 $Y=3.195
+ $X2=9.68 $Y2=2.565
r119 9 41 95.2352 $w=5e-07 $l=8.9e-07 $layer=POLY_cond $X=9.68 $Y=0.93 $X2=9.68
+ $Y2=1.82
r120 2 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.47
+ $Y=2.695 $X2=7.61 $Y2=2.84
r121 2 17 600 $w=1.7e-07 $l=7.41704e-07 $layer=licon1_PDIFF $count=1 $X=7.47
+ $Y=2.695 $X2=7.61 $Y2=3.37
r122 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.565
+ $Y=0.555 $X2=7.705 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%A_2365_443# 1 2 9 13 17 21 27 28 30 31
r49 28 34 25.2235 $w=5.55e-07 $l=2.55e-07 $layer=POLY_cond $X=13.227 $Y=1.83
+ $X2=13.227 $Y2=2.085
r50 28 33 25.2235 $w=5.55e-07 $l=2.55e-07 $layer=POLY_cond $X=13.227 $Y=1.83
+ $X2=13.227 $Y2=1.575
r51 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.135
+ $Y=1.83 $X2=13.135 $Y2=1.83
r52 25 31 1.23199 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=12.135 $Y=1.83
+ $X2=11.97 $Y2=1.83
r53 25 27 34.9225 $w=3.28e-07 $l=1e-06 $layer=LI1_cond $X=12.135 $Y=1.83
+ $X2=13.135 $Y2=1.83
r54 23 31 5.29963 $w=3.2e-07 $l=1.69926e-07 $layer=LI1_cond $X=11.96 $Y=1.995
+ $X2=11.97 $Y2=1.83
r55 23 30 7.43512 $w=3.08e-07 $l=2e-07 $layer=LI1_cond $X=11.96 $Y=1.995
+ $X2=11.96 $Y2=2.195
r56 19 31 5.29963 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=11.97 $Y=1.665
+ $X2=11.97 $Y2=1.83
r57 19 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.97 $Y=1.665
+ $X2=11.97 $Y2=1.235
r58 17 30 5.81909 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.95 $Y=2.36
+ $X2=11.95 $Y2=2.195
r59 13 33 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=13.255 $Y=1.07
+ $X2=13.255 $Y2=1.575
r60 9 34 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=13.235 $Y=2.965
+ $X2=13.235 $Y2=2.085
r61 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=11.825
+ $Y=2.215 $X2=11.95 $Y2=2.36
r62 1 21 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=11.845
+ $Y=1.025 $X2=11.97 $Y2=1.235
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%VPWR 1 2 3 4 5 6 19 22 29 42 46 57 65 73
r98 71 73 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=12.41 $Y=3.63
+ $X2=13.13 $Y2=3.63
r99 70 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.13 $Y=3.59
+ $X2=13.13 $Y2=3.59
r100 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.41 $Y=3.59
+ $X2=12.41 $Y2=3.59
r101 68 70 5.32947 $w=9.48e-07 $l=4.15e-07 $layer=LI1_cond $X=12.77 $Y=3.175
+ $X2=12.77 $Y2=3.59
r102 65 68 10.7232 $w=9.48e-07 $l=8.35e-07 $layer=LI1_cond $X=12.77 $Y=2.34
+ $X2=12.77 $Y2=3.175
r103 62 71 0.343595 $w=3.7e-07 $l=8.95e-07 $layer=MET1_cond $X=11.515 $Y=3.63
+ $X2=12.41 $Y2=3.63
r104 60 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.515 $Y=3.59
+ $X2=11.515 $Y2=3.59
r105 57 60 27.0515 $w=5.33e-07 $l=1.21e-06 $layer=LI1_cond $X=11.337 $Y=2.36
+ $X2=11.337 $Y2=3.57
r106 54 62 0.834994 $w=3.7e-07 $l=2.175e-06 $layer=MET1_cond $X=9.34 $Y=3.63
+ $X2=11.515 $Y2=3.63
r107 52 54 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.62 $Y=3.63
+ $X2=9.34 $Y2=3.63
r108 51 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.34 $Y=3.6
+ $X2=9.34 $Y2=3.6
r109 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.62 $Y=3.6
+ $X2=8.62 $Y2=3.6
r110 49 51 5.20105 $w=9.48e-07 $l=4.05e-07 $layer=LI1_cond $X=8.98 $Y=3.195
+ $X2=8.98 $Y2=3.6
r111 46 49 4.55895 $w=9.48e-07 $l=3.55e-07 $layer=LI1_cond $X=8.98 $Y=2.84
+ $X2=8.98 $Y2=3.195
r112 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.1 $Y=3.59
+ $X2=6.1 $Y2=3.59
r113 40 42 0.819232 $w=7.28e-07 $l=5e-08 $layer=LI1_cond $X=6.05 $Y=3.35 $X2=6.1
+ $Y2=3.35
r114 37 43 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.38 $Y=3.63
+ $X2=6.1 $Y2=3.63
r115 36 40 10.9777 $w=7.28e-07 $l=6.7e-07 $layer=LI1_cond $X=5.38 $Y=3.35
+ $X2=6.05 $Y2=3.35
r116 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.38 $Y=3.59
+ $X2=5.38 $Y2=3.59
r117 33 37 0.946327 $w=3.7e-07 $l=2.465e-06 $layer=MET1_cond $X=2.915 $Y=3.63
+ $X2=5.38 $Y2=3.63
r118 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.915 $Y=3.59
+ $X2=2.915 $Y2=3.59
r119 29 32 15.4587 $w=5.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2.735 $Y=2.905
+ $X2=2.735 $Y2=3.59
r120 26 33 0.717903 $w=3.7e-07 $l=1.87e-06 $layer=MET1_cond $X=1.045 $Y=3.63
+ $X2=2.915 $Y2=3.63
r121 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.045 $Y=3.59
+ $X2=1.045 $Y2=3.59
r122 22 25 20.7793 $w=5.88e-07 $l=1.025e-06 $layer=LI1_cond $X=0.865 $Y=2.565
+ $X2=0.865 $Y2=3.59
r123 19 52 0.637283 $w=3.7e-07 $l=1.66e-06 $layer=MET1_cond $X=6.96 $Y=3.63
+ $X2=8.62 $Y2=3.63
r124 19 43 0.330159 $w=3.7e-07 $l=8.6e-07 $layer=MET1_cond $X=6.96 $Y=3.63
+ $X2=6.1 $Y2=3.63
r125 6 68 300 $w=1.7e-07 $l=1.08e-06 $layer=licon1_PDIFF $count=2 $X=12.59
+ $Y=2.215 $X2=12.845 $Y2=3.175
r126 6 65 300 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=2 $X=12.59
+ $Y=2.215 $X2=12.845 $Y2=2.34
r127 5 60 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=11.26
+ $Y=2.215 $X2=11.4 $Y2=3.57
r128 5 57 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=11.26
+ $Y=2.215 $X2=11.4 $Y2=2.36
r129 4 49 300 $w=1.7e-07 $l=6.06218e-07 $layer=licon1_PDIFF $count=2 $X=9.055
+ $Y=2.695 $X2=9.29 $Y2=3.195
r130 4 46 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=9.055
+ $Y=2.695 $X2=9.29 $Y2=2.84
r131 3 40 300 $w=1.7e-07 $l=4.78278e-07 $layer=licon1_PDIFF $count=2 $X=5.815
+ $Y=2.695 $X2=6.05 $Y2=3.07
r132 2 29 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=2.695 $X2=2.905 $Y2=2.905
r133 1 22 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.935
+ $Y=2.44 $X2=1.075 $Y2=2.565
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%A_709_111# 1 2 9 11 14 17
r31 16 17 112.214 $w=1.68e-07 $l=1.72e-06 $layer=LI1_cond $X=3.615 $Y=0.935
+ $X2=3.615 $Y2=2.655
r32 14 16 8.28756 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.685 $Y=0.775
+ $X2=3.685 $Y2=0.935
r33 9 17 6.75802 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=3.65 $Y=2.775
+ $X2=3.65 $Y2=2.655
r34 9 11 6.2424 $w=2.38e-07 $l=1.3e-07 $layer=LI1_cond $X=3.65 $Y=2.775 $X2=3.65
+ $Y2=2.905
r35 2 11 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.545
+ $Y=2.695 $X2=3.685 $Y2=2.905
r36 1 14 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=3.545
+ $Y=0.555 $X2=3.685 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%Q 1 2 7 8 9 10 11 12 13 25 46 50 54
r31 50 51 7.61291 $w=4.33e-07 $l=1.65e-07 $layer=LI1_cond $X=10.672 $Y=2.36
+ $X2=10.672 $Y2=2.195
r32 36 54 0.185451 $w=4.33e-07 $l=7e-09 $layer=LI1_cond $X=10.672 $Y=2.412
+ $X2=10.672 $Y2=2.405
r33 23 46 1.24517 $w=4.33e-07 $l=4.7e-08 $layer=LI1_cond $X=10.672 $Y=1.248
+ $X2=10.672 $Y2=1.295
r34 13 43 11.2595 $w=4.33e-07 $l=4.25e-07 $layer=LI1_cond $X=10.672 $Y=3.145
+ $X2=10.672 $Y2=3.57
r35 12 13 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=10.672 $Y=2.775
+ $X2=10.672 $Y2=3.145
r36 11 54 1.03322 $w=4.33e-07 $l=3.9e-08 $layer=LI1_cond $X=10.672 $Y=2.366
+ $X2=10.672 $Y2=2.405
r37 11 50 0.158958 $w=4.33e-07 $l=6e-09 $layer=LI1_cond $X=10.672 $Y=2.366
+ $X2=10.672 $Y2=2.36
r38 11 12 8.58371 $w=4.33e-07 $l=3.24e-07 $layer=LI1_cond $X=10.672 $Y=2.451
+ $X2=10.672 $Y2=2.775
r39 11 36 1.03322 $w=4.33e-07 $l=3.9e-08 $layer=LI1_cond $X=10.672 $Y=2.451
+ $X2=10.672 $Y2=2.412
r40 10 51 8.65632 $w=2.03e-07 $l=1.6e-07 $layer=LI1_cond $X=10.787 $Y=2.035
+ $X2=10.787 $Y2=2.195
r41 9 10 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=10.787 $Y=1.665
+ $X2=10.787 $Y2=2.035
r42 9 48 10.8204 $w=2.03e-07 $l=2e-07 $layer=LI1_cond $X=10.787 $Y=1.665
+ $X2=10.787 $Y2=1.465
r43 8 48 7.24201 $w=4.33e-07 $l=1.51e-07 $layer=LI1_cond $X=10.672 $Y=1.314
+ $X2=10.672 $Y2=1.465
r44 8 46 0.503366 $w=4.33e-07 $l=1.9e-08 $layer=LI1_cond $X=10.672 $Y=1.314
+ $X2=10.672 $Y2=1.295
r45 8 23 0.503366 $w=4.33e-07 $l=1.9e-08 $layer=LI1_cond $X=10.672 $Y=1.229
+ $X2=10.672 $Y2=1.248
r46 7 8 8.05385 $w=4.33e-07 $l=3.04e-07 $layer=LI1_cond $X=10.672 $Y=0.925
+ $X2=10.672 $Y2=1.229
r47 7 25 2.2519 $w=4.33e-07 $l=8.5e-08 $layer=LI1_cond $X=10.672 $Y=0.925
+ $X2=10.672 $Y2=0.84
r48 2 50 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=10.495
+ $Y=2.215 $X2=10.62 $Y2=2.36
r49 2 43 300 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_PDIFF $count=2 $X=10.495
+ $Y=2.215 $X2=10.62 $Y2=3.57
r50 1 25 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=10.495
+ $Y=0.695 $X2=10.62 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%Q_N 1 2 7 8 9 10 11 12 13 35
r16 33 35 1.81098 $w=3.48e-07 $l=5.5e-08 $layer=LI1_cond $X=13.635 $Y=2.35
+ $X2=13.635 $Y2=2.405
r17 13 42 14.6525 $w=3.48e-07 $l=4.45e-07 $layer=LI1_cond $X=13.635 $Y=3.145
+ $X2=13.635 $Y2=3.59
r18 12 13 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=13.635 $Y=2.775
+ $X2=13.635 $Y2=3.145
r19 11 33 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=13.635 $Y=2.335
+ $X2=13.635 $Y2=2.35
r20 11 45 5.31946 $w=3.48e-07 $l=1.6e-07 $layer=LI1_cond $X=13.635 $Y=2.335
+ $X2=13.635 $Y2=2.175
r21 11 12 11.6891 $w=3.48e-07 $l=3.55e-07 $layer=LI1_cond $X=13.635 $Y=2.42
+ $X2=13.635 $Y2=2.775
r22 11 35 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=13.635 $Y=2.42
+ $X2=13.635 $Y2=2.405
r23 10 45 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=13.645 $Y=2.035
+ $X2=13.645 $Y2=2.175
r24 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.645 $Y=1.665
+ $X2=13.645 $Y2=2.035
r25 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.645 $Y=1.295
+ $X2=13.645 $Y2=1.665
r26 7 8 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=13.645 $Y=0.84
+ $X2=13.645 $Y2=1.295
r27 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=13.485
+ $Y=2.215 $X2=13.625 $Y2=2.34
r28 2 42 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=13.485
+ $Y=2.215 $X2=13.625 $Y2=3.59
r29 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.505
+ $Y=0.695 $X2=13.645 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXBP_1%VGND 1 2 3 4 5 6 19 22 31 47 50 61 68 72
r101 74 76 6.42105 $w=9.48e-07 $l=5e-07 $layer=LI1_cond $X=12.79 $Y=0.82
+ $X2=12.79 $Y2=1.32
r102 69 72 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=12.43 $Y=0.44
+ $X2=13.15 $Y2=0.44
r103 68 74 4.36632 $w=9.48e-07 $l=3.4e-07 $layer=LI1_cond $X=12.79 $Y=0.48
+ $X2=12.79 $Y2=0.82
r104 68 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.15 $Y=0.48
+ $X2=13.15 $Y2=0.48
r105 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.43 $Y=0.48
+ $X2=12.43 $Y2=0.48
r106 62 69 0.347434 $w=3.7e-07 $l=9.05e-07 $layer=MET1_cond $X=11.525 $Y=0.44
+ $X2=12.43 $Y2=0.44
r107 61 65 7.32733 $w=5.53e-07 $l=3.4e-07 $layer=LI1_cond $X=11.347 $Y=0.48
+ $X2=11.347 $Y2=0.82
r108 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.525 $Y=0.48
+ $X2=11.525 $Y2=0.48
r109 56 58 5.90737 $w=9.48e-07 $l=4.6e-07 $layer=LI1_cond $X=9.25 $Y=0.7
+ $X2=9.25 $Y2=1.16
r110 54 62 0.735179 $w=3.7e-07 $l=1.915e-06 $layer=MET1_cond $X=9.61 $Y=0.44
+ $X2=11.525 $Y2=0.44
r111 51 54 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.89 $Y=0.44
+ $X2=9.61 $Y2=0.44
r112 50 56 2.82526 $w=9.48e-07 $l=2.2e-07 $layer=LI1_cond $X=9.25 $Y=0.48
+ $X2=9.25 $Y2=0.7
r113 50 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.61 $Y=0.48
+ $X2=9.61 $Y2=0.48
r114 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.89 $Y=0.48
+ $X2=8.89 $Y2=0.48
r115 44 47 0.512605 $w=6.98e-07 $l=3e-08 $layer=LI1_cond $X=6.02 $Y=0.715
+ $X2=6.05 $Y2=0.715
r116 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.02 $Y=0.48
+ $X2=6.02 $Y2=0.48
r117 41 45 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.3 $Y=0.44
+ $X2=6.02 $Y2=0.44
r118 40 44 12.3025 $w=6.98e-07 $l=7.2e-07 $layer=LI1_cond $X=5.3 $Y=0.715
+ $X2=6.02 $Y2=0.715
r119 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.3 $Y=0.48
+ $X2=5.3 $Y2=0.48
r120 35 41 0.919453 $w=3.7e-07 $l=2.395e-06 $layer=MET1_cond $X=2.905 $Y=0.44
+ $X2=5.3 $Y2=0.44
r121 32 35 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.185 $Y=0.44
+ $X2=2.905 $Y2=0.44
r122 31 37 3.90674 $w=8.88e-07 $l=2.85e-07 $layer=LI1_cond $X=2.545 $Y=0.48
+ $X2=2.545 $Y2=0.765
r123 31 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.905 $Y=0.48
+ $X2=2.905 $Y2=0.48
r124 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.185 $Y=0.48
+ $X2=2.185 $Y2=0.48
r125 26 32 0.280251 $w=3.7e-07 $l=7.3e-07 $layer=MET1_cond $X=1.455 $Y=0.44
+ $X2=2.185 $Y2=0.44
r126 23 26 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.735 $Y=0.44
+ $X2=1.455 $Y2=0.44
r127 22 28 3.72421 $w=9.48e-07 $l=2.9e-07 $layer=LI1_cond $X=1.095 $Y=0.48
+ $X2=1.095 $Y2=0.77
r128 22 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.455 $Y=0.48
+ $X2=1.455 $Y2=0.48
r129 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.735 $Y=0.48
+ $X2=0.735 $Y2=0.48
r130 19 51 0.740937 $w=3.7e-07 $l=1.93e-06 $layer=MET1_cond $X=6.96 $Y=0.44
+ $X2=8.89 $Y2=0.44
r131 19 45 0.360871 $w=3.7e-07 $l=9.4e-07 $layer=MET1_cond $X=6.96 $Y=0.44
+ $X2=6.02 $Y2=0.44
r132 6 76 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=12.61
+ $Y=1.025 $X2=12.865 $Y2=1.32
r133 6 74 182 $w=1.7e-07 $l=3.42491e-07 $layer=licon1_NDIFF $count=1 $X=12.61
+ $Y=1.025 $X2=12.865 $Y2=0.82
r134 5 65 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=11.26
+ $Y=0.695 $X2=11.4 $Y2=0.82
r135 4 58 182 $w=1.7e-07 $l=7.12881e-07 $layer=licon1_NDIFF $count=1 $X=9.055
+ $Y=0.555 $X2=9.29 $Y2=1.16
r136 4 56 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=9.055
+ $Y=0.555 $X2=9.29 $Y2=0.7
r137 3 47 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=5.815
+ $Y=0.555 $X2=6.05 $Y2=0.8
r138 2 37 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.68
+ $Y=0.555 $X2=2.825 $Y2=0.765
r139 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.915
+ $Y=0.56 $X2=1.055 $Y2=0.77
.ends

