* File: sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3.spice
* Created: Fri Aug 28 09:37:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3.pex.spice"
.subckt sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3  VNB VPB LVPWR VGND SLEEP_B A
+ X VPWR
* 
* VPWR	VPWR
* X	X
* A	A
* SLEEP_B	SLEEP_B
* VGND	VGND
* LVPWR	LVPWR
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_A_3617_1198#_M1018_g N_A_528_1171#_M1018_s N_VNB_M1018_b
+ NSHORT L=0.15 W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_528_1171#_M1007_g N_A_1472_1171#_M1007_s N_VNB_M1018_b
+ NSHORT L=0.15 W=0.74 AD=0.2331 AS=0.1184 PD=2.11 PS=1.06 NRD=4.86 NRS=6.48 M=1
+ R=4.93333 SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_A_3617_1198#_M1019_g N_A_528_1171#_M1018_s N_VNB_M1018_b
+ NSHORT L=0.15 W=0.74 AD=0.1221 AS=0.1036 PD=1.07 PS=1.02 NRD=8.1 NRS=0 M=1
+ R=4.93333 SA=75000.6 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_528_1171#_M1009_g N_A_1472_1171#_M1007_s N_VNB_M1018_b
+ NSHORT L=0.15 W=0.74 AD=0.1221 AS=0.1184 PD=1.07 PS=1.06 NRD=0 NRS=0 M=1
+ R=4.93333 SA=75000.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1019_d N_A_3617_1198#_M1027_g N_A_528_1171#_M1027_s N_VNB_M1018_b
+ NSHORT L=0.15 W=0.74 AD=0.1221 AS=0.1184 PD=1.07 PS=1.06 NRD=0 NRS=0 M=1
+ R=4.93333 SA=75001.1 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1009_d N_A_528_1171#_M1014_g N_A_1472_1171#_M1014_s N_VNB_M1018_b
+ NSHORT L=0.15 W=0.74 AD=0.1221 AS=0.1036 PD=1.07 PS=1.02 NRD=8.1 NRS=0 M=1
+ R=4.93333 SA=75001.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1033 N_VGND_M1033_d N_A_3617_1198#_M1033_g N_A_528_1171#_M1027_s N_VNB_M1018_b
+ NSHORT L=0.15 W=0.74 AD=0.2331 AS=0.1184 PD=2.11 PS=1.06 NRD=4.86 NRS=6.48 M=1
+ R=4.93333 SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_A_528_1171#_M1016_g N_A_1472_1171#_M1014_s N_VNB_M1018_b
+ NSHORT L=0.15 W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1
+ R=4.93333 SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1024_d N_A_M1024_g N_A_3617_1198#_M1024_s N_VNB_M1018_b NSHORT
+ L=0.15 W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1046 N_VGND_M1046_d N_A_M1046_g N_A_3617_1198#_M1024_s N_VNB_M1018_b NSHORT
+ L=0.15 W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_262_107#_M1008_g N_X_M1008_s N_VNB_M1018_b NHV L=0.5
+ W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=2 SA=250000 SB=250002
+ A=0.5 P=3 MULT=1
MM1000 N_A_362_1243#_M1000_d N_VGND_M1000_g N_VGND_M1000_s N_VNB_M1018_b NHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1030 N_VGND_M1008_d N_A_262_107#_M1030_g N_X_M1030_s N_VNB_M1018_b NHV L=0.5
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=2 SA=250001 SB=250001
+ A=0.5 P=3 MULT=1
MM1047 N_VGND_M1047_d N_A_262_107#_M1047_g N_X_M1030_s N_VNB_M1018_b NHV L=0.5
+ W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=2 SA=250002 SB=250000
+ A=0.5 P=3 MULT=1
MM1012 N_VGND_M1012_d N_A_840_107#_M1012_g N_A_262_107#_M1012_s N_VNB_M1018_b
+ NHV L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=2 SA=250000
+ SB=250001 A=0.5 P=3 MULT=1
MM1034 N_VGND_M1012_d N_A_840_107#_M1034_g N_A_262_107#_M1034_s N_VNB_M1018_b
+ NHV L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=2 SA=250001
+ SB=250000 A=0.5 P=3 MULT=1
MM1002 N_VGND_M1002_d N_A_2092_381#_M1002_g N_A_840_107#_M1002_s N_VNB_M1018_b
+ NHV L=0.5 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1045 N_VGND_M1045_d N_SLEEP_B_M1045_g N_A_2092_381#_M1045_s N_VNB_M1018_b NHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1004 N_VGND_M1004_d N_A_528_1171#_M1004_g N_A_362_1243#_M1004_s N_VNB_M1018_b
+ NHVNATIVE L=0.9 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=1.11111
+ SA=450000 SB=450008 A=0.9 P=3.8 MULT=1
MM1010 N_VGND_M1010_d N_A_528_1171#_M1010_g N_A_362_1243#_M1004_s N_VNB_M1018_b
+ NHVNATIVE L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=1.11111
+ SA=450001 SB=450007 A=0.9 P=3.8 MULT=1
MM1023 N_VGND_M1010_d N_A_528_1171#_M1023_g N_A_362_1243#_M1023_s N_VNB_M1018_b
+ NHVNATIVE L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=1.11111
+ SA=450002 SB=450006 A=0.9 P=3.8 MULT=1
MM1040 N_VGND_M1040_d N_A_528_1171#_M1040_g N_A_362_1243#_M1023_s N_VNB_M1018_b
+ NHVNATIVE L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=1.11111
+ SA=450003 SB=450005 A=0.9 P=3.8 MULT=1
MM1001 N_VGND_M1040_d N_A_1472_1171#_M1001_g N_A_840_107#_M1001_s N_VNB_M1018_b
+ NHVNATIVE L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=1.11111
+ SA=450005 SB=450003 A=0.9 P=3.8 MULT=1
MM1029 N_VGND_M1029_d N_A_1472_1171#_M1029_g N_A_840_107#_M1001_s N_VNB_M1018_b
+ NHVNATIVE L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=1.11111
+ SA=450006 SB=450002 A=0.9 P=3.8 MULT=1
MM1032 N_VGND_M1029_d N_A_1472_1171#_M1032_g N_A_840_107#_M1032_s N_VNB_M1018_b
+ NHVNATIVE L=0.9 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=1.11111
+ SA=450007 SB=450001 A=0.9 P=3.8 MULT=1
MM1041 N_VGND_M1041_d N_A_1472_1171#_M1041_g N_A_840_107#_M1032_s N_VNB_M1018_b
+ NHVNATIVE L=0.9 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=1.11111
+ SA=450008 SB=450000 A=0.9 P=3.8 MULT=1
MM1006 N_A_528_1171#_M1006_d N_A_3617_1198#_M1006_g N_LVPWR_M1006_s
+ N_LVPWR_M1006_b PHIGHVT L=0.15 W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83
+ NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.2 SB=75001.6 A=0.168 P=2.54
+ MULT=1
MM1003 N_A_1472_1171#_M1003_d N_A_528_1171#_M1003_g N_LVPWR_M1003_s
+ N_LVPWR_M1006_b PHIGHVT L=0.15 W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83
+ NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.2 SB=75001.6 A=0.168 P=2.54
+ MULT=1
MM1013 N_A_528_1171#_M1006_d N_A_3617_1198#_M1013_g N_LVPWR_M1013_s
+ N_LVPWR_M1006_b PHIGHVT L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42
+ NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.7 SB=75001.1 A=0.168 P=2.54
+ MULT=1
MM1026 N_A_1472_1171#_M1003_d N_A_528_1171#_M1026_g N_LVPWR_M1026_s
+ N_LVPWR_M1006_b PHIGHVT L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42
+ NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.7 SB=75001.1 A=0.168 P=2.54
+ MULT=1
MM1015 N_A_528_1171#_M1015_d N_A_3617_1198#_M1015_g N_LVPWR_M1013_s
+ N_LVPWR_M1006_b PHIGHVT L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42
+ NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.1 SB=75000.7 A=0.168 P=2.54
+ MULT=1
MM1035 N_A_1472_1171#_M1035_d N_A_528_1171#_M1035_g N_LVPWR_M1026_s
+ N_LVPWR_M1006_b PHIGHVT L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42
+ NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.1 SB=75000.7 A=0.168 P=2.54
+ MULT=1
MM1025 N_A_528_1171#_M1015_d N_A_3617_1198#_M1025_g N_LVPWR_M1025_s
+ N_LVPWR_M1006_b PHIGHVT L=0.15 W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83
+ NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.6 SB=75000.2 A=0.168 P=2.54
+ MULT=1
MM1038 N_A_1472_1171#_M1035_d N_A_528_1171#_M1038_g N_LVPWR_M1038_s
+ N_LVPWR_M1006_b PHIGHVT L=0.15 W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83
+ NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.6 SB=75000.2 A=0.168 P=2.54
+ MULT=1
MM1031 N_A_3617_1198#_M1031_d N_A_M1031_g N_LVPWR_M1031_s N_LVPWR_M1006_b
+ PHIGHVT L=0.15 W=1.12 AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533
+ M=1 R=7.46667 SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1044 N_A_3617_1198#_M1031_d N_A_M1044_g N_LVPWR_M1044_s N_LVPWR_M1006_b
+ PHIGHVT L=0.15 W=1.12 AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533
+ M=1 R=7.46667 SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_A_262_107#_M1005_g N_X_M1005_s N_VPB_M1005_b PHV L=0.5
+ W=3 AD=0.42 AS=0.795 PD=3.28 PS=6.53 NRD=0 NRS=0 M=1 R=6 SA=250000 SB=250002
+ A=1.5 P=7 MULT=1
MM1011 N_VPWR_M1005_d N_A_262_107#_M1011_g N_X_M1011_s N_VPB_M1005_b PHV L=0.5
+ W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 M=1 R=6 SA=250001 SB=250001
+ A=1.5 P=7 MULT=1
MM1036 N_VPWR_M1036_d N_A_262_107#_M1036_g N_X_M1011_s N_VPB_M1005_b PHV L=0.5
+ W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=6 SA=250002 SB=250000
+ A=1.5 P=7 MULT=1
MM39_noxref N_VPWR_M39_noxref_d N_A_840_107#_M39_noxref_g
+ N_A_262_107#_M39_noxref_s N_VPB_M1005_b PHV L=0.5 W=1.5 AD=0.21 AS=0.3975
+ PD=1.78 PS=3.53 NRD=0 NRS=0 M=1 R=3 SA=250000 SB=250001 A=0.75 P=4 MULT=1
MM40_noxref N_A_262_107#_M40_noxref_d N_A_840_107#_M40_noxref_g
+ N_VPWR_M39_noxref_d N_VPB_M1005_b PHV L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53
+ PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001 SB=250000 A=0.75 P=4 MULT=1
MM1022 N_A_1410_571#_M1022_d N_A_840_107#_M1022_g N_A_362_1243#_M1022_s
+ N_VPB_M1005_b PHV L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0
+ M=1 R=3 SA=250000 SB=250001 A=0.75 P=4 MULT=1
MM1043 N_A_840_107#_M1043_d N_A_362_1243#_M1043_g N_A_1410_571#_M1022_d
+ N_VPB_M1005_b PHV L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0
+ M=1 R=3 SA=250001 SB=250000 A=0.75 P=4 MULT=1
MM43_noxref N_A_1410_571#_M43_noxref_d N_A_2092_381#_M43_noxref_g
+ N_VPWR_M43_noxref_s N_VPB_M1005_b PHV L=0.5 W=3 AD=0.42 AS=0.795 PD=3.28
+ PS=6.53 NRD=0 NRS=0 M=1 R=6 SA=250000 SB=250002 A=1.5 P=7 MULT=1
MM44_noxref N_VPWR_M44_noxref_d N_A_2092_381#_M44_noxref_g
+ N_A_1410_571#_M43_noxref_d N_VPB_M1005_b PHV L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28
+ PS=3.28 NRD=0 NRS=0 M=1 R=6 SA=250001 SB=250002 A=1.5 P=7 MULT=1
MM45_noxref N_A_1410_571#_M45_noxref_d N_A_2092_381#_M45_noxref_g
+ N_VPWR_M44_noxref_d N_VPB_M1005_b PHV L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28
+ PS=3.28 NRD=0 NRS=0 M=1 R=6 SA=250002 SB=250001 A=1.5 P=7 MULT=1
MM46_noxref N_VPWR_M46_noxref_d N_A_2092_381#_M46_noxref_g
+ N_A_1410_571#_M45_noxref_d N_VPB_M1005_b PHV L=0.5 W=3 AD=0.795 AS=0.42
+ PD=6.53 PS=3.28 NRD=0 NRS=0 M=1 R=6 SA=250002 SB=250000 A=1.5 P=7 MULT=1
MM1020 N_VPWR_M1020_d N_SLEEP_B_M1020_g N_A_2092_381#_M1020_s N_VPB_M1005_b PHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
DX48_noxref N_VNB_M1018_b N_VPB_M1005_b NWDIODE A=60.4821 P=40.97
DX49_noxref N_VNB_M1018_b N_LVPWR_M1006_b NWDIODE A=17.415 P=16.7
*
.include "sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3.pxi.spice"
*
.ends
*
*
