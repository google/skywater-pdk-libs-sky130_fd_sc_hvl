* File: sky130_fd_sc_hvl__sdlxtp_1.spice
* Created: Wed Sep  2 09:10:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__sdlxtp_1.pex.spice"
.subckt sky130_fd_sc_hvl__sdlxtp_1  VNB VPB SCE D SCD GATE VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE	GATE
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_SCE_M1004_g N_A_30_587#_M1004_s N_VNB_M1004_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250004 A=0.21 P=1.84 MULT=1
MM1015 A_347_107# N_D_M1015_g N_VGND_M1004_d N_VNB_M1004_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84 SA=250001
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1016 N_A_489_107#_M1016_d N_A_30_587#_M1016_g A_347_107# N_VNB_M1004_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1008 A_645_107# N_SCE_M1008_g N_A_489_107#_M1016_d N_VNB_M1004_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1009 N_VGND_M1009_d N_SCD_M1009_g A_645_107# N_VNB_M1004_b NHV L=0.5 W=0.42
+ AD=0.05985 AS=0.0441 PD=0.705 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250003
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1006 N_A_944_107#_M1006_d N_GATE_M1006_g N_VGND_M1009_d N_VNB_M1004_b NHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.05985 PD=1.37 PS=0.705 NRD=0 NRS=1.3566 M=1 R=0.84
+ SA=250004 SB=250000 A=0.21 P=1.84 MULT=1
MM1005 N_A_1214_107#_M1005_d N_A_944_107#_M1005_g N_VGND_M1005_s N_VNB_M1004_b
+ NHV L=0.5 W=0.42 AD=0.1113 AS=0.1197 PD=1.37 PS=1.41 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1002 N_A_1480_107#_M1002_d N_A_1214_107#_M1002_g N_A_489_107#_M1002_s
+ N_VNB_M1004_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1019 A_1636_107# N_A_944_107#_M1019_g N_A_1480_107#_M1002_d N_VNB_M1004_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1022 N_VGND_M1022_d N_A_1678_81#_M1022_g A_1636_107# N_VNB_M1004_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1013 N_VGND_M1013_d N_A_1480_107#_M1013_g N_A_1678_81#_M1013_s N_VNB_M1004_b
+ NHV L=0.5 W=0.42 AD=0.0879308 AS=0.1113 PD=0.807692 PS=1.37 NRD=25.7754 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1020 N_Q_M1020_d N_A_1480_107#_M1020_g N_VGND_M1013_d N_VNB_M1004_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.157019 PD=2.03 PS=1.44231 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1018 N_VPWR_M1018_d N_SCE_M1018_g N_A_30_587#_M1018_s N_VPB_M1018_b PHV L=0.5
+ W=0.42 AD=0.0879308 AS=0.1197 PD=0.807692 PS=1.41 NRD=43.1851 NRS=0 M=1 R=0.84
+ SA=250000 SB=250004 A=0.21 P=1.84 MULT=1
MM1010 A_362_587# N_SCE_M1010_g N_VPWR_M1018_d N_VPB_M1018_b PHV L=0.5 W=0.75
+ AD=0.07875 AS=0.157019 PD=0.96 PS=1.44231 NRD=12.7206 NRS=0 M=1 R=1.5
+ SA=250001 SB=250003 A=0.375 P=2.5 MULT=1
MM1017 N_A_489_107#_M1017_d N_D_M1017_g A_362_587# N_VPB_M1018_b PHV L=0.5
+ W=0.75 AD=0.105 AS=0.07875 PD=1.03 PS=0.96 NRD=0 NRS=12.7206 M=1 R=1.5
+ SA=250001 SB=250002 A=0.375 P=2.5 MULT=1
MM1003 A_660_587# N_A_30_587#_M1003_g N_A_489_107#_M1017_d N_VPB_M1018_b PHV
+ L=0.5 W=0.75 AD=0.07875 AS=0.105 PD=0.96 PS=1.03 NRD=12.7206 NRS=0 M=1 R=1.5
+ SA=250002 SB=250002 A=0.375 P=2.5 MULT=1
MM1012 N_VPWR_M1012_d N_SCD_M1012_g A_660_587# N_VPB_M1018_b PHV L=0.5 W=0.75
+ AD=0.105 AS=0.07875 PD=1.03 PS=0.96 NRD=0 NRS=12.7206 M=1 R=1.5 SA=250003
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1023 N_A_944_107#_M1023_d N_GATE_M1023_g N_VPWR_M1012_d N_VPB_M1018_b PHV
+ L=0.5 W=0.75 AD=0.21375 AS=0.105 PD=2.07 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250003 SB=250000 A=0.375 P=2.5 MULT=1
MM1014 N_A_1214_107#_M1014_d N_A_944_107#_M1014_g N_VPWR_M1014_s N_VPB_M1018_b
+ PHV L=0.5 W=0.75 AD=0.21375 AS=0.21375 PD=2.07 PS=2.07 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1007 N_A_1480_107#_M1007_d N_A_944_107#_M1007_g N_A_489_107#_M1007_s
+ N_VPB_M1018_b PHV L=0.5 W=0.75 AD=0.166635 AS=0.21375 PD=1.46795 PS=2.07 NRD=0
+ NRS=0 M=1 R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1000 A_1724_593# N_A_1214_107#_M1000_g N_A_1480_107#_M1007_d N_VPB_M1018_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0933154 PD=0.63 PS=0.822051 NRD=22.729 NRS=52.2958
+ M=1 R=0.84 SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1001 N_VPWR_M1001_d N_A_1678_81#_M1001_g A_1724_593# N_VPB_M1018_b PHV L=0.5
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1011 N_VPWR_M1011_d N_A_1480_107#_M1011_g N_A_1678_81#_M1011_s N_VPB_M1018_b
+ PHV L=0.5 W=0.42 AD=0.103622 AS=0.1197 PD=0.829062 PS=1.41 NRD=54.5687 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1021 N_Q_M1021_d N_A_1480_107#_M1021_g N_VPWR_M1011_d N_VPB_M1018_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.370078 PD=3.57 PS=2.96094 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
DX24_noxref N_VNB_M1004_b N_VPB_M1018_b NWDIODE A=31.668 P=29.56
*
.include "sky130_fd_sc_hvl__sdlxtp_1.pxi.spice"
*
.ends
*
*
