* File: sky130_fd_sc_hvl__diode_2.pxi.spice
* Created: Wed Sep  2 09:05:41 2020
* 
x_PM_SKY130_FD_SC_HVL__DIODE_2%VNB N_VNB_D0_noxref_pos VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__DIODE_2%VNB
x_PM_SKY130_FD_SC_HVL__DIODE_2%VPB N_VPB_X1_noxref_D1 VPB N_VPB_c_8_p VPB
+ PM_SKY130_FD_SC_HVL__DIODE_2%VPB
x_PM_SKY130_FD_SC_HVL__DIODE_2%DIODE N_DIODE_D0_noxref_neg DIODE DIODE DIODE
+ DIODE DIODE DIODE DIODE N_DIODE_c_9_n PM_SKY130_FD_SC_HVL__DIODE_2%DIODE
cc_1 N_VNB_D0_noxref_pos N_DIODE_c_9_n 0.146106f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=0.68
cc_2 N_VNB_c_2_p N_DIODE_c_9_n 0.00170391f $X=0.72 $Y=0 $X2=0.665 $Y2=0.68
cc_3 N_VNB_D0_noxref_pos VGND 0.0504029f $X=-0.33 $Y=-0.265 $X2=0.15 $Y2=0.535
cc_4 N_VNB_c_2_p VGND 0.102741f $X=0.72 $Y=0 $X2=0.15 $Y2=0.535
cc_5 N_VPB_X1_noxref_D1 N_DIODE_c_9_n 0.16193f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=0.68
cc_6 N_VPB_X1_noxref_D1 VPWR 0.0563655f $X=-0.33 $Y=1.885 $X2=0.15 $Y2=0.535
cc_7 VPB VPWR 0.102779f $X=0 $Y=3.955 $X2=0.15 $Y2=0.535
cc_8 N_VPB_c_8_p VPWR 0.00735982f $X=0.72 $Y=4.07 $X2=0.15 $Y2=0.535
cc_9 N_DIODE_c_9_n VGND 0.0697846f $X=0.665 $Y=0.68 $X2=0 $Y2=0
cc_10 N_DIODE_c_9_n VPWR 0.0431015f $X=0.665 $Y=0.68 $X2=0 $Y2=0
