* File: sky130_fd_sc_hvl__dfrtp_1.pex.spice
* Created: Fri Aug 28 09:34:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%VNB 5 7 11
r98 7 11 0.000463867 $w=1.536e-05 $l=5.7e-08 $layer=MET1_cond $X=7.68 $Y=0.057
+ $X2=7.68 $Y2=0
r99 5 11 0.58125 $w=1.7e-07 $l=2.72e-06 $layer=mcon $count=16 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r100 5 11 0.58125 $w=1.7e-07 $l=2.72e-06 $layer=mcon $count=16 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%VPB 4 6 14
c162 4 0 1.9686e-19 $X=-0.33 $Y=1.885
r163 10 14 0.58125 $w=1.7e-07 $l=2.72e-06 $layer=mcon $count=16 $X=15.12 $Y=4.07
+ $X2=15.12 $Y2=4.07
r164 9 14 970.781 $w=1.68e-07 $l=1.488e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=15.12 $Y2=4.07
r165 9 10 0.58125 $w=1.7e-07 $l=2.72e-06 $layer=mcon $count=16 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r166 6 10 0.000463867 $w=1.536e-05 $l=5.7e-08 $layer=MET1_cond $X=7.68 $Y=4.013
+ $X2=7.68 $Y2=4.07
r167 4 14 11.375 $w=1.7e-07 $l=1.51624e-05 $layer=licon1_NTAP_notbjt $count=16
+ $X=0 $Y=3.985 $X2=15.12 $Y2=4.07
r168 4 9 11.375 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=16
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%CLK 3 7 9 10 11 16
c30 16 0 3.93823e-20 $X=0.725 $Y=1.34
r31 16 19 54.0174 $w=5.2e-07 $l=5.25e-07 $layer=POLY_cond $X=0.675 $Y=1.34
+ $X2=0.675 $Y2=1.865
r32 16 18 26.237 $w=5.2e-07 $l=2.55e-07 $layer=POLY_cond $X=0.675 $Y=1.34
+ $X2=0.675 $Y2=1.085
r33 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.725 $Y=1.665
+ $X2=0.725 $Y2=2.035
r34 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.725 $Y=1.295
+ $X2=0.725 $Y2=1.665
r35 9 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.725
+ $Y=1.34 $X2=0.725 $Y2=1.34
r36 7 18 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.685 $Y=0.745 $X2=0.685
+ $Y2=1.085
r37 3 19 127.872 $w=5e-07 $l=1.195e-06 $layer=POLY_cond $X=0.665 $Y=3.06
+ $X2=0.665 $Y2=1.865
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%A_30_107# 1 2 9 13 15 17 19 21 22 24 31 34
+ 38 40 44 45 48 49 50 52 53 54 56 57 58 59 60 61 64 65 66 68 69 70 74 75 76 77
+ 80 81 83 84 87 91
c283 75 0 1.75956e-19 $X=9.165 $Y=2.05
c284 66 0 1.18092e-19 $X=6.75 $Y=3.72
c285 58 0 1.03544e-19 $X=3.7 $Y=3.72
c286 57 0 1.47925e-19 $X=5.1 $Y=3.72
c287 49 0 1.03544e-19 $X=2.67 $Y=3.72
c288 44 0 3.93823e-20 $X=1.405 $Y=2.02
c289 31 0 1.30273e-19 $X=10.195 $Y=1.185
c290 22 0 8.40164e-20 $X=10.195 $Y=0.935
r291 87 91 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=5.135 $Y=2.835
+ $X2=5.135 $Y2=3.37
r292 86 88 4.84127 $w=3.15e-07 $l=1.25e-07 $layer=LI1_cond $X=5.145 $Y=2.835
+ $X2=5.145 $Y2=2.96
r293 86 87 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.145
+ $Y=2.835 $X2=5.145 $Y2=2.835
r294 80 81 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.13
+ $Y=1.25 $X2=10.13 $Y2=1.25
r295 78 80 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=10.107 $Y=1.585
+ $X2=10.107 $Y2=1.25
r296 76 78 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=9.965 $Y=1.67
+ $X2=10.107 $Y2=1.585
r297 76 77 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=9.965 $Y=1.67
+ $X2=9.25 $Y2=1.67
r298 74 75 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.165
+ $Y=2.05 $X2=9.165 $Y2=2.05
r299 72 74 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=9.165 $Y=3.105
+ $X2=9.165 $Y2=2.05
r300 71 77 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.165 $Y=1.755
+ $X2=9.25 $Y2=1.67
r301 71 74 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.165 $Y=1.755
+ $X2=9.165 $Y2=2.05
r302 69 72 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.08 $Y=3.19
+ $X2=9.165 $Y2=3.105
r303 69 70 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=9.08 $Y=3.19
+ $X2=7.61 $Y2=3.19
r304 67 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.525 $Y=3.275
+ $X2=7.61 $Y2=3.19
r305 67 68 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.525 $Y=3.275
+ $X2=7.525 $Y2=3.635
r306 65 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.44 $Y=3.72
+ $X2=7.525 $Y2=3.635
r307 65 66 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.44 $Y=3.72
+ $X2=6.75 $Y2=3.72
r308 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.665 $Y=3.635
+ $X2=6.75 $Y2=3.72
r309 63 64 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.665 $Y=3.045
+ $X2=6.665 $Y2=3.635
r310 62 88 4.34843 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.31 $Y=2.96
+ $X2=5.145 $Y2=2.96
r311 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.58 $Y=2.96
+ $X2=6.665 $Y2=3.045
r312 61 62 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=6.58 $Y=2.96
+ $X2=5.31 $Y2=2.96
r313 59 88 5.86024 $w=3.15e-07 $l=1.03078e-07 $layer=LI1_cond $X=5.185 $Y=3.045
+ $X2=5.145 $Y2=2.96
r314 59 60 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.185 $Y=3.045
+ $X2=5.185 $Y2=3.635
r315 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.1 $Y=3.72
+ $X2=5.185 $Y2=3.635
r316 57 58 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=5.1 $Y=3.72 $X2=3.7
+ $Y2=3.72
r317 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.615 $Y=3.635
+ $X2=3.7 $Y2=3.72
r318 55 56 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.615 $Y=3.19
+ $X2=3.615 $Y2=3.635
r319 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.53 $Y=3.105
+ $X2=3.615 $Y2=3.19
r320 53 54 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.53 $Y=3.105
+ $X2=2.84 $Y2=3.105
r321 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.755 $Y=3.19
+ $X2=2.84 $Y2=3.105
r322 51 52 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.755 $Y=3.19
+ $X2=2.755 $Y2=3.635
r323 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.67 $Y=3.72
+ $X2=2.755 $Y2=3.635
r324 49 50 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=2.67 $Y=3.72
+ $X2=1.57 $Y2=3.72
r325 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.485 $Y=3.635
+ $X2=1.57 $Y2=3.72
r326 47 84 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.485 $Y=2.525
+ $X2=1.405 $Y2=2.44
r327 47 48 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=1.485 $Y=2.525
+ $X2=1.485 $Y2=3.635
r328 45 99 55.0463 $w=5.2e-07 $l=5.35e-07 $layer=POLY_cond $X=1.455 $Y=2.02
+ $X2=1.455 $Y2=2.555
r329 45 98 19.0347 $w=5.2e-07 $l=1.85e-07 $layer=POLY_cond $X=1.455 $Y=2.02
+ $X2=1.455 $Y2=1.835
r330 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.405
+ $Y=2.02 $X2=1.405 $Y2=2.02
r331 42 84 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.405 $Y=2.355
+ $X2=1.405 $Y2=2.44
r332 42 44 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.405 $Y=2.355
+ $X2=1.405 $Y2=2.02
r333 41 83 3.44808 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.44 $Y=2.44
+ $X2=0.275 $Y2=2.44
r334 40 84 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=2.44
+ $X2=1.405 $Y2=2.44
r335 40 41 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.24 $Y=2.44 $X2=0.44
+ $Y2=2.44
r336 36 83 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.275 $Y=2.525
+ $X2=0.275 $Y2=2.44
r337 36 38 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.275 $Y=2.525
+ $X2=0.275 $Y2=2.83
r338 32 83 3.14896 $w=3e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.245 $Y=2.355
+ $X2=0.275 $Y2=2.44
r339 32 34 68.7197 $w=2.68e-07 $l=1.61e-06 $layer=LI1_cond $X=0.245 $Y=2.355
+ $X2=0.245 $Y2=0.745
r340 31 81 7.24519 $w=4.8e-07 $l=6.5e-08 $layer=POLY_cond $X=10.205 $Y=1.185
+ $X2=10.205 $Y2=1.25
r341 29 75 65.3939 $w=4.55e-07 $l=5.35e-07 $layer=POLY_cond $X=9.102 $Y=2.585
+ $X2=9.102 $Y2=2.05
r342 27 87 17.656 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.135 $Y=2.67
+ $X2=5.135 $Y2=2.835
r343 22 31 26.7515 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=10.195 $Y=0.935
+ $X2=10.195 $Y2=1.185
r344 22 24 18.316 $w=5e-07 $l=1.9e-07 $layer=POLY_cond $X=10.195 $Y=0.935
+ $X2=10.195 $Y2=0.745
r345 19 29 27.2903 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=9.125 $Y=2.835
+ $X2=9.125 $Y2=2.585
r346 19 21 36.632 $w=5e-07 $l=3.8e-07 $layer=POLY_cond $X=9.125 $Y=2.835
+ $X2=9.125 $Y2=3.215
r347 15 27 91.9946 $w=3.72e-07 $l=7.1e-07 $layer=POLY_cond $X=4.425 $Y=2.372
+ $X2=5.135 $Y2=2.372
r348 15 17 107.006 $w=5e-07 $l=1e-06 $layer=POLY_cond $X=4.425 $Y=2.075
+ $X2=4.425 $Y2=1.075
r349 13 98 116.636 $w=5e-07 $l=1.09e-06 $layer=POLY_cond $X=1.465 $Y=0.745
+ $X2=1.465 $Y2=1.835
r350 9 99 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.445 $Y=3.06
+ $X2=1.445 $Y2=2.555
r351 2 38 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.685 $X2=0.275 $Y2=2.83
r352 1 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.535 $X2=0.295 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%RESET_B 3 7 10 13 16 20 24 25 28 29 31 32
+ 33 34 37 40 42 43 44 46 47 48 53 54 55 56 58 59 60 63 68
c192 56 0 4.39293e-20 $X=8.375 $Y=1.21
c193 53 0 3.10406e-20 $X=2.86 $Y=1.785
c194 48 0 1.30273e-19 $X=10.95 $Y=1.18
c195 42 0 1.7921e-20 $X=8.375 $Y=1.825
c196 34 0 1.02712e-19 $X=8.29 $Y=1.91
c197 33 0 9.70453e-20 $X=6.01 $Y=1.21
c198 3 0 1.03544e-19 $X=2.795 $Y=3.37
r199 59 69 50.2236 $w=5.7e-07 $l=5.25e-07 $layer=POLY_cond $X=11.65 $Y=1.23
+ $X2=11.65 $Y2=1.755
r200 59 68 16.4322 $w=5.7e-07 $l=1.65e-07 $layer=POLY_cond $X=11.65 $Y=1.23
+ $X2=11.65 $Y2=1.065
r201 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.62
+ $Y=1.23 $X2=11.62 $Y2=1.23
r202 54 64 46.5943 $w=6.4e-07 $l=5.25e-07 $layer=POLY_cond $X=2.865 $Y=1.785
+ $X2=2.865 $Y2=2.31
r203 54 63 35.3085 $w=6.4e-07 $l=3.9e-07 $layer=POLY_cond $X=2.865 $Y=1.785
+ $X2=2.865 $Y2=1.395
r204 53 55 9.76796 $w=5.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=1.785
+ $X2=2.965 $Y2=1.62
r205 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.86
+ $Y=1.785 $X2=2.86 $Y2=1.785
r206 51 60 11.407 $w=5.38e-07 $l=5.15e-07 $layer=LI1_cond $X=2.965 $Y=1.89
+ $X2=2.965 $Y2=2.405
r207 51 53 2.32571 $w=5.38e-07 $l=1.05e-07 $layer=LI1_cond $X=2.965 $Y=1.89
+ $X2=2.965 $Y2=1.785
r208 47 58 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.455 $Y=1.18
+ $X2=11.62 $Y2=1.18
r209 47 48 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=11.455 $Y=1.18
+ $X2=10.95 $Y2=1.18
r210 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.865 $Y=1.095
+ $X2=10.95 $Y2=1.18
r211 45 46 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=10.865 $Y=0.435
+ $X2=10.865 $Y2=1.095
r212 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.78 $Y=0.35
+ $X2=10.865 $Y2=0.435
r213 43 44 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=10.78 $Y=0.35
+ $X2=8.46 $Y2=0.35
r214 41 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.375 $Y=1.295
+ $X2=8.375 $Y2=1.21
r215 41 42 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.375 $Y=1.295
+ $X2=8.375 $Y2=1.825
r216 40 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.375 $Y=1.125
+ $X2=8.375 $Y2=1.21
r217 39 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.375 $Y=0.435
+ $X2=8.46 $Y2=0.35
r218 39 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.375 $Y=0.435
+ $X2=8.375 $Y2=1.125
r219 37 66 18.4754 $w=5.55e-07 $l=1.85e-07 $layer=POLY_cond $X=6.677 $Y=1.91
+ $X2=6.677 $Y2=1.725
r220 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.77
+ $Y=1.91 $X2=6.77 $Y2=1.91
r221 34 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.29 $Y=1.91
+ $X2=8.375 $Y2=1.825
r222 34 36 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=8.29 $Y=1.91
+ $X2=6.77 $Y2=1.91
r223 32 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.29 $Y=1.21
+ $X2=8.375 $Y2=1.21
r224 32 33 148.749 $w=1.68e-07 $l=2.28e-06 $layer=LI1_cond $X=8.29 $Y=1.21
+ $X2=6.01 $Y2=1.21
r225 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.925 $Y=1.125
+ $X2=6.01 $Y2=1.21
r226 30 31 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.925 $Y=0.63
+ $X2=5.925 $Y2=1.125
r227 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.84 $Y=0.545
+ $X2=5.925 $Y2=0.63
r228 28 29 169.952 $w=1.68e-07 $l=2.605e-06 $layer=LI1_cond $X=5.84 $Y=0.545
+ $X2=3.235 $Y2=0.545
r229 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.15 $Y=0.63
+ $X2=3.235 $Y2=0.545
r230 26 55 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=3.15 $Y=0.63
+ $X2=3.15 $Y2=1.62
r231 24 68 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.685 $Y=0.745
+ $X2=11.685 $Y2=1.065
r232 20 69 125.197 $w=5e-07 $l=1.17e-06 $layer=POLY_cond $X=11.615 $Y=2.925
+ $X2=11.615 $Y2=1.755
r233 16 25 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.705 $Y=3.37
+ $X2=6.705 $Y2=3.03
r234 13 25 27.3444 $w=5.55e-07 $l=2.77e-07 $layer=POLY_cond $X=6.677 $Y=2.753
+ $X2=6.677 $Y2=3.03
r235 12 37 8.86896 $w=5.55e-07 $l=9.2e-08 $layer=POLY_cond $X=6.677 $Y=2.002
+ $X2=6.677 $Y2=1.91
r236 12 13 72.3977 $w=5.55e-07 $l=7.51e-07 $layer=POLY_cond $X=6.677 $Y=2.002
+ $X2=6.677 $Y2=2.753
r237 10 66 69.5538 $w=5e-07 $l=6.5e-07 $layer=POLY_cond $X=6.65 $Y=1.075
+ $X2=6.65 $Y2=1.725
r238 7 63 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.935 $Y=1.075
+ $X2=2.935 $Y2=1.395
r239 3 64 113.426 $w=5e-07 $l=1.06e-06 $layer=POLY_cond $X=2.795 $Y=3.37
+ $X2=2.795 $Y2=2.31
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%D 3 6 7 8 9 14
c38 6 0 1.03544e-19 $X=3.61 $Y=3.05
r39 14 17 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.645 $Y=1.075
+ $X2=3.645 $Y2=1.6
r40 9 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.58 $Y=1.6
+ $X2=3.58 $Y2=1.6
r41 8 9 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.58 $Y=1.295
+ $X2=3.58 $Y2=1.6
r42 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.58 $Y=0.925 $X2=3.58
+ $Y2=1.295
r43 5 17 101.656 $w=5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.645 $Y=2.55 $X2=3.645
+ $Y2=1.6
r44 5 6 46.9324 $w=5.7e-07 $l=5e-07 $layer=POLY_cond $X=3.61 $Y=2.55 $X2=3.61
+ $Y2=3.05
r45 3 6 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.575 $Y=3.37 $X2=3.575
+ $Y2=3.05
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%A_339_537# 1 2 7 9 14 18 22 25 28 34 37 39
+ 40 41 43 44 45 46 47 48 51 57 58 63 66 71 73
c198 66 0 9.70453e-20 $X=5.205 $Y=1.075
c199 57 0 7.32434e-20 $X=9.84 $Y=2.035
c200 47 0 8.07904e-20 $X=9.695 $Y=2.035
c201 18 0 8.85078e-20 $X=9.647 $Y=1.525
c202 7 0 6.18503e-20 $X=9.195 $Y=1.395
r203 71 74 16.7639 $w=7.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.905 $Y=2.27
+ $X2=9.905 $Y2=2.435
r204 71 73 41.3539 $w=7.3e-07 $l=1.85e-07 $layer=POLY_cond $X=9.905 $Y=2.27
+ $X2=9.905 $Y2=2.085
r205 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.79
+ $Y=2.27 $X2=9.79 $Y2=2.27
r206 58 72 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=9.79 $Y=2.035
+ $X2=9.79 $Y2=2.27
r207 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=2.035
+ $X2=9.84 $Y2=2.035
r208 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=2.035
+ $X2=4.56 $Y2=2.035
r209 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=2.035
+ $X2=2.16 $Y2=2.035
r210 48 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=2.035
+ $X2=4.56 $Y2=2.035
r211 47 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=2.035
+ $X2=9.84 $Y2=2.035
r212 47 48 6.17573 $w=1.4e-07 $l=4.99e-06 $layer=MET1_cond $X=9.695 $Y=2.035
+ $X2=4.705 $Y2=2.035
r213 46 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=2.035
+ $X2=2.16 $Y2=2.035
r214 45 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.415 $Y=2.035
+ $X2=4.56 $Y2=2.035
r215 45 46 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=4.415 $Y=2.035
+ $X2=2.305 $Y2=2.035
r216 44 55 20.7941 $w=2.28e-07 $l=4.15e-07 $layer=LI1_cond $X=4.975 $Y=2.035
+ $X2=4.56 $Y2=2.035
r217 43 55 5.51168 $w=2.28e-07 $l=1.1e-07 $layer=LI1_cond $X=4.45 $Y=2.035
+ $X2=4.56 $Y2=2.035
r218 40 63 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=4.355 $Y=2.835
+ $X2=4.355 $Y2=3.37
r219 39 41 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=4.34 $Y=2.835
+ $X2=4.34 $Y2=2.67
r220 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.34
+ $Y=2.835 $X2=4.34 $Y2=2.835
r221 35 66 52.9679 $w=5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.205 $Y=1.57
+ $X2=5.205 $Y2=1.075
r222 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.14
+ $Y=1.57 $X2=5.14 $Y2=1.57
r223 32 44 7.10306 $w=2.3e-07 $l=2.14942e-07 $layer=LI1_cond $X=5.14 $Y=1.92
+ $X2=4.975 $Y2=2.035
r224 32 34 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=5.14 $Y=1.92
+ $X2=5.14 $Y2=1.57
r225 30 43 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.365 $Y=2.15
+ $X2=4.45 $Y2=2.035
r226 30 41 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.365 $Y=2.15
+ $X2=4.365 $Y2=2.67
r227 26 80 0.201461 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=1.875 $Y=2.15
+ $X2=1.875 $Y2=2.035
r228 26 28 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=1.875 $Y=2.15
+ $X2=1.875 $Y2=2.83
r229 25 51 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.885 $Y=2.035
+ $X2=2.16 $Y2=2.035
r230 25 80 0.501062 $w=2.28e-07 $l=1e-08 $layer=LI1_cond $X=1.885 $Y=2.035
+ $X2=1.875 $Y2=2.035
r231 25 37 39.4818 $w=2.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.885 $Y=1.92
+ $X2=1.885 $Y2=0.995
r232 20 37 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0.83
+ $X2=1.855 $Y2=0.995
r233 20 22 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=0.83
+ $X2=1.855 $Y2=0.745
r234 14 74 52.4329 $w=5e-07 $l=4.9e-07 $layer=POLY_cond $X=10.02 $Y=2.925
+ $X2=10.02 $Y2=2.435
r235 10 18 7.41015 $w=2.15e-07 $l=1.3e-07 $layer=POLY_cond $X=9.647 $Y=1.655
+ $X2=9.647 $Y2=1.525
r236 10 73 128.343 $w=2.15e-07 $l=4.3e-07 $layer=POLY_cond $X=9.647 $Y=1.655
+ $X2=9.647 $Y2=2.085
r237 7 18 107.982 $w=2.6e-07 $l=4.52e-07 $layer=POLY_cond $X=9.195 $Y=1.525
+ $X2=9.647 $Y2=1.525
r238 7 9 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.195 $Y=1.395
+ $X2=9.195 $Y2=0.91
r239 2 28 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=2.685 $X2=1.835 $Y2=2.83
r240 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.715
+ $Y=0.535 $X2=1.855 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%A_1119_506# 1 2 9 13 16 17 18 21 22 24 25
+ 28 32 35 36 37
c95 36 0 1.65819e-19 $X=8.735 $Y=2.26
c96 16 0 2.39819e-20 $X=5.892 $Y=3.03
c97 9 0 2.66018e-19 $X=5.845 $Y=3.37
r98 35 36 3.19717 $w=2.95e-07 $l=1.00995e-07 $layer=LI1_cond $X=8.77 $Y=2.175
+ $X2=8.735 $Y2=2.26
r99 35 37 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=8.77 $Y=2.175
+ $X2=8.77 $Y2=1.325
r100 30 37 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.805 $Y=1.16
+ $X2=8.805 $Y2=1.325
r101 30 32 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=8.805 $Y=1.16
+ $X2=8.805 $Y2=0.7
r102 26 36 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=8.735 $Y=2.345
+ $X2=8.735 $Y2=2.26
r103 26 28 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=8.735 $Y=2.345
+ $X2=8.735 $Y2=2.84
r104 24 36 3.3845 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.57 $Y=2.26
+ $X2=8.735 $Y2=2.26
r105 24 25 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=8.57 $Y=2.26
+ $X2=6.17 $Y2=2.26
r106 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.005
+ $Y=1.915 $X2=6.005 $Y2=1.915
r107 19 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.005 $Y=2.175
+ $X2=6.17 $Y2=2.26
r108 19 21 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=6.005 $Y=2.175
+ $X2=6.005 $Y2=1.915
r109 17 22 26.2929 $w=5.25e-07 $l=2.58e-07 $layer=POLY_cond $X=5.927 $Y=1.657
+ $X2=5.927 $Y2=1.915
r110 17 18 26.8714 $w=5.25e-07 $l=2.62e-07 $layer=POLY_cond $X=5.927 $Y=1.657
+ $X2=5.927 $Y2=1.395
r111 15 22 62.6749 $w=5.25e-07 $l=6.15e-07 $layer=POLY_cond $X=5.927 $Y=2.53
+ $X2=5.927 $Y2=1.915
r112 15 16 51.126 $w=5.25e-07 $l=5e-07 $layer=POLY_cond $X=5.892 $Y=2.53
+ $X2=5.892 $Y2=3.03
r113 13 18 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.915 $Y=1.075
+ $X2=5.915 $Y2=1.395
r114 9 16 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.845 $Y=3.37 $X2=5.845
+ $Y2=3.03
r115 2 28 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=8.595
+ $Y=2.715 $X2=8.735 $Y2=2.84
r116 1 32 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=8.665
+ $Y=0.535 $X2=8.805 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%A_921_632# 1 2 3 12 14 16 19 20 21 24 26 29
+ 32 36 39 40 43 47 48 54
r137 53 54 7.49041 $w=5e-07 $l=7e-08 $layer=POLY_cond $X=8.345 $Y=1.645
+ $X2=8.415 $Y2=1.645
r138 48 49 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.575 $Y=2.415
+ $X2=5.575 $Y2=2.61
r139 43 45 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.815 $Y=1.075
+ $X2=4.815 $Y2=1.16
r140 39 40 7.06528 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=4.745 $Y=3.325
+ $X2=4.745 $Y2=3.2
r141 34 36 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=7.095 $Y=2.695
+ $X2=7.095 $Y2=3.325
r142 33 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.66 $Y=2.61
+ $X2=5.575 $Y2=2.61
r143 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.93 $Y=2.61
+ $X2=7.095 $Y2=2.695
r144 32 33 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=6.93 $Y=2.61
+ $X2=5.66 $Y2=2.61
r145 30 53 42.8024 $w=5e-07 $l=4e-07 $layer=POLY_cond $X=7.945 $Y=1.645
+ $X2=8.345 $Y2=1.645
r146 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.945
+ $Y=1.56 $X2=7.945 $Y2=1.56
r147 27 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.66 $Y=1.56
+ $X2=5.575 $Y2=1.56
r148 27 29 149.075 $w=1.68e-07 $l=2.285e-06 $layer=LI1_cond $X=5.66 $Y=1.56
+ $X2=7.945 $Y2=1.56
r149 26 48 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.575 $Y=2.33
+ $X2=5.575 $Y2=2.415
r150 25 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.575 $Y=1.645
+ $X2=5.575 $Y2=1.56
r151 25 26 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.575 $Y=1.645
+ $X2=5.575 $Y2=2.33
r152 24 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.575 $Y=1.475
+ $X2=5.575 $Y2=1.56
r153 23 24 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.575 $Y=1.245
+ $X2=5.575 $Y2=1.475
r154 22 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.98 $Y=1.16
+ $X2=4.815 $Y2=1.16
r155 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.49 $Y=1.16
+ $X2=5.575 $Y2=1.245
r156 21 22 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.49 $Y=1.16
+ $X2=4.98 $Y2=1.16
r157 19 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.49 $Y=2.415
+ $X2=5.575 $Y2=2.415
r158 19 20 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.49 $Y=2.415
+ $X2=4.8 $Y2=2.415
r159 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.715 $Y=2.5
+ $X2=4.8 $Y2=2.415
r160 17 40 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.715 $Y=2.5
+ $X2=4.715 $Y2=3.2
r161 14 54 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.415 $Y=1.395
+ $X2=8.415 $Y2=1.645
r162 14 16 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=8.415 $Y=1.395
+ $X2=8.415 $Y2=0.91
r163 10 53 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.345 $Y=1.895
+ $X2=8.345 $Y2=1.645
r164 10 12 141.248 $w=5e-07 $l=1.32e-06 $layer=POLY_cond $X=8.345 $Y=1.895
+ $X2=8.345 $Y2=3.215
r165 3 36 600 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=6.955
+ $Y=3.16 $X2=7.095 $Y2=3.325
r166 2 39 600 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=4.605
+ $Y=3.16 $X2=4.745 $Y2=3.325
r167 1 43 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.675
+ $Y=0.865 $X2=4.815 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%A_2096_417# 1 2 9 13 16 19 20 23 25 26 29
+ 32 34 35 36 38
c88 9 0 1.88037e-19 $X=10.73 $Y=2.925
r89 33 36 4.55203 $w=1.97e-07 $l=9.80051e-08 $layer=LI1_cond $X=12.76 $Y=2.005
+ $X2=12.732 $Y2=1.92
r90 33 34 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=12.76 $Y=2.005
+ $X2=12.76 $Y2=2.535
r91 32 36 4.55203 $w=1.97e-07 $l=8.5e-08 $layer=LI1_cond $X=12.732 $Y=1.835
+ $X2=12.732 $Y2=1.92
r92 32 35 43.0245 $w=2.23e-07 $l=8.4e-07 $layer=LI1_cond $X=12.732 $Y=1.835
+ $X2=12.732 $Y2=0.995
r93 27 35 6.93655 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.785 $Y=0.83
+ $X2=12.785 $Y2=0.995
r94 27 29 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=12.785 $Y=0.83
+ $X2=12.785 $Y2=0.745
r95 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.675 $Y=2.62
+ $X2=12.76 $Y2=2.535
r96 25 26 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=12.675 $Y=2.62
+ $X2=12.09 $Y2=2.62
r97 21 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=11.965 $Y=2.705
+ $X2=12.09 $Y2=2.62
r98 21 23 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=11.965 $Y=2.705
+ $X2=11.965 $Y2=2.925
r99 19 36 1.88765 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=12.62 $Y=1.92
+ $X2=12.732 $Y2=1.92
r100 19 20 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=12.62 $Y=1.92
+ $X2=11.135 $Y2=1.92
r101 17 38 86.6748 $w=5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.905 $Y=1.555
+ $X2=10.905 $Y2=0.745
r102 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.97
+ $Y=1.555 $X2=10.97 $Y2=1.555
r103 14 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.97 $Y=1.835
+ $X2=11.135 $Y2=1.92
r104 14 16 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=10.97 $Y=1.835
+ $X2=10.97 $Y2=1.555
r105 12 17 56.7131 $w=5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.905 $Y=2.085
+ $X2=10.905 $Y2=1.555
r106 12 13 39.6318 $w=6.75e-07 $l=5e-07 $layer=POLY_cond $X=10.817 $Y=2.085
+ $X2=10.817 $Y2=2.585
r107 9 13 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=10.73 $Y=2.925
+ $X2=10.73 $Y2=2.585
r108 2 23 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.865
+ $Y=2.715 $X2=12.005 $Y2=2.925
r109 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.645
+ $Y=0.535 $X2=12.785 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%A_1875_543# 1 2 9 11 15 19 22 23 24 26 28
+ 30 32 34 37 39 40 42 43 54
c133 39 0 8.85078e-20 $X=10.515 $Y=2.185
c134 32 0 5.68085e-20 $X=10.135 $Y=2.76
r135 49 51 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.22 $Y=2.27
+ $X2=10.515 $Y2=2.27
r136 43 54 70.0889 $w=5e-07 $l=6.55e-07 $layer=POLY_cond $X=12.395 $Y=2.27
+ $X2=12.395 $Y2=2.925
r137 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.33
+ $Y=2.27 $X2=12.33 $Y2=2.27
r138 40 51 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=10.6 $Y=2.27
+ $X2=10.515 $Y2=2.27
r139 40 42 112.866 $w=1.68e-07 $l=1.73e-06 $layer=LI1_cond $X=10.6 $Y=2.27
+ $X2=12.33 $Y2=2.27
r140 39 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.515 $Y=2.185
+ $X2=10.515 $Y2=2.27
r141 38 39 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=10.515 $Y=0.785
+ $X2=10.515 $Y2=2.185
r142 36 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.22 $Y=2.355
+ $X2=10.22 $Y2=2.27
r143 36 37 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.22 $Y=2.355
+ $X2=10.22 $Y2=2.675
r144 35 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.76 $Y=0.7
+ $X2=9.595 $Y2=0.7
r145 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.43 $Y=0.7
+ $X2=10.515 $Y2=0.785
r146 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.43 $Y=0.7
+ $X2=9.76 $Y2=0.7
r147 33 48 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.68 $Y=2.76
+ $X2=9.555 $Y2=2.76
r148 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.135 $Y=2.76
+ $X2=10.22 $Y2=2.675
r149 32 33 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=10.135 $Y=2.76
+ $X2=9.68 $Y2=2.76
r150 28 48 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.555 $Y=2.845
+ $X2=9.555 $Y2=2.76
r151 28 30 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=9.555 $Y=2.845
+ $X2=9.555 $Y2=3.215
r152 24 46 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.595 $Y=0.785
+ $X2=9.595 $Y2=0.7
r153 24 26 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=9.595 $Y=0.785
+ $X2=9.595 $Y2=1.16
r154 21 43 19.7961 $w=5e-07 $l=1.85e-07 $layer=POLY_cond $X=12.395 $Y=2.085
+ $X2=12.395 $Y2=2.27
r155 21 22 20.4101 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=12.395 $Y=2.085
+ $X2=12.395 $Y2=1.835
r156 17 23 20.4101 $w=5e-07 $l=2.59808e-07 $layer=POLY_cond $X=13.82 $Y=2.085
+ $X2=13.8 $Y2=1.835
r157 17 19 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=13.82 $Y=2.085
+ $X2=13.82 $Y2=2.59
r158 13 23 20.4101 $w=5e-07 $l=2.59808e-07 $layer=POLY_cond $X=13.78 $Y=1.585
+ $X2=13.8 $Y2=1.835
r159 13 15 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=13.78 $Y=1.585
+ $X2=13.78 $Y2=1.245
r160 12 22 5.30422 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=12.645 $Y=1.835
+ $X2=12.395 $Y2=1.835
r161 11 23 5.30422 $w=5e-07 $l=2.7e-07 $layer=POLY_cond $X=13.53 $Y=1.835
+ $X2=13.8 $Y2=1.835
r162 11 12 94.7002 $w=5e-07 $l=8.85e-07 $layer=POLY_cond $X=13.53 $Y=1.835
+ $X2=12.645 $Y2=1.835
r163 7 22 20.4101 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=12.395 $Y=1.585
+ $X2=12.395 $Y2=1.835
r164 7 9 89.8849 $w=5e-07 $l=8.4e-07 $layer=POLY_cond $X=12.395 $Y=1.585
+ $X2=12.395 $Y2=0.745
r165 2 48 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=9.375
+ $Y=2.715 $X2=9.515 $Y2=2.84
r166 2 30 300 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_PDIFF $count=2 $X=9.375
+ $Y=2.715 $X2=9.515 $Y2=3.215
r167 1 46 182 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_NDIFF $count=1 $X=9.445
+ $Y=0.535 $X2=9.595 $Y2=0.7
r168 1 26 182 $w=1.7e-07 $l=6.95971e-07 $layer=licon1_NDIFF $count=1 $X=9.445
+ $Y=0.535 $X2=9.595 $Y2=1.16
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%A_2649_207# 1 2 9 13 17 20 23 27 28 30 31
r52 28 34 23.8503 $w=5.75e-07 $l=2.45e-07 $layer=POLY_cond $X=14.657 $Y=1.84
+ $X2=14.657 $Y2=2.085
r53 28 33 24.7808 $w=5.75e-07 $l=2.55e-07 $layer=POLY_cond $X=14.657 $Y=1.84
+ $X2=14.657 $Y2=1.585
r54 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.555
+ $Y=1.84 $X2=14.555 $Y2=1.84
r55 25 31 0.0811015 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=13.595 $Y=1.84
+ $X2=13.47 $Y2=1.84
r56 25 27 33.5256 $w=3.28e-07 $l=9.6e-07 $layer=LI1_cond $X=13.595 $Y=1.84
+ $X2=14.555 $Y2=1.84
r57 21 31 6.89714 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=13.47 $Y=2.005
+ $X2=13.47 $Y2=1.84
r58 21 23 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=13.47 $Y=2.005
+ $X2=13.47 $Y2=2.34
r59 20 31 6.89714 $w=2.3e-07 $l=1.74714e-07 $layer=LI1_cond $X=13.45 $Y=1.675
+ $X2=13.47 $Y2=1.84
r60 20 30 9.50649 $w=2.08e-07 $l=1.8e-07 $layer=LI1_cond $X=13.45 $Y=1.675
+ $X2=13.45 $Y2=1.495
r61 15 30 7.28026 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.39 $Y=1.33
+ $X2=13.39 $Y2=1.495
r62 15 17 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=13.39 $Y=1.33
+ $X2=13.39 $Y2=1.245
r63 13 34 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=14.695 $Y=2.965
+ $X2=14.695 $Y2=2.085
r64 9 33 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=14.675 $Y=1.08
+ $X2=14.675 $Y2=1.585
r65 2 23 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=13.285
+ $Y=2.215 $X2=13.43 $Y2=2.34
r66 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=13.245
+ $Y=1.035 $X2=13.39 $Y2=1.245
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%VPWR 1 2 3 4 5 6 7 22 25 32 44 53 57 66 75
+ 83
c124 83 0 1.88037e-19 $X=14.605 $Y=3.59
r125 81 83 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=13.885 $Y=3.63
+ $X2=14.605 $Y2=3.63
r126 80 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.605 $Y=3.59
+ $X2=14.605 $Y2=3.59
r127 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.885 $Y=3.59
+ $X2=13.885 $Y2=3.59
r128 78 80 5.42222 $w=9.43e-07 $l=4.2e-07 $layer=LI1_cond $X=14.247 $Y=3.17
+ $X2=14.247 $Y2=3.59
r129 75 78 10.4571 $w=9.43e-07 $l=8.1e-07 $layer=LI1_cond $X=14.247 $Y=2.36
+ $X2=14.247 $Y2=3.17
r130 72 81 0.310963 $w=3.7e-07 $l=8.1e-07 $layer=MET1_cond $X=13.075 $Y=3.63
+ $X2=13.885 $Y2=3.63
r131 70 72 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=12.355 $Y=3.63
+ $X2=13.075 $Y2=3.63
r132 69 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.075 $Y=3.59
+ $X2=13.075 $Y2=3.59
r133 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.355 $Y=3.59
+ $X2=12.355 $Y2=3.59
r134 66 69 8.17877 $w=8.93e-07 $l=6e-07 $layer=LI1_cond $X=12.717 $Y=2.99
+ $X2=12.717 $Y2=3.59
r135 63 70 0.397342 $w=3.7e-07 $l=1.035e-06 $layer=MET1_cond $X=11.32 $Y=3.63
+ $X2=12.355 $Y2=3.63
r136 61 63 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.6 $Y=3.63
+ $X2=11.32 $Y2=3.63
r137 60 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.32 $Y=3.59
+ $X2=11.32 $Y2=3.59
r138 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.6 $Y=3.59
+ $X2=10.6 $Y2=3.59
r139 57 60 8.54 $w=9.48e-07 $l=6.65e-07 $layer=LI1_cond $X=10.96 $Y=2.925
+ $X2=10.96 $Y2=3.59
r140 54 61 0.758213 $w=3.7e-07 $l=1.975e-06 $layer=MET1_cond $X=8.625 $Y=3.63
+ $X2=10.6 $Y2=3.63
r141 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.625 $Y=3.59
+ $X2=8.625 $Y2=3.59
r142 49 54 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.905 $Y=3.63
+ $X2=8.625 $Y2=3.63
r143 48 53 27.6586 $w=2.98e-07 $l=7.2e-07 $layer=LI1_cond $X=7.905 $Y=3.605
+ $X2=8.625 $Y2=3.605
r144 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.905 $Y=3.59
+ $X2=7.905 $Y2=3.59
r145 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.285 $Y=3.59
+ $X2=6.285 $Y2=3.59
r146 42 44 1.24592 $w=4.78e-07 $l=5e-08 $layer=LI1_cond $X=6.235 $Y=3.465
+ $X2=6.285 $Y2=3.465
r147 39 45 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.565 $Y=3.63
+ $X2=6.285 $Y2=3.63
r148 38 42 16.6953 $w=4.78e-07 $l=6.7e-07 $layer=LI1_cond $X=5.565 $Y=3.465
+ $X2=6.235 $Y2=3.465
r149 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.565 $Y=3.59
+ $X2=5.565 $Y2=3.59
r150 35 39 0.93289 $w=3.7e-07 $l=2.43e-06 $layer=MET1_cond $X=3.135 $Y=3.63
+ $X2=5.565 $Y2=3.63
r151 32 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.135 $Y=3.59
+ $X2=3.135 $Y2=3.59
r152 29 35 0.779328 $w=3.7e-07 $l=2.03e-06 $layer=MET1_cond $X=1.105 $Y=3.63
+ $X2=3.135 $Y2=3.63
r153 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.105 $Y=3.59
+ $X2=1.105 $Y2=3.59
r154 25 28 15.8126 $w=5.88e-07 $l=7.8e-07 $layer=LI1_cond $X=0.925 $Y=2.81
+ $X2=0.925 $Y2=3.59
r155 22 49 0.0863787 $w=3.7e-07 $l=2.25e-07 $layer=MET1_cond $X=7.68 $Y=3.63
+ $X2=7.905 $Y2=3.63
r156 22 45 0.535548 $w=3.7e-07 $l=1.395e-06 $layer=MET1_cond $X=7.68 $Y=3.63
+ $X2=6.285 $Y2=3.63
r157 7 78 300 $w=1.7e-07 $l=1.06604e-06 $layer=licon1_PDIFF $count=2 $X=14.07
+ $Y=2.215 $X2=14.305 $Y2=3.17
r158 7 75 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=14.07
+ $Y=2.215 $X2=14.305 $Y2=2.36
r159 6 66 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=12.645
+ $Y=2.715 $X2=12.785 $Y2=2.99
r160 5 57 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=10.98
+ $Y=2.715 $X2=11.12 $Y2=2.925
r161 4 48 600 $w=1.7e-07 $l=9.19647e-07 $layer=licon1_PDIFF $count=1 $X=7.81
+ $Y=2.715 $X2=7.955 $Y2=3.565
r162 3 42 600 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=6.095
+ $Y=3.16 $X2=6.235 $Y2=3.38
r163 2 32 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=3.16 $X2=3.185 $Y2=3.455
r164 1 25 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.915
+ $Y=2.685 $X2=1.055 $Y2=2.81
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%A_452_632# 1 2 3 12 14 15 17 20 24 28 29 30
+ 31
r63 28 29 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=3.99 $Y=2.32
+ $X2=3.99 $Y2=2.49
r64 28 31 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=4.015 $Y=2.32
+ $X2=4.015 $Y2=1.325
r65 22 31 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.065 $Y=1.19
+ $X2=4.065 $Y2=1.325
r66 22 24 4.90855 $w=2.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.065 $Y=1.19
+ $X2=4.065 $Y2=1.075
r67 18 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.965 $Y=2.84
+ $X2=3.965 $Y2=2.755
r68 18 20 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.965 $Y=2.84
+ $X2=3.965 $Y2=3.285
r69 17 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.965 $Y=2.67
+ $X2=3.965 $Y2=2.755
r70 17 29 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.965 $Y=2.67
+ $X2=3.965 $Y2=2.49
r71 14 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=2.755
+ $X2=3.965 $Y2=2.755
r72 14 15 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=3.88 $Y=2.755
+ $X2=2.49 $Y2=2.755
r73 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.365 $Y=2.84
+ $X2=2.49 $Y2=2.755
r74 10 12 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.365 $Y=2.84
+ $X2=2.365 $Y2=3.285
r75 3 20 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.825
+ $Y=3.16 $X2=3.965 $Y2=3.285
r76 2 12 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.26
+ $Y=3.16 $X2=2.405 $Y2=3.285
r77 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.895
+ $Y=0.865 $X2=4.035 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%Q 1 2 7 8 9 10 11 12 13 22
r12 13 40 14.6205 $w=3.33e-07 $l=4.25e-07 $layer=LI1_cond $X=15.067 $Y=3.145
+ $X2=15.067 $Y2=3.57
r13 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=15.067 $Y=2.775
+ $X2=15.067 $Y2=3.145
r14 11 12 14.2765 $w=3.33e-07 $l=4.15e-07 $layer=LI1_cond $X=15.067 $Y=2.36
+ $X2=15.067 $Y2=2.775
r15 10 11 11.1804 $w=3.33e-07 $l=3.25e-07 $layer=LI1_cond $X=15.067 $Y=2.035
+ $X2=15.067 $Y2=2.36
r16 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=15.067 $Y=1.665
+ $X2=15.067 $Y2=2.035
r17 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=15.067 $Y=1.295
+ $X2=15.067 $Y2=1.665
r18 7 8 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=15.067 $Y=0.925
+ $X2=15.067 $Y2=1.295
r19 7 22 3.26812 $w=3.33e-07 $l=9.5e-08 $layer=LI1_cond $X=15.067 $Y=0.925
+ $X2=15.067 $Y2=0.83
r20 2 40 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=14.945
+ $Y=2.215 $X2=15.085 $Y2=3.57
r21 2 11 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=14.945
+ $Y=2.215 $X2=15.085 $Y2=2.36
r22 1 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=14.925
+ $Y=0.705 $X2=15.065 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_HVL__DFRTP_1%VGND 1 2 3 4 5 16 19 28 41 51 55 59
c87 51 0 8.40164e-20 $X=11.965 $Y=0.48
r88 61 63 6.42105 $w=9.48e-07 $l=5e-07 $layer=LI1_cond $X=14.21 $Y=0.83
+ $X2=14.21 $Y2=1.33
r89 56 59 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=13.85 $Y=0.44
+ $X2=14.57 $Y2=0.44
r90 55 61 4.49474 $w=9.48e-07 $l=3.5e-07 $layer=LI1_cond $X=14.21 $Y=0.48
+ $X2=14.21 $Y2=0.83
r91 55 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.57 $Y=0.48
+ $X2=14.57 $Y2=0.48
r92 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.85 $Y=0.48
+ $X2=13.85 $Y2=0.48
r93 52 56 0.723662 $w=3.7e-07 $l=1.885e-06 $layer=MET1_cond $X=11.965 $Y=0.44
+ $X2=13.85 $Y2=0.44
r94 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.965 $Y=0.48
+ $X2=11.965 $Y2=0.48
r95 49 51 14.5704 $w=5.48e-07 $l=6.7e-07 $layer=LI1_cond $X=11.295 $Y=0.64
+ $X2=11.965 $Y2=0.64
r96 46 52 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=11.245 $Y=0.44
+ $X2=11.965 $Y2=0.44
r97 45 49 1.08734 $w=5.48e-07 $l=5e-08 $layer=LI1_cond $X=11.245 $Y=0.64
+ $X2=11.295 $Y2=0.64
r98 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.245 $Y=0.48
+ $X2=11.245 $Y2=0.48
r99 42 46 1.24769 $w=3.7e-07 $l=3.25e-06 $layer=MET1_cond $X=7.995 $Y=0.44
+ $X2=11.245 $Y2=0.44
r100 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.995 $Y=0.48
+ $X2=7.995 $Y2=0.48
r101 39 41 1.0311 $w=5.78e-07 $l=5e-08 $layer=LI1_cond $X=7.945 $Y=0.655
+ $X2=7.995 $Y2=0.655
r102 35 39 13.8168 $w=5.78e-07 $l=6.7e-07 $layer=LI1_cond $X=7.275 $Y=0.655
+ $X2=7.945 $Y2=0.655
r103 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.275 $Y=0.48
+ $X2=7.275 $Y2=0.48
r104 29 36 1.76596 $w=3.7e-07 $l=4.6e-06 $layer=MET1_cond $X=2.675 $Y=0.44
+ $X2=7.275 $Y2=0.44
r105 28 32 12.0621 $w=5.88e-07 $l=5.95e-07 $layer=LI1_cond $X=2.495 $Y=0.48
+ $X2=2.495 $Y2=1.075
r106 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.675 $Y=0.48
+ $X2=2.675 $Y2=0.48
r107 23 29 0.491399 $w=3.7e-07 $l=1.28e-06 $layer=MET1_cond $X=1.395 $Y=0.44
+ $X2=2.675 $Y2=0.44
r108 20 23 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.675 $Y=0.44
+ $X2=1.395 $Y2=0.44
r109 19 25 3.40316 $w=9.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.035 $Y=0.48
+ $X2=1.035 $Y2=0.745
r110 19 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.395 $Y=0.48
+ $X2=1.395 $Y2=0.48
r111 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.675 $Y=0.48
+ $X2=0.675 $Y2=0.48
r112 16 42 0.12093 $w=3.7e-07 $l=3.15e-07 $layer=MET1_cond $X=7.68 $Y=0.44
+ $X2=7.995 $Y2=0.44
r113 16 36 0.155482 $w=3.7e-07 $l=4.05e-07 $layer=MET1_cond $X=7.68 $Y=0.44
+ $X2=7.275 $Y2=0.44
r114 5 63 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=14.03
+ $Y=1.035 $X2=14.285 $Y2=1.33
r115 5 61 182 $w=1.7e-07 $l=3.42491e-07 $layer=licon1_NDIFF $count=1 $X=14.03
+ $Y=1.035 $X2=14.285 $Y2=0.83
r116 4 49 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.155
+ $Y=0.535 $X2=11.295 $Y2=0.745
r117 3 39 182 $w=1.7e-07 $l=1.09624e-06 $layer=licon1_NDIFF $count=1 $X=6.9
+ $Y=0.865 $X2=7.945 $Y2=0.76
r118 2 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.4
+ $Y=0.865 $X2=2.545 $Y2=1.075
r119 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.935
+ $Y=0.535 $X2=1.075 $Y2=0.745
.ends

