* File: sky130_fd_sc_hvl__a22oi_1.pex.spice
* Created: Fri Aug 28 09:32:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__A22OI_1%VNB 5 7 11 25
r23 7 25 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=0.057
+ $X2=1.92 $Y2=0.058
r24 7 11 0.00185547 $w=3.84e-06 $l=5.7e-08 $layer=MET1_cond $X=1.92 $Y=0.057
+ $X2=1.92 $Y2=0
r25 5 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r26 5 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__A22OI_1%VPB 4 6 14 21
r36 10 21 0.00185547 $w=3.84e-06 $l=5.7e-08 $layer=MET1_cond $X=1.92 $Y=4.07
+ $X2=1.92 $Y2=4.013
r37 10 14 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=4.07
+ $X2=3.6 $Y2=4.07
r38 9 14 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=3.6
+ $Y2=4.07
r39 9 10 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r40 6 21 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=4.012
+ $X2=1.92 $Y2=4.013
r41 4 14 45.5 $w=1.7e-07 $l=3.64225e-06 $layer=licon1_NTAP_notbjt $count=4 $X=0
+ $Y=3.985 $X2=3.6 $Y2=4.07
r42 4 9 45.5 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=4 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__A22OI_1%B2 3 7 9 10 14
r29 14 17 39.8984 $w=5.7e-07 $l=4.15e-07 $layer=POLY_cond $X=0.735 $Y=1.67
+ $X2=0.735 $Y2=2.085
r30 14 16 24.8801 $w=5.7e-07 $l=2.55e-07 $layer=POLY_cond $X=0.735 $Y=1.67
+ $X2=0.735 $Y2=1.415
r31 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=1.67 $X2=0.635 $Y2=1.67
r32 9 10 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=0.24 $Y=1.67
+ $X2=0.635 $Y2=1.67
r33 7 16 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.77 $Y=0.91 $X2=0.77
+ $Y2=1.415
r34 3 17 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.7 $Y=2.965 $X2=0.7
+ $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_HVL__A22OI_1%B1 3 7 9 12
r40 12 15 28.1653 $w=5.7e-07 $l=2.9e-07 $layer=POLY_cond $X=1.515 $Y=1.625
+ $X2=1.515 $Y2=1.915
r41 12 14 20.6562 $w=5.7e-07 $l=2.1e-07 $layer=POLY_cond $X=1.515 $Y=1.625
+ $X2=1.515 $Y2=1.415
r42 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.625 $X2=1.63 $Y2=1.625
r43 7 15 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=1.48 $Y=2.965 $X2=1.48
+ $Y2=1.915
r44 3 14 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.48 $Y=0.91 $X2=1.48
+ $Y2=1.415
.ends

.subckt PM_SKY130_FD_SC_HVL__A22OI_1%A1 1 2 6 12
c27 6 0 1.4473e-19 $X=2.26 $Y=0.91
r28 9 12 142.853 $w=5e-07 $l=1.335e-06 $layer=POLY_cond $X=2.26 $Y=1.63 $X2=2.26
+ $Y2=2.965
r29 6 9 77.0442 $w=5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.26 $Y=0.91 $X2=2.26
+ $Y2=1.63
r30 1 2 22.5785 $w=2.43e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.627 $X2=2.64
+ $Y2=1.627
r31 1 9 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21 $Y=1.63
+ $X2=2.21 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HVL__A22OI_1%A2 3 7 9 10 14
c21 10 0 1.4473e-19 $X=3.6 $Y=1.665
r22 14 17 43.653 $w=5.7e-07 $l=4.55e-07 $layer=POLY_cond $X=3.005 $Y=1.63
+ $X2=3.005 $Y2=2.085
r23 14 16 21.1255 $w=5.7e-07 $l=2.15e-07 $layer=POLY_cond $X=3.005 $Y=1.63
+ $X2=3.005 $Y2=1.415
r24 9 10 23.2841 $w=2.43e-07 $l=4.95e-07 $layer=LI1_cond $X=3.105 $Y=1.627
+ $X2=3.6 $Y2=1.627
r25 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.105
+ $Y=1.63 $X2=3.105 $Y2=1.63
r26 7 17 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.04 $Y=2.965 $X2=3.04
+ $Y2=2.085
r27 3 16 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.97 $Y=0.91 $X2=2.97
+ $Y2=1.415
.ends

.subckt PM_SKY130_FD_SC_HVL__A22OI_1%A_33_443# 1 2 3 12 16 17 21 24 25 28
r47 28 30 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=3.43 $Y=2.34
+ $X2=3.43 $Y2=3.59
r48 26 28 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.43 $Y=2.1 $X2=3.43
+ $Y2=2.34
r49 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.265 $Y=2.015
+ $X2=3.43 $Y2=2.1
r50 24 25 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=3.265 $Y=2.015
+ $X2=1.955 $Y2=2.015
r51 21 23 57.6222 $w=2.48e-07 $l=1.25e-06 $layer=LI1_cond $X=1.83 $Y=2.34
+ $X2=1.83 $Y2=3.59
r52 19 23 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=1.83 $Y=3.635
+ $X2=1.83 $Y2=3.59
r53 18 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.83 $Y=2.1
+ $X2=1.955 $Y2=2.015
r54 18 21 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=1.83 $Y=2.1 $X2=1.83
+ $Y2=2.34
r55 16 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.705 $Y=3.72
+ $X2=1.83 $Y2=3.635
r56 16 17 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=1.705 $Y=3.72
+ $X2=0.475 $Y2=3.72
r57 12 15 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=0.31 $Y=2.34
+ $X2=0.31 $Y2=3.59
r58 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.31 $Y=3.635
+ $X2=0.475 $Y2=3.72
r59 10 15 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.31 $Y=3.635
+ $X2=0.31 $Y2=3.59
r60 3 30 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=3.29
+ $Y=2.215 $X2=3.43 $Y2=3.59
r61 3 28 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=3.29
+ $Y=2.215 $X2=3.43 $Y2=2.34
r62 2 23 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.73
+ $Y=2.215 $X2=1.87 $Y2=3.59
r63 2 21 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.73
+ $Y=2.215 $X2=1.87 $Y2=2.34
r64 1 15 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=2.215 $X2=0.31 $Y2=3.59
r65 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=2.215 $X2=0.31 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__A22OI_1%Y 1 2 9 13 14 15 16 17 18 19 20 21 32 43
r46 41 59 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=1.105 $Y=2.355
+ $X2=1.105 $Y2=2.34
r47 41 43 1.60062 $w=3.58e-07 $l=5e-08 $layer=LI1_cond $X=1.105 $Y=2.355
+ $X2=1.105 $Y2=2.405
r48 21 50 7.20277 $w=3.58e-07 $l=2.25e-07 $layer=LI1_cond $X=1.105 $Y=3.145
+ $X2=1.105 $Y2=3.37
r49 20 21 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.105 $Y=2.775
+ $X2=1.105 $Y2=3.145
r50 19 59 0.0960369 $w=3.58e-07 $l=3e-09 $layer=LI1_cond $X=1.105 $Y=2.337
+ $X2=1.105 $Y2=2.34
r51 19 57 7.44475 $w=3.58e-07 $l=1.62e-07 $layer=LI1_cond $X=1.105 $Y=2.337
+ $X2=1.105 $Y2=2.175
r52 19 20 11.3003 $w=3.58e-07 $l=3.53e-07 $layer=LI1_cond $X=1.105 $Y=2.422
+ $X2=1.105 $Y2=2.775
r53 19 43 0.544209 $w=3.58e-07 $l=1.7e-08 $layer=LI1_cond $X=1.105 $Y=2.422
+ $X2=1.105 $Y2=2.405
r54 18 57 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=1.185 $Y=2.035
+ $X2=1.185 $Y2=2.175
r55 17 18 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.185 $Y=1.665
+ $X2=1.185 $Y2=2.035
r56 16 17 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.185 $Y=1.295
+ $X2=1.185 $Y2=1.665
r57 15 32 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.895
+ $X2=1.185 $Y2=0.98
r58 15 16 16.6364 $w=1.98e-07 $l=3e-07 $layer=LI1_cond $X=1.185 $Y=0.995
+ $X2=1.185 $Y2=1.295
r59 15 32 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.185 $Y=0.995
+ $X2=1.185 $Y2=0.98
r60 13 15 16.9204 $w=3.08e-07 $l=4.2e-07 $layer=LI1_cond $X=1.705 $Y=0.895
+ $X2=1.285 $Y2=0.895
r61 13 14 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.705 $Y=0.895
+ $X2=1.83 $Y2=0.895
r62 7 14 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=0.81 $X2=1.83
+ $Y2=0.895
r63 7 9 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=1.83 $Y=0.81 $X2=1.83
+ $Y2=0.66
r64 2 59 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.95
+ $Y=2.215 $X2=1.09 $Y2=2.34
r65 2 50 300 $w=1.7e-07 $l=1.223e-06 $layer=licon1_PDIFF $count=2 $X=0.95
+ $Y=2.215 $X2=1.09 $Y2=3.37
r66 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.73
+ $Y=0.535 $X2=1.87 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__A22OI_1%VPWR 1 4 7 14
r25 11 14 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.25 $Y=3.63
+ $X2=2.97 $Y2=3.63
r26 10 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.97 $Y=3.59
+ $X2=2.97 $Y2=3.59
r27 10 11 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.25 $Y=3.59
+ $X2=2.25 $Y2=3.59
r28 7 10 15.7316 $w=9.48e-07 $l=1.225e-06 $layer=LI1_cond $X=2.61 $Y=2.365
+ $X2=2.61 $Y2=3.59
r29 4 11 0.126689 $w=3.7e-07 $l=3.3e-07 $layer=MET1_cond $X=1.92 $Y=3.63
+ $X2=2.25 $Y2=3.63
r30 1 10 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.51
+ $Y=2.215 $X2=2.65 $Y2=3.59
r31 1 7 300 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=2 $X=2.51
+ $Y=2.215 $X2=2.65 $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_HVL__A22OI_1%VGND 1 2 7 10 17 21
r29 18 21 0.552824 $w=3.7e-07 $l=1.44e-06 $layer=MET1_cond $X=2.22 $Y=0.44
+ $X2=3.66 $Y2=0.44
r30 17 23 1.35975 $w=1.613e-06 $l=1.8e-07 $layer=LI1_cond $X=2.942 $Y=0.48
+ $X2=2.942 $Y2=0.66
r31 17 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.66 $Y=0.48
+ $X2=3.66 $Y2=0.48
r32 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.22 $Y=0.48
+ $X2=2.22 $Y2=0.48
r33 10 14 3.64905 $w=5.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.385 $Y=0.48
+ $X2=0.385 $Y2=0.66
r34 10 11 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.565 $Y=0.48
+ $X2=0.565 $Y2=0.48
r35 7 18 0.115172 $w=3.7e-07 $l=3e-07 $layer=MET1_cond $X=1.92 $Y=0.44 $X2=2.22
+ $Y2=0.44
r36 7 11 0.520192 $w=3.7e-07 $l=1.355e-06 $layer=MET1_cond $X=1.92 $Y=0.44
+ $X2=0.565 $Y2=0.44
r37 2 23 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.22
+ $Y=0.535 $X2=3.36 $Y2=0.66
r38 1 14 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.235
+ $Y=0.535 $X2=0.38 $Y2=0.66
.ends

