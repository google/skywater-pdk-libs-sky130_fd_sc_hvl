* NGSPICE file created from sky130_fd_sc_hvl__dfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
M1000 a_1494_539# a_30_112# a_1063_85# VPB phv w=1e+06u l=500000u
+  ad=3.112e+11p pd=2.75e+06u as=2.8e+11p ps=2.56e+06u
M1001 VPWR a_1711_85# Q VPB phv w=1.5e+06u l=500000u
+  ad=1.8596e+12p pd=1.629e+07u as=3.975e+11p ps=3.53e+06u
M1002 a_1669_539# a_339_112# a_1494_539# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1003 a_1711_85# a_1494_539# VPWR VPB phv w=1e+06u l=500000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1004 a_339_112# a_30_112# VGND VNB nhv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=1.2345e+12p ps=1.183e+07u
M1005 VPWR a_1711_85# a_2365_443# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u
M1006 a_709_111# D VPWR VPB phv w=420000u l=500000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1007 a_1669_111# a_30_112# a_1494_539# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1008 VPWR a_1711_85# a_1669_539# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1711_85# a_1494_539# VGND VNB nhv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
M1010 VGND a_1711_85# Q VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u
M1011 a_1021_539# a_30_112# a_865_111# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1012 VPWR CLK a_30_112# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=2.1375e+11p ps=2.07e+06u
M1013 a_709_111# D VGND VNB nhv w=420000u l=500000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1014 VGND a_1711_85# a_2365_443# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1015 VPWR a_1063_85# a_1021_539# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_1711_85# a_1669_111# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1063_85# a_865_111# VPWR VPB phv w=1e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1021_111# a_339_112# a_865_111# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1019 a_865_111# a_339_112# a_709_111# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Q_N a_2365_443# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=0p ps=0u
M1021 VGND a_1063_85# a_1021_111# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_339_112# a_30_112# VPWR VPB phv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
M1023 a_1063_85# a_865_111# VGND VNB nhv w=750000u l=500000u
+  ad=2.4495e+11p pd=2.25e+06u as=0p ps=0u
M1024 a_1494_539# a_339_112# a_1063_85# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND CLK a_30_112# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1026 a_865_111# a_30_112# a_709_111# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q_N a_2365_443# VGND VNB nhv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
.ends

