* File: sky130_fd_sc_hvl__xnor2_1.spice
* Created: Fri Aug 28 09:40:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__xnor2_1.pex.spice"
.subckt sky130_fd_sc_hvl__xnor2_1  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1004 A_222_107# N_B_M1004_g N_A_30_107#_M1004_s N_VNB_M1004_b NHV L=0.5 W=0.75
+ AD=0.07875 AS=0.345 PD=0.96 PS=2.42 NRD=7.5924 NRS=29.64 M=1 R=1.5 SA=250000
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g A_222_107# N_VNB_M1004_b NHV L=0.5 W=0.75
+ AD=0.110625 AS=0.07875 PD=1.045 PS=0.96 NRD=0 NRS=7.5924 M=1 R=1.5 SA=250001
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1008 N_A_523_107#_M1008_d N_A_M1008_g N_VGND_M1005_d N_VNB_M1004_b NHV L=0.5
+ W=0.75 AD=0.10875 AS=0.110625 PD=1.04 PS=1.045 NRD=0 NRS=2.2686 M=1 R=1.5
+ SA=250002 SB=250001 A=0.375 P=2.5 MULT=1
MM1006 N_VGND_M1006_d N_B_M1006_g N_A_523_107#_M1008_d N_VNB_M1004_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.10875 PD=2.07 PS=1.04 NRD=0 NRS=1.5162 M=1 R=1.5
+ SA=250003 SB=250000 A=0.375 P=2.5 MULT=1
MM1002 N_Y_M1002_d N_A_30_107#_M1002_g N_A_523_107#_M1002_s N_VNB_M1004_b NHV
+ L=0.5 W=0.75 AD=0.21375 AS=0.21375 PD=2.07 PS=2.07 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1009 N_A_30_107#_M1009_d N_B_M1009_g N_VPWR_M1009_s N_VPB_M1009_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.4275 PD=1.78 PS=3.57 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250004 A=0.75 P=4 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_30_107#_M1009_d N_VPB_M1009_b PHV L=0.5
+ W=1.5 AD=0.22875 AS=0.21 PD=1.805 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001
+ SB=250003 A=0.75 P=4 MULT=1
MM1000 A_539_443# N_A_M1000_g N_VPWR_M1003_d N_VPB_M1009_b PHV L=0.5 W=1.5
+ AD=0.1575 AS=0.22875 PD=1.71 PS=1.805 NRD=6.3603 NRS=3.1706 M=1 R=3 SA=250002
+ SB=250002 A=0.75 P=4 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g A_539_443# N_VPB_M1009_b PHV L=0.5 W=1.5
+ AD=0.63375 AS=0.1575 PD=2.345 PS=1.71 NRD=71.9306 NRS=6.3603 M=1 R=3 SA=250002
+ SB=250001 A=0.75 P=4 MULT=1
MM1007 N_VPWR_M1007_d N_A_30_107#_M1007_g N_Y_M1001_d N_VPB_M1009_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.63375 PD=3.57 PS=2.345 NRD=0 NRS=0 M=1 R=3 SA=250004
+ SB=250000 A=0.75 P=4 MULT=1
DX10_noxref N_VNB_M1004_b N_VPB_M1009_b NWDIODE A=15.444 P=17.08
*
.include "sky130_fd_sc_hvl__xnor2_1.pxi.spice"
*
.ends
*
*
