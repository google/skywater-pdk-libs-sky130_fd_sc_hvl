# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__inv_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__inv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  9.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.310000 1.580000 6.760000 1.815000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.520000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.195000 0.730000 1.405000 1.230000 ;
        RECT 1.195000 1.230000 7.110000 1.395000 ;
        RECT 1.195000 1.395000 6.225000 1.400000 ;
        RECT 1.275000 2.035000 7.110000 2.205000 ;
        RECT 1.275000 2.205000 1.605000 3.445000 ;
        RECT 2.755000 0.730000 2.965000 1.230000 ;
        RECT 2.835000 2.205000 3.165000 3.445000 ;
        RECT 4.315000 0.730000 4.525000 1.230000 ;
        RECT 4.395000 2.205000 4.725000 3.445000 ;
        RECT 5.915000 0.730000 6.565000 1.225000 ;
        RECT 5.915000 1.225000 7.110000 1.230000 ;
        RECT 5.955000 2.205000 6.285000 3.445000 ;
        RECT 6.940000 1.395000 7.110000 2.035000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.380000 7.105000 0.550000 ;
        RECT 0.095000 0.550000 0.985000 1.385000 ;
        RECT 1.575000 0.550000 2.585000 1.045000 ;
        RECT 3.135000 0.550000 4.145000 1.045000 ;
        RECT 4.695000 0.550000 5.745000 1.045000 ;
        RECT 6.735000 0.550000 7.105000 1.045000 ;
      LAYER mcon ;
        RECT 0.455000 0.380000 0.625000 0.550000 ;
        RECT 0.815000 0.380000 0.985000 0.550000 ;
        RECT 1.175000 0.380000 1.345000 0.550000 ;
        RECT 1.535000 0.380000 1.705000 0.550000 ;
        RECT 1.895000 0.380000 2.065000 0.550000 ;
        RECT 2.255000 0.380000 2.425000 0.550000 ;
        RECT 2.615000 0.380000 2.785000 0.550000 ;
        RECT 2.975000 0.380000 3.145000 0.550000 ;
        RECT 3.335000 0.380000 3.505000 0.550000 ;
        RECT 3.695000 0.380000 3.865000 0.550000 ;
        RECT 4.055000 0.380000 4.225000 0.550000 ;
        RECT 4.415000 0.380000 4.585000 0.550000 ;
        RECT 4.775000 0.380000 4.945000 0.550000 ;
        RECT 5.135000 0.380000 5.305000 0.550000 ;
        RECT 5.495000 0.380000 5.665000 0.550000 ;
        RECT 5.855000 0.380000 6.025000 0.550000 ;
        RECT 6.215000 0.380000 6.385000 0.550000 ;
        RECT 6.575000 0.380000 6.745000 0.550000 ;
        RECT 6.935000 0.380000 7.105000 0.550000 ;
      LAYER met1 ;
        RECT 0.000000 0.255000 7.200000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.200000 0.085000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.115000 7.200000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 7.200000 4.155000 ;
      LAYER mcon ;
        RECT 0.155000 3.985000 0.325000 4.155000 ;
        RECT 0.635000 3.985000 0.805000 4.155000 ;
        RECT 1.115000 3.985000 1.285000 4.155000 ;
        RECT 1.595000 3.985000 1.765000 4.155000 ;
        RECT 2.075000 3.985000 2.245000 4.155000 ;
        RECT 2.555000 3.985000 2.725000 4.155000 ;
        RECT 3.035000 3.985000 3.205000 4.155000 ;
        RECT 3.515000 3.985000 3.685000 4.155000 ;
        RECT 3.995000 3.985000 4.165000 4.155000 ;
        RECT 4.475000 3.985000 4.645000 4.155000 ;
        RECT 4.955000 3.985000 5.125000 4.155000 ;
        RECT 5.435000 3.985000 5.605000 4.155000 ;
        RECT 5.915000 3.985000 6.085000 4.155000 ;
        RECT 6.395000 3.985000 6.565000 4.155000 ;
        RECT 6.875000 3.985000 7.045000 4.155000 ;
      LAYER met1 ;
        RECT 0.000000 3.955000 7.200000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095000 2.445000 0.985000 3.625000 ;
        RECT 0.095000 3.625000 7.025000 3.795000 ;
        RECT 1.775000 2.385000 2.665000 3.625000 ;
        RECT 3.335000 2.385000 4.225000 3.625000 ;
        RECT 4.895000 2.385000 5.785000 3.625000 ;
        RECT 6.455000 2.385000 7.025000 3.625000 ;
      LAYER mcon ;
        RECT 0.095000 3.475000 0.265000 3.645000 ;
        RECT 0.455000 3.475000 0.625000 3.645000 ;
        RECT 0.815000 3.475000 0.985000 3.645000 ;
        RECT 1.775000 3.475000 1.945000 3.645000 ;
        RECT 2.135000 3.475000 2.305000 3.645000 ;
        RECT 2.495000 3.475000 2.665000 3.645000 ;
        RECT 3.335000 3.475000 3.505000 3.645000 ;
        RECT 3.695000 3.475000 3.865000 3.645000 ;
        RECT 4.055000 3.475000 4.225000 3.645000 ;
        RECT 4.895000 3.475000 5.065000 3.645000 ;
        RECT 5.255000 3.475000 5.425000 3.645000 ;
        RECT 5.615000 3.475000 5.785000 3.645000 ;
        RECT 6.455000 3.475000 6.625000 3.645000 ;
        RECT 6.855000 3.475000 7.025000 3.645000 ;
      LAYER met1 ;
        RECT 0.000000 3.445000 7.200000 3.815000 ;
    END
  END VPWR
END sky130_fd_sc_hvl__inv_8
