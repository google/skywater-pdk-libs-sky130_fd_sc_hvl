# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__decap_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__decap_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.170000 0.365000 1.780000 0.845000 ;
        RECT 0.475000 0.845000 1.780000 1.250000 ;
        RECT 0.475000 1.250000 0.805000 2.030000 ;
      LAYER mcon ;
        RECT 0.215000 0.395000 0.385000 0.565000 ;
        RECT 0.655000 0.395000 0.825000 0.565000 ;
        RECT 1.095000 0.395000 1.265000 0.565000 ;
        RECT 1.510000 0.395000 1.680000 0.565000 ;
      LAYER met1 ;
        RECT 0.000000 0.255000 1.920000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 1.920000 0.085000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.115000 1.920000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 1.920000 4.155000 ;
      LAYER mcon ;
        RECT 0.155000 3.985000 0.325000 4.155000 ;
        RECT 0.635000 3.985000 0.805000 4.155000 ;
        RECT 1.115000 3.985000 1.285000 4.155000 ;
        RECT 1.595000 3.985000 1.765000 4.155000 ;
      LAYER met1 ;
        RECT 0.000000 3.955000 1.920000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.250000 2.685000 1.700000 3.755000 ;
        RECT 1.015000 1.700000 1.345000 2.685000 ;
      LAYER mcon ;
        RECT 0.495000 3.560000 0.665000 3.730000 ;
        RECT 0.860000 3.560000 1.030000 3.730000 ;
        RECT 1.300000 3.560000 1.470000 3.730000 ;
      LAYER met1 ;
        RECT 0.000000 3.445000 1.920000 3.815000 ;
    END
  END VPWR
END sky130_fd_sc_hvl__decap_4
