* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 VGND A2 a_36_113# VNB nhv w=750000u l=500000u
+  ad=2.85e+11p pd=2.26e+06u as=6.375e+11p ps=6.2e+06u
M1001 a_36_113# B2 Y VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=2.1e+11p ps=2.06e+06u
M1002 a_207_443# B1 VPWR VPB phv w=1.5e+06u l=500000u
+  ad=3.15e+11p pd=3.42e+06u as=8.55e+11p ps=7.14e+06u
M1003 Y B2 a_207_443# VPB phv w=1.5e+06u l=500000u
+  ad=5.325e+11p pd=3.71e+06u as=0p ps=0u
M1004 a_520_443# A2 Y VPB phv w=1.5e+06u l=500000u
+  ad=3.15e+11p pd=3.42e+06u as=0p ps=0u
M1005 VPWR A1 a_520_443# VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B1 a_36_113# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_36_113# A1 VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
