* File: sky130_fd_sc_hvl__dfstp_1.pxi.spice
* Created: Wed Sep  2 09:05:19 2020
* 
x_PM_SKY130_FD_SC_HVL__DFSTP_1%VNB N_VNB_M1017_b VNB N_VNB_c_2_p
+ PM_SKY130_FD_SC_HVL__DFSTP_1%VNB
x_PM_SKY130_FD_SC_HVL__DFSTP_1%VPB N_VPB_M1016_b VPB N_VPB_c_105_p
+ PM_SKY130_FD_SC_HVL__DFSTP_1%VPB
x_PM_SKY130_FD_SC_HVL__DFSTP_1%CLK N_CLK_M1016_g N_CLK_M1017_g CLK N_CLK_c_262_n
+ PM_SKY130_FD_SC_HVL__DFSTP_1%CLK
x_PM_SKY130_FD_SC_HVL__DFSTP_1%A_30_131# N_A_30_131#_M1017_s N_A_30_131#_M1016_s
+ N_A_30_131#_M1028_g N_A_30_131#_M1029_g N_A_30_131#_M1021_g
+ N_A_30_131#_c_310_n N_A_30_131#_M1014_g N_A_30_131#_M1018_g
+ N_A_30_131#_c_286_n N_A_30_131#_c_288_n N_A_30_131#_c_289_n
+ N_A_30_131#_c_290_n N_A_30_131#_c_291_n N_A_30_131#_c_293_n
+ N_A_30_131#_c_295_n N_A_30_131#_c_296_n N_A_30_131#_c_297_n
+ N_A_30_131#_c_298_n N_A_30_131#_c_317_n N_A_30_131#_c_320_n
+ N_A_30_131#_c_299_n N_A_30_131#_c_324_n N_A_30_131#_c_327_n
+ N_A_30_131#_c_330_n N_A_30_131#_c_300_n N_A_30_131#_c_332_n
+ N_A_30_131#_c_333_n N_A_30_131#_c_301_n N_A_30_131#_c_353_n
+ N_A_30_131#_c_302_n N_A_30_131#_c_335_n N_A_30_131#_c_303_n
+ N_A_30_131#_c_338_n N_A_30_131#_c_304_n N_A_30_131#_M1006_g
+ N_A_30_131#_c_340_n PM_SKY130_FD_SC_HVL__DFSTP_1%A_30_131#
x_PM_SKY130_FD_SC_HVL__DFSTP_1%D N_D_M1027_g N_D_c_525_n N_D_M1002_g D
+ PM_SKY130_FD_SC_HVL__DFSTP_1%D
x_PM_SKY130_FD_SC_HVL__DFSTP_1%A_340_593# N_A_340_593#_M1029_d
+ N_A_340_593#_M1028_d N_A_340_593#_M1024_g N_A_340_593#_M1023_g
+ N_A_340_593#_c_558_n N_A_340_593#_M1015_g N_A_340_593#_c_568_n
+ N_A_340_593#_c_571_n N_A_340_593#_c_560_n N_A_340_593#_c_575_n
+ N_A_340_593#_c_576_n N_A_340_593#_c_623_n N_A_340_593#_c_674_p
+ N_A_340_593#_c_561_n N_A_340_593#_c_562_n N_A_340_593#_c_581_n
+ N_A_340_593#_c_563_n N_A_340_593#_c_639_n N_A_340_593#_c_564_n
+ N_A_340_593#_c_642_n N_A_340_593#_c_645_n N_A_340_593#_c_583_n
+ N_A_340_593#_c_586_n N_A_340_593#_c_589_n N_A_340_593#_c_590_n
+ N_A_340_593#_c_591_n N_A_340_593#_c_565_n N_A_340_593#_c_655_n
+ N_A_340_593#_c_566_n N_A_340_593#_M1030_g
+ PM_SKY130_FD_SC_HVL__DFSTP_1%A_340_593#
x_PM_SKY130_FD_SC_HVL__DFSTP_1%A_1000_81# N_A_1000_81#_M1025_s
+ N_A_1000_81#_M1009_d N_A_1000_81#_M1003_g N_A_1000_81#_c_769_n
+ N_A_1000_81#_c_770_n N_A_1000_81#_c_771_n N_A_1000_81#_c_772_n
+ N_A_1000_81#_c_775_n N_A_1000_81#_c_777_n N_A_1000_81#_c_787_n
+ N_A_1000_81#_c_789_n N_A_1000_81#_c_791_n N_A_1000_81#_c_778_n
+ N_A_1000_81#_M1000_g PM_SKY130_FD_SC_HVL__DFSTP_1%A_1000_81#
x_PM_SKY130_FD_SC_HVL__DFSTP_1%SET_B N_SET_B_M1022_g N_SET_B_M1026_g
+ N_SET_B_c_842_n N_SET_B_c_843_n N_SET_B_M1010_g N_SET_B_c_855_n
+ N_SET_B_c_844_n N_SET_B_c_845_n N_SET_B_c_868_n N_SET_B_c_884_p SET_B SET_B
+ SET_B SET_B SET_B SET_B N_SET_B_c_847_n N_SET_B_c_892_p N_SET_B_M1020_g
+ N_SET_B_c_849_n N_SET_B_c_850_n N_SET_B_c_886_p
+ PM_SKY130_FD_SC_HVL__DFSTP_1%SET_B
x_PM_SKY130_FD_SC_HVL__DFSTP_1%A_798_107# N_A_798_107#_M1006_d
+ N_A_798_107#_M1024_d N_A_798_107#_c_935_n N_A_798_107#_M1025_g
+ N_A_798_107#_M1009_g N_A_798_107#_c_938_n N_A_798_107#_M1013_g
+ N_A_798_107#_M1011_g N_A_798_107#_c_940_n N_A_798_107#_c_951_n
+ N_A_798_107#_c_941_n N_A_798_107#_c_954_n N_A_798_107#_c_955_n
+ N_A_798_107#_c_943_n N_A_798_107#_c_944_n N_A_798_107#_c_946_n
+ N_A_798_107#_c_947_n PM_SKY130_FD_SC_HVL__DFSTP_1%A_798_107#
x_PM_SKY130_FD_SC_HVL__DFSTP_1%A_2031_177# N_A_2031_177#_M1007_d
+ N_A_2031_177#_M1012_s N_A_2031_177#_c_1055_n N_A_2031_177#_c_1060_n
+ N_A_2031_177#_c_1061_n N_A_2031_177#_c_1064_n N_A_2031_177#_c_1056_n
+ N_A_2031_177#_c_1057_n N_A_2031_177#_c_1067_n N_A_2031_177#_c_1058_n
+ N_A_2031_177#_M1019_g N_A_2031_177#_M1031_g
+ PM_SKY130_FD_SC_HVL__DFSTP_1%A_2031_177#
x_PM_SKY130_FD_SC_HVL__DFSTP_1%A_1787_137# N_A_1787_137#_M1015_d
+ N_A_1787_137#_M1014_d N_A_1787_137#_M1010_d N_A_1787_137#_M1007_g
+ N_A_1787_137#_M1012_g N_A_1787_137#_c_1133_n N_A_1787_137#_M1004_g
+ N_A_1787_137#_c_1135_n N_A_1787_137#_M1005_g N_A_1787_137#_c_1138_n
+ N_A_1787_137#_c_1139_n N_A_1787_137#_c_1142_n N_A_1787_137#_c_1131_n
+ N_A_1787_137#_c_1143_n N_A_1787_137#_c_1144_n N_A_1787_137#_c_1155_n
+ N_A_1787_137#_c_1145_n N_A_1787_137#_c_1146_n N_A_1787_137#_c_1147_n
+ N_A_1787_137#_c_1148_n PM_SKY130_FD_SC_HVL__DFSTP_1%A_1787_137#
x_PM_SKY130_FD_SC_HVL__DFSTP_1%A_2553_203# N_A_2553_203#_M1004_s
+ N_A_2553_203#_M1005_s N_A_2553_203#_M1008_g N_A_2553_203#_M1001_g
+ N_A_2553_203#_c_1256_n N_A_2553_203#_c_1264_n N_A_2553_203#_c_1257_n
+ N_A_2553_203#_c_1258_n N_A_2553_203#_c_1266_n N_A_2553_203#_c_1268_n
+ N_A_2553_203#_c_1290_n N_A_2553_203#_c_1259_n N_A_2553_203#_c_1260_n
+ N_A_2553_203#_c_1276_n PM_SKY130_FD_SC_HVL__DFSTP_1%A_2553_203#
x_PM_SKY130_FD_SC_HVL__DFSTP_1%VPWR N_VPWR_M1016_d N_VPWR_M1002_s N_VPWR_M1000_d
+ N_VPWR_M1026_d N_VPWR_M1031_d N_VPWR_M1012_d N_VPWR_M1005_d VPWR
+ N_VPWR_c_1317_n N_VPWR_c_1320_n N_VPWR_c_1323_n N_VPWR_c_1326_n
+ N_VPWR_c_1329_n N_VPWR_c_1332_n N_VPWR_c_1335_n N_VPWR_c_1338_n
+ PM_SKY130_FD_SC_HVL__DFSTP_1%VPWR
x_PM_SKY130_FD_SC_HVL__DFSTP_1%A_642_107# N_A_642_107#_M1027_d
+ N_A_642_107#_M1002_d N_A_642_107#_c_1438_n N_A_642_107#_c_1439_n
+ PM_SKY130_FD_SC_HVL__DFSTP_1%A_642_107#
x_PM_SKY130_FD_SC_HVL__DFSTP_1%Q N_Q_M1008_d N_Q_M1001_d Q Q Q Q Q Q Q
+ N_Q_c_1461_n PM_SKY130_FD_SC_HVL__DFSTP_1%Q
x_PM_SKY130_FD_SC_HVL__DFSTP_1%VGND N_VGND_M1017_d N_VGND_M1027_s N_VGND_M1003_d
+ N_VGND_M1022_d N_VGND_M1020_d N_VGND_M1004_d VGND N_VGND_c_1476_n
+ N_VGND_c_1478_n N_VGND_c_1480_n N_VGND_c_1482_n N_VGND_c_1484_n
+ N_VGND_c_1486_n N_VGND_c_1488_n PM_SKY130_FD_SC_HVL__DFSTP_1%VGND
cc_1 N_VNB_M1017_b N_CLK_M1017_g 0.107853f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=0.865
cc_2 N_VNB_c_2_p N_CLK_M1017_g 5.52994e-19 $X=0.24 $Y=0 $X2=0.685 $Y2=0.865
cc_3 N_VNB_M1017_b N_A_30_131#_M1029_g 0.0451994f $X=-0.33 $Y=-0.265 $X2=0.71
+ $Y2=2.24
cc_4 N_VNB_c_2_p N_A_30_131#_M1029_g 5.14587e-19 $X=0.24 $Y=0 $X2=0.71 $Y2=2.24
cc_5 N_VNB_M1017_b N_A_30_131#_M1018_g 0.0587138f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_M1017_b N_A_30_131#_c_286_n 0.0361636f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_7 N_VNB_c_2_p N_A_30_131#_c_286_n 5.2203e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_8 N_VNB_M1017_b N_A_30_131#_c_288_n 0.022226f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_M1017_b N_A_30_131#_c_289_n 0.0132081f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_10 N_VNB_M1017_b N_A_30_131#_c_290_n 0.00110658f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1017_b N_A_30_131#_c_291_n 0.0656548f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_c_2_p N_A_30_131#_c_291_n 0.00262311f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_13 N_VNB_M1017_b N_A_30_131#_c_293_n 0.0141601f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_c_2_p N_A_30_131#_c_293_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_15 N_VNB_M1017_b N_A_30_131#_c_295_n 0.0154161f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_16 N_VNB_M1017_b N_A_30_131#_c_296_n 0.011832f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_17 N_VNB_M1017_b N_A_30_131#_c_297_n 0.00919848f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1017_b N_A_30_131#_c_298_n 0.00168577f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_19 N_VNB_M1017_b N_A_30_131#_c_299_n 0.00171491f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_20 N_VNB_M1017_b N_A_30_131#_c_300_n 0.00206039f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_21 N_VNB_M1017_b N_A_30_131#_c_301_n 0.00841486f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_22 N_VNB_M1017_b N_A_30_131#_c_302_n 0.0726517f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_23 N_VNB_M1017_b N_A_30_131#_c_303_n 0.00132349f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_24 N_VNB_M1017_b N_A_30_131#_c_304_n 0.0269613f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_25 N_VNB_M1017_b N_A_30_131#_M1006_g 0.119559f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_26 N_VNB_c_2_p N_A_30_131#_M1006_g 0.0023273f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_27 N_VNB_M1017_b N_D_M1027_g 0.0679612f $X=-0.33 $Y=-0.265 $X2=0.67 $Y2=3.34
cc_28 N_VNB_c_2_p N_D_M1027_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.67 $Y2=3.34
cc_29 N_VNB_M1017_b N_D_c_525_n 0.082187f $X=-0.33 $Y=-0.265 $X2=0.685 $Y2=1.95
cc_30 N_VNB_M1017_b N_A_340_593#_M1023_g 0.0830299f $X=-0.33 $Y=-0.265 $X2=0.71
+ $Y2=2.24
cc_31 N_VNB_c_2_p N_A_340_593#_M1023_g 0.0023273f $X=0.24 $Y=0 $X2=0.71 $Y2=2.24
cc_32 N_VNB_M1017_b N_A_340_593#_c_558_n 0.0782083f $X=-0.33 $Y=-0.265 $X2=0.677
+ $Y2=2.45
cc_33 N_VNB_c_2_p N_A_340_593#_c_558_n 0.00196852f $X=0.24 $Y=0 $X2=0.677
+ $Y2=2.45
cc_34 N_VNB_M1017_b N_A_340_593#_c_560_n 0.0116605f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_35 N_VNB_M1017_b N_A_340_593#_c_561_n 0.0420074f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_36 N_VNB_M1017_b N_A_340_593#_c_562_n 0.0210183f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_37 N_VNB_M1017_b N_A_340_593#_c_563_n 0.00479192f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_38 N_VNB_M1017_b N_A_340_593#_c_564_n 0.00936135f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_39 N_VNB_M1017_b N_A_340_593#_c_565_n 0.00301816f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_M1017_b N_A_340_593#_c_566_n 0.00223646f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_41 N_VNB_M1017_b N_A_1000_81#_M1003_g 0.0654634f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=2.32
cc_42 N_VNB_M1017_b N_A_1000_81#_c_769_n 0.016635f $X=-0.33 $Y=-0.265 $X2=0.71
+ $Y2=2.24
cc_43 N_VNB_M1017_b N_A_1000_81#_c_770_n 0.026493f $X=-0.33 $Y=-0.265 $X2=0.677
+ $Y2=1.95
cc_44 N_VNB_M1017_b N_A_1000_81#_c_771_n 0.024696f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_45 N_VNB_M1017_b N_A_1000_81#_c_772_n 0.00123723f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_M1017_b N_SET_B_M1026_g 0.00959969f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=0.865
cc_47 N_VNB_M1017_b N_SET_B_c_842_n 0.026363f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_48 N_VNB_M1017_b N_SET_B_c_843_n 0.00320809f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=2.32
cc_49 N_VNB_M1017_b N_SET_B_c_844_n 0.0039534f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_50 N_VNB_M1017_b N_SET_B_c_845_n 0.0508166f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_51 N_VNB_M1017_b SET_B 0.0383962f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_52 N_VNB_M1017_b N_SET_B_c_847_n 0.100674f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_53 N_VNB_c_2_p N_SET_B_c_847_n 0.00221559f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_54 N_VNB_M1017_b N_SET_B_c_849_n 0.0301704f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_55 N_VNB_M1017_b N_SET_B_c_850_n 0.0661431f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_56 N_VNB_c_2_p N_SET_B_c_850_n 0.00779379f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_57 N_VNB_M1017_b N_A_798_107#_c_935_n 0.134293f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=0.865
cc_58 N_VNB_c_2_p N_A_798_107#_c_935_n 0.0456632f $X=0.24 $Y=0 $X2=0.685
+ $Y2=0.865
cc_59 N_VNB_M1017_b N_A_798_107#_M1025_g 0.0753615f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_60 N_VNB_M1017_b N_A_798_107#_c_938_n 0.1786f $X=-0.33 $Y=-0.265 $X2=0.677
+ $Y2=2.45
cc_61 N_VNB_M1017_b N_A_798_107#_M1013_g 0.048566f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_62 N_VNB_M1017_b N_A_798_107#_c_940_n 0.0651255f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_63 N_VNB_M1017_b N_A_798_107#_c_941_n 0.00892207f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_64 N_VNB_c_2_p N_A_798_107#_c_941_n 6.3194e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_65 N_VNB_M1017_b N_A_798_107#_c_943_n 0.011738f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_66 N_VNB_M1017_b N_A_798_107#_c_944_n 0.0208715f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_67 N_VNB_c_2_p N_A_798_107#_c_944_n 0.00157832f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_68 N_VNB_M1017_b N_A_798_107#_c_946_n 0.00237943f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_69 N_VNB_M1017_b N_A_798_107#_c_947_n 0.00814527f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_70 N_VNB_M1017_b N_A_2031_177#_c_1055_n 0.0114464f $X=-0.33 $Y=-0.265
+ $X2=0.685 $Y2=0.865
cc_71 N_VNB_M1017_b N_A_2031_177#_c_1056_n 0.0128128f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_72 N_VNB_M1017_b N_A_2031_177#_c_1057_n 0.00111476f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_73 N_VNB_M1017_b N_A_2031_177#_c_1058_n 0.0106953f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_74 N_VNB_M1017_b N_A_2031_177#_M1019_g 0.0618424f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_75 N_VNB_M1017_b N_A_1787_137#_M1007_g 0.0742443f $X=-0.33 $Y=-0.265 $X2=0.71
+ $Y2=2.24
cc_76 N_VNB_M1017_b N_A_1787_137#_M1004_g 0.078102f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_77 N_VNB_M1017_b N_A_1787_137#_c_1131_n 0.00433734f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_78 N_VNB_M1017_b N_A_2553_203#_M1008_g 0.0490494f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=2.32
cc_79 N_VNB_c_2_p N_A_2553_203#_M1008_g 9.48828e-19 $X=0.24 $Y=0 $X2=0.635
+ $Y2=2.32
cc_80 N_VNB_M1017_b N_A_2553_203#_c_1256_n 0.0340466f $X=-0.33 $Y=-0.265
+ $X2=0.677 $Y2=2.45
cc_81 N_VNB_M1017_b N_A_2553_203#_c_1257_n 0.00823078f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_82 N_VNB_M1017_b N_A_2553_203#_c_1258_n 0.005082f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_83 N_VNB_M1017_b N_A_2553_203#_c_1259_n 0.00357789f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_84 N_VNB_M1017_b N_A_2553_203#_c_1260_n 0.00354733f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_85 N_VNB_M1017_b N_A_642_107#_c_1438_n 0.00716869f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=2.32
cc_86 N_VNB_M1017_b N_A_642_107#_c_1439_n 0.0175182f $X=-0.33 $Y=-0.265 $X2=0.71
+ $Y2=2.24
cc_87 N_VNB_c_2_p N_A_642_107#_c_1439_n 9.59404e-19 $X=0.24 $Y=0 $X2=0.71
+ $Y2=2.24
cc_88 N_VNB_M1017_b N_Q_c_1461_n 0.0589273f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_89 N_VNB_M1017_b N_VGND_c_1476_n 0.0346157f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_90 N_VNB_c_2_p N_VGND_c_1476_n 0.00166879f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_91 N_VNB_M1017_b N_VGND_c_1478_n 0.0294265f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_92 N_VNB_c_2_p N_VGND_c_1478_n 0.00151451f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_93 N_VNB_M1017_b N_VGND_c_1480_n 0.0510207f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_94 N_VNB_c_2_p N_VGND_c_1480_n 0.00271305f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_95 N_VNB_M1017_b N_VGND_c_1482_n 0.0419228f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_96 N_VNB_c_2_p N_VGND_c_1482_n 0.00449559f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_97 N_VNB_M1017_b N_VGND_c_1484_n 0.0500643f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_98 N_VNB_c_2_p N_VGND_c_1484_n 0.00166879f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_99 N_VNB_M1017_b N_VGND_c_1486_n 0.0822184f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_100 N_VNB_c_2_p N_VGND_c_1486_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_101 N_VNB_M1017_b N_VGND_c_1488_n 0.246678f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_102 N_VNB_c_2_p N_VGND_c_1488_n 1.58776f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_103 N_VPB_M1016_b N_CLK_M1016_g 0.0762003f $X=-0.33 $Y=1.885 $X2=0.67
+ $Y2=3.34
cc_104 VPB N_CLK_M1016_g 0.00970178f $X=0 $Y=3.955 $X2=0.67 $Y2=3.34
cc_105 N_VPB_c_105_p N_CLK_M1016_g 0.0152133f $X=14.64 $Y=4.07 $X2=0.67 $Y2=3.34
cc_106 N_VPB_M1016_b N_CLK_M1017_g 0.00606517f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=0.865
cc_107 N_VPB_M1016_b N_CLK_c_262_n 0.0500026f $X=-0.33 $Y=1.885 $X2=0.71
+ $Y2=2.24
cc_108 N_VPB_M1016_b N_A_30_131#_M1028_g 0.128625f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=2.32
cc_109 VPB N_A_30_131#_M1028_g 0.00970178f $X=0 $Y=3.955 $X2=0.635 $Y2=2.32
cc_110 N_VPB_c_105_p N_A_30_131#_M1028_g 0.015886f $X=14.64 $Y=4.07 $X2=0.635
+ $Y2=2.32
cc_111 N_VPB_M1016_b N_A_30_131#_c_310_n 0.0365205f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=2.41
cc_112 VPB N_A_30_131#_c_310_n 0.00109097f $X=0 $Y=3.955 $X2=0.72 $Y2=2.41
cc_113 N_VPB_c_105_p N_A_30_131#_c_310_n 0.00680566f $X=14.64 $Y=4.07 $X2=0.72
+ $Y2=2.41
cc_114 N_VPB_M1016_b N_A_30_131#_c_288_n 0.0800752f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_115 VPB N_A_30_131#_c_288_n 7.36921e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_116 N_VPB_c_105_p N_A_30_131#_c_288_n 0.0120479f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_117 N_VPB_M1016_b N_A_30_131#_c_298_n 0.00393926f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_118 N_VPB_M1016_b N_A_30_131#_c_317_n 0.00699855f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_119 VPB N_A_30_131#_c_317_n 0.00223977f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_120 N_VPB_c_105_p N_A_30_131#_c_317_n 0.0146189f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_121 N_VPB_M1016_b N_A_30_131#_c_320_n 0.00114907f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_122 VPB N_A_30_131#_c_320_n 7.77907e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_123 N_VPB_c_105_p N_A_30_131#_c_320_n 0.00472626f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_124 N_VPB_M1016_b N_A_30_131#_c_299_n 0.00234604f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_125 N_VPB_M1016_b N_A_30_131#_c_324_n 0.00714348f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_126 VPB N_A_30_131#_c_324_n 0.00409757f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_127 N_VPB_c_105_p N_A_30_131#_c_324_n 0.0324095f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_128 N_VPB_M1016_b N_A_30_131#_c_327_n 0.0600418f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_129 VPB N_A_30_131#_c_327_n 0.00249404f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_130 N_VPB_c_105_p N_A_30_131#_c_327_n 0.00802262f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_131 N_VPB_M1016_b N_A_30_131#_c_330_n 0.00618221f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_132 N_VPB_M1016_b N_A_30_131#_c_300_n 0.00680814f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_133 N_VPB_M1016_b N_A_30_131#_c_332_n 0.00415379f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_134 N_VPB_M1016_b N_A_30_131#_c_333_n 0.0208985f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_135 N_VPB_M1016_b N_A_30_131#_c_302_n 0.00946949f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_136 VPB N_A_30_131#_c_335_n 7.77907e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_137 N_VPB_c_105_p N_A_30_131#_c_335_n 0.00472626f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_138 N_VPB_M1016_b N_A_30_131#_c_303_n 0.00156775f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_139 N_VPB_M1016_b N_A_30_131#_c_338_n 0.00243944f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_140 N_VPB_M1016_b N_A_30_131#_c_304_n 0.119203f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_141 N_VPB_M1016_b N_A_30_131#_c_340_n 0.0318185f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_142 N_VPB_M1016_b N_D_c_525_n 0.104197f $X=-0.33 $Y=1.885 $X2=0.685 $Y2=1.95
cc_143 N_VPB_M1016_b N_D_M1002_g 0.0332879f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=0.865
cc_144 N_VPB_M1016_b N_A_340_593#_M1024_g 0.0419988f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_145 N_VPB_M1016_b N_A_340_593#_c_568_n 0.174029f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=2.41
cc_146 VPB N_A_340_593#_c_568_n 0.0287467f $X=0 $Y=3.955 $X2=0.72 $Y2=2.41
cc_147 N_VPB_c_105_p N_A_340_593#_c_568_n 0.0481497f $X=14.64 $Y=4.07 $X2=0.72
+ $Y2=2.41
cc_148 N_VPB_M1016_b N_A_340_593#_c_571_n 0.00924525f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_149 VPB N_A_340_593#_c_571_n 0.00101808f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_150 N_VPB_c_105_p N_A_340_593#_c_571_n 0.0158392f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_151 N_VPB_M1016_b N_A_340_593#_c_560_n 0.00566483f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_152 N_VPB_M1016_b N_A_340_593#_c_575_n 0.0285328f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_153 N_VPB_M1016_b N_A_340_593#_c_576_n 0.00699264f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_154 VPB N_A_340_593#_c_576_n 8.06243e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_155 N_VPB_c_105_p N_A_340_593#_c_576_n 0.00821266f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_156 N_VPB_M1016_b N_A_340_593#_c_561_n 0.115025f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_157 N_VPB_M1016_b N_A_340_593#_c_562_n 0.00311247f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_158 N_VPB_M1016_b N_A_340_593#_c_581_n 0.00774819f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_159 N_VPB_M1016_b N_A_340_593#_c_563_n 0.00578113f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_160 N_VPB_M1016_b N_A_340_593#_c_583_n 0.00189949f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_161 VPB N_A_340_593#_c_583_n 5.70856e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_162 N_VPB_c_105_p N_A_340_593#_c_583_n 0.0114989f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_163 N_VPB_M1016_b N_A_340_593#_c_586_n 0.00526822f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_164 VPB N_A_340_593#_c_586_n 0.00363331f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_165 N_VPB_c_105_p N_A_340_593#_c_586_n 0.0621681f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_166 N_VPB_M1016_b N_A_340_593#_c_589_n 0.00368911f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_167 N_VPB_M1016_b N_A_340_593#_c_590_n 0.00798422f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_168 N_VPB_M1016_b N_A_340_593#_c_591_n 0.00343325f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_169 N_VPB_M1016_b N_A_340_593#_M1030_g 0.121574f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_170 VPB N_A_340_593#_M1030_g 0.00983156f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_171 N_VPB_c_105_p N_A_340_593#_M1030_g 0.0153362f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_172 N_VPB_M1016_b N_A_1000_81#_c_769_n 0.00877413f $X=-0.33 $Y=1.885 $X2=0.71
+ $Y2=2.24
cc_173 N_VPB_M1016_b N_A_1000_81#_c_770_n 0.00314481f $X=-0.33 $Y=1.885
+ $X2=0.677 $Y2=1.95
cc_174 VPB N_A_1000_81#_c_775_n 0.00105511f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_175 N_VPB_c_105_p N_A_1000_81#_c_775_n 0.00534802f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_176 N_VPB_M1016_b N_A_1000_81#_c_777_n 0.00206039f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_177 N_VPB_M1016_b N_A_1000_81#_c_778_n 0.00416532f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_178 N_VPB_M1016_b N_A_1000_81#_M1000_g 0.107439f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_179 VPB N_A_1000_81#_M1000_g 0.00228906f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_180 N_VPB_c_105_p N_A_1000_81#_M1000_g 0.00956687f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_181 N_VPB_M1016_b N_SET_B_M1026_g 0.0722637f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=0.865
cc_182 N_VPB_M1016_b N_SET_B_c_843_n 0.0258514f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=2.32
cc_183 N_VPB_M1016_b N_SET_B_M1010_g 0.039574f $X=-0.33 $Y=1.885 $X2=0.71
+ $Y2=2.24
cc_184 N_VPB_M1016_b N_SET_B_c_855_n 0.0271489f $X=-0.33 $Y=1.885 $X2=0.71
+ $Y2=2.41
cc_185 N_VPB_M1016_b N_SET_B_c_845_n 0.0122535f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_186 N_VPB_M1016_b N_A_798_107#_M1009_g 0.0441707f $X=-0.33 $Y=1.885 $X2=0.71
+ $Y2=2.24
cc_187 N_VPB_M1016_b N_A_798_107#_M1013_g 0.018704f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_188 N_VPB_M1016_b N_A_798_107#_c_940_n 0.0364677f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_189 N_VPB_M1016_b N_A_798_107#_c_951_n 0.0739074f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_190 VPB N_A_798_107#_c_951_n 0.00117695f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_191 N_VPB_c_105_p N_A_798_107#_c_951_n 0.00737898f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_192 N_VPB_M1016_b N_A_798_107#_c_954_n 0.00240186f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_193 N_VPB_M1016_b N_A_798_107#_c_955_n 0.00300364f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_194 N_VPB_M1016_b N_A_798_107#_c_947_n 0.00669708f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_195 N_VPB_M1016_b N_A_2031_177#_c_1060_n 0.00647095f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=2.32
cc_196 N_VPB_M1016_b N_A_2031_177#_c_1061_n 0.00504927f $X=-0.33 $Y=1.885
+ $X2=0.677 $Y2=2.24
cc_197 VPB N_A_2031_177#_c_1061_n 7.61228e-19 $X=0 $Y=3.955 $X2=0.677 $Y2=2.24
cc_198 N_VPB_c_105_p N_A_2031_177#_c_1061_n 0.0130842f $X=14.64 $Y=4.07
+ $X2=0.677 $Y2=2.24
cc_199 N_VPB_M1016_b N_A_2031_177#_c_1064_n 0.0114864f $X=-0.33 $Y=1.885
+ $X2=0.71 $Y2=2.24
cc_200 N_VPB_M1016_b N_A_2031_177#_c_1057_n 0.0122649f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_201 N_VPB_M1016_b N_A_2031_177#_M1019_g 0.0857562f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_202 N_VPB_M1016_b N_A_1787_137#_M1007_g 0.00954856f $X=-0.33 $Y=1.885
+ $X2=0.71 $Y2=2.24
cc_203 N_VPB_M1016_b N_A_1787_137#_c_1133_n 0.0887975f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_204 N_VPB_M1016_b N_A_1787_137#_M1004_g 0.0102558f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_205 N_VPB_M1016_b N_A_1787_137#_c_1135_n 0.0396135f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_206 VPB N_A_1787_137#_c_1135_n 7.77452e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_207 N_VPB_c_105_p N_A_1787_137#_c_1135_n 0.00424836f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_208 N_VPB_M1016_b N_A_1787_137#_c_1138_n 0.0460947f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_209 N_VPB_M1016_b N_A_1787_137#_c_1139_n 0.0670309f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_210 VPB N_A_1787_137#_c_1139_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_211 N_VPB_c_105_p N_A_1787_137#_c_1139_n 0.0138108f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_212 N_VPB_M1016_b N_A_1787_137#_c_1142_n 0.0392751f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_213 N_VPB_M1016_b N_A_1787_137#_c_1143_n 0.00499359f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_214 N_VPB_M1016_b N_A_1787_137#_c_1144_n 0.00151296f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_215 N_VPB_M1016_b N_A_1787_137#_c_1145_n 0.0190576f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_216 N_VPB_M1016_b N_A_1787_137#_c_1146_n 8.47737e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_217 N_VPB_M1016_b N_A_1787_137#_c_1147_n 0.047392f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_218 N_VPB_M1016_b N_A_1787_137#_c_1148_n 0.00522035f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_219 N_VPB_M1016_b N_A_2553_203#_M1001_g 0.0452815f $X=-0.33 $Y=1.885 $X2=0.71
+ $Y2=2.24
cc_220 VPB N_A_2553_203#_M1001_g 0.00250311f $X=0 $Y=3.955 $X2=0.71 $Y2=2.24
cc_221 N_VPB_c_105_p N_A_2553_203#_M1001_g 0.00978839f $X=14.64 $Y=4.07 $X2=0.71
+ $Y2=2.24
cc_222 N_VPB_M1016_b N_A_2553_203#_c_1264_n 0.0324487f $X=-0.33 $Y=1.885
+ $X2=0.72 $Y2=2.41
cc_223 N_VPB_M1016_b N_A_2553_203#_c_1258_n 0.00115485f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_224 N_VPB_M1016_b N_A_2553_203#_c_1266_n 0.0039009f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_225 N_VPB_c_105_p N_A_2553_203#_c_1266_n 0.00327732f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_226 N_VPB_M1016_b N_A_2553_203#_c_1268_n 0.0131103f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_227 N_VPB_M1016_b N_A_2553_203#_c_1259_n 0.0323565f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_228 N_VPB_M1016_b N_VPWR_c_1317_n 0.0122659f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1317_n 0.00406397f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_230 N_VPB_c_105_p N_VPWR_c_1317_n 0.047451f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_231 N_VPB_M1016_b N_VPWR_c_1320_n 0.0222993f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1320_n 7.03841e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_233 N_VPB_c_105_p N_VPWR_c_1320_n 0.0107249f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_234 N_VPB_M1016_b N_VPWR_c_1323_n 0.0192629f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1323_n 9.30887e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_236 N_VPB_c_105_p N_VPWR_c_1323_n 0.0141846f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_237 N_VPB_M1016_b N_VPWR_c_1326_n 0.0239632f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1326_n 0.00318418f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_239 N_VPB_c_105_p N_VPWR_c_1326_n 0.0399652f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_240 N_VPB_M1016_b N_VPWR_c_1329_n 0.030607f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1329_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_242 N_VPB_c_105_p N_VPWR_c_1329_n 0.0409968f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_243 N_VPB_M1016_b N_VPWR_c_1332_n 0.0128579f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1332_n 0.00361638f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_245 N_VPB_c_105_p N_VPWR_c_1332_n 0.0437252f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_246 N_VPB_M1016_b N_VPWR_c_1335_n 0.00983222f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1335_n 0.00319858f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_248 N_VPB_c_105_p N_VPWR_c_1335_n 0.0396892f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_249 N_VPB_M1016_b N_VPWR_c_1338_n 0.146979f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1338_n 1.5855f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_251 N_VPB_c_105_p N_VPWR_c_1338_n 0.0729226f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_252 N_VPB_M1016_b N_A_642_107#_c_1438_n 0.0155615f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=2.32
cc_253 N_VPB_M1016_b N_Q_c_1461_n 0.0675129f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_254 VPB N_Q_c_1461_n 9.56025e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_255 N_VPB_c_105_p N_Q_c_1461_n 0.0108986f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_256 N_CLK_M1016_g N_A_30_131#_M1028_g 0.0404347f $X=0.67 $Y=3.34 $X2=0 $Y2=0
cc_257 CLK N_A_30_131#_M1028_g 0.00427882f $X=0.635 $Y=2.32 $X2=0 $Y2=0
cc_258 N_CLK_c_262_n N_A_30_131#_M1028_g 0.0294745f $X=0.71 $Y=2.24 $X2=0 $Y2=0
cc_259 N_CLK_M1017_g N_A_30_131#_M1029_g 0.01416f $X=0.685 $Y=0.865 $X2=0 $Y2=0
cc_260 N_CLK_M1017_g N_A_30_131#_c_286_n 0.0114062f $X=0.685 $Y=0.865 $X2=0
+ $Y2=0
cc_261 N_CLK_M1017_g N_A_30_131#_c_288_n 0.0222295f $X=0.685 $Y=0.865 $X2=0
+ $Y2=0
cc_262 CLK N_A_30_131#_c_288_n 0.04973f $X=0.635 $Y=2.32 $X2=0 $Y2=0
cc_263 N_CLK_c_262_n N_A_30_131#_c_288_n 0.0370442f $X=0.71 $Y=2.24 $X2=0 $Y2=0
cc_264 N_CLK_M1017_g N_A_30_131#_c_289_n 0.0407169f $X=0.685 $Y=0.865 $X2=0
+ $Y2=0
cc_265 CLK N_A_30_131#_c_289_n 0.00866996f $X=0.635 $Y=2.32 $X2=0 $Y2=0
cc_266 N_CLK_c_262_n N_A_30_131#_c_289_n 4.47249e-19 $X=0.71 $Y=2.24 $X2=0 $Y2=0
cc_267 N_CLK_M1017_g N_A_30_131#_c_290_n 0.0012582f $X=0.685 $Y=0.865 $X2=0
+ $Y2=0
cc_268 N_CLK_M1017_g N_A_30_131#_c_353_n 0.00300946f $X=0.685 $Y=0.865 $X2=0
+ $Y2=0
cc_269 N_CLK_M1017_g N_A_30_131#_c_302_n 0.0497206f $X=0.685 $Y=0.865 $X2=0
+ $Y2=0
cc_270 N_CLK_M1016_g N_VPWR_c_1317_n 0.0466884f $X=0.67 $Y=3.34 $X2=0 $Y2=0
cc_271 CLK N_VPWR_c_1317_n 0.0264328f $X=0.635 $Y=2.32 $X2=0 $Y2=0
cc_272 N_CLK_c_262_n N_VPWR_c_1317_n 5.26683e-19 $X=0.71 $Y=2.24 $X2=0 $Y2=0
cc_273 N_CLK_M1016_g N_VPWR_c_1338_n 0.00853624f $X=0.67 $Y=3.34 $X2=0 $Y2=0
cc_274 N_CLK_M1017_g N_VGND_c_1476_n 0.0401717f $X=0.685 $Y=0.865 $X2=0 $Y2=0
cc_275 N_CLK_M1017_g N_VGND_c_1488_n 0.00911864f $X=0.685 $Y=0.865 $X2=0 $Y2=0
cc_276 N_A_30_131#_c_295_n N_D_M1027_g 0.00661619f $X=2.205 $Y=1.175 $X2=0 $Y2=0
cc_277 N_A_30_131#_c_296_n N_D_M1027_g 0.0176119f $X=3.015 $Y=1.26 $X2=0 $Y2=0
cc_278 N_A_30_131#_M1006_g N_D_M1027_g 0.0448742f $X=3.74 $Y=0.745 $X2=0 $Y2=0
cc_279 N_A_30_131#_c_296_n N_D_c_525_n 0.021192f $X=3.015 $Y=1.26 $X2=-0.33
+ $Y2=-0.265
cc_280 N_A_30_131#_c_298_n N_D_c_525_n 0.0492454f $X=3.1 $Y=3.285 $X2=-0.33
+ $Y2=-0.265
cc_281 N_A_30_131#_c_298_n N_D_M1002_g 0.0280422f $X=3.1 $Y=3.285 $X2=0 $Y2=0
cc_282 N_A_30_131#_c_317_n N_D_M1002_g 0.00327289f $X=3.715 $Y=3.45 $X2=0 $Y2=0
cc_283 N_A_30_131#_c_299_n N_D_M1002_g 6.51992e-19 $X=3.8 $Y=1.25 $X2=0 $Y2=0
cc_284 N_A_30_131#_c_296_n D 0.02351f $X=3.015 $Y=1.26 $X2=0 $Y2=0
cc_285 N_A_30_131#_c_298_n D 0.0397145f $X=3.1 $Y=3.285 $X2=0 $Y2=0
cc_286 N_A_30_131#_c_298_n N_A_340_593#_M1024_g 0.00255985f $X=3.1 $Y=3.285
+ $X2=0.24 $Y2=0
cc_287 N_A_30_131#_c_317_n N_A_340_593#_M1024_g 0.0100258f $X=3.715 $Y=3.45
+ $X2=0.24 $Y2=0
cc_288 N_A_30_131#_c_299_n N_A_340_593#_M1024_g 0.0300556f $X=3.8 $Y=1.25
+ $X2=0.24 $Y2=0
cc_289 N_A_30_131#_c_324_n N_A_340_593#_M1024_g 0.0126546f $X=4.835 $Y=3.45
+ $X2=0.24 $Y2=0
cc_290 N_A_30_131#_c_327_n N_A_340_593#_M1024_g 0.023367f $X=4.565 $Y=3.45
+ $X2=0.24 $Y2=0
cc_291 N_A_30_131#_c_335_n N_A_340_593#_M1024_g 0.00190495f $X=3.8 $Y=3.45
+ $X2=0.24 $Y2=0
cc_292 N_A_30_131#_c_340_n N_A_340_593#_M1024_g 0.00996342f $X=4.645 $Y=3.175
+ $X2=0.24 $Y2=0
cc_293 N_A_30_131#_M1006_g N_A_340_593#_M1023_g 0.027534f $X=3.74 $Y=0.745 $X2=0
+ $Y2=0
cc_294 N_A_30_131#_M1018_g N_A_340_593#_c_558_n 0.0190146f $X=9.695 $Y=1.225
+ $X2=0 $Y2=0
cc_295 N_A_30_131#_c_333_n N_A_340_593#_c_558_n 0.00104755f $X=8.63 $Y=2.41
+ $X2=0 $Y2=0
cc_296 N_A_30_131#_c_338_n N_A_340_593#_c_558_n 6.22195e-19 $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_297 N_A_30_131#_c_304_n N_A_340_593#_c_558_n 0.0307035f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_298 N_A_30_131#_c_317_n N_A_340_593#_c_568_n 0.0221786f $X=3.715 $Y=3.45
+ $X2=0 $Y2=0
cc_299 N_A_30_131#_c_320_n N_A_340_593#_c_568_n 0.00896514f $X=3.185 $Y=3.45
+ $X2=0 $Y2=0
cc_300 N_A_30_131#_c_324_n N_A_340_593#_c_568_n 0.00912415f $X=4.835 $Y=3.45
+ $X2=0 $Y2=0
cc_301 N_A_30_131#_c_335_n N_A_340_593#_c_568_n 0.00546828f $X=3.8 $Y=3.45 $X2=0
+ $Y2=0
cc_302 N_A_30_131#_M1028_g N_A_340_593#_c_571_n 0.0143195f $X=1.45 $Y=3.34
+ $X2=7.44 $Y2=0
cc_303 N_A_30_131#_M1028_g N_A_340_593#_c_560_n 0.0205072f $X=1.45 $Y=3.34 $X2=0
+ $Y2=0
cc_304 N_A_30_131#_M1029_g N_A_340_593#_c_560_n 0.013512f $X=1.465 $Y=0.865
+ $X2=0 $Y2=0
cc_305 N_A_30_131#_c_290_n N_A_340_593#_c_560_n 0.0452134f $X=1.425 $Y=1.295
+ $X2=0 $Y2=0
cc_306 N_A_30_131#_c_291_n N_A_340_593#_c_560_n 0.0168914f $X=2.12 $Y=0.35 $X2=0
+ $Y2=0
cc_307 N_A_30_131#_c_295_n N_A_340_593#_c_560_n 0.0409957f $X=2.205 $Y=1.175
+ $X2=0 $Y2=0
cc_308 N_A_30_131#_c_297_n N_A_340_593#_c_560_n 0.0141596f $X=2.29 $Y=1.26 $X2=0
+ $Y2=0
cc_309 N_A_30_131#_c_353_n N_A_340_593#_c_560_n 0.0428495f $X=1.345 $Y=1.425
+ $X2=0 $Y2=0
cc_310 N_A_30_131#_c_302_n N_A_340_593#_c_560_n 0.028362f $X=1.345 $Y=1.425
+ $X2=0 $Y2=0
cc_311 N_A_30_131#_c_298_n N_A_340_593#_c_575_n 0.0123662f $X=3.1 $Y=3.285 $X2=0
+ $Y2=0
cc_312 N_A_30_131#_c_298_n N_A_340_593#_c_576_n 0.054934f $X=3.1 $Y=3.285 $X2=0
+ $Y2=0
cc_313 N_A_30_131#_c_320_n N_A_340_593#_c_576_n 0.0231191f $X=3.185 $Y=3.45
+ $X2=0 $Y2=0
cc_314 N_A_30_131#_c_332_n N_A_340_593#_c_623_n 7.9431e-19 $X=5.005 $Y=2.24
+ $X2=0 $Y2=0
cc_315 N_A_30_131#_c_340_n N_A_340_593#_c_623_n 0.0015369f $X=4.645 $Y=3.175
+ $X2=0 $Y2=0
cc_316 N_A_30_131#_c_299_n N_A_340_593#_c_561_n 0.0224585f $X=3.8 $Y=1.25 $X2=0
+ $Y2=0
cc_317 N_A_30_131#_c_330_n N_A_340_593#_c_561_n 9.1835e-19 $X=4.92 $Y=3.285
+ $X2=0 $Y2=0
cc_318 N_A_30_131#_c_332_n N_A_340_593#_c_561_n 0.00187353f $X=5.005 $Y=2.24
+ $X2=0 $Y2=0
cc_319 N_A_30_131#_M1006_g N_A_340_593#_c_561_n 0.0435877f $X=3.74 $Y=0.745
+ $X2=0 $Y2=0
cc_320 N_A_30_131#_c_340_n N_A_340_593#_c_561_n 0.0214977f $X=4.645 $Y=3.175
+ $X2=0 $Y2=0
cc_321 N_A_30_131#_c_300_n N_A_340_593#_c_562_n 0.0974818f $X=6.465 $Y=2.24
+ $X2=0 $Y2=0
cc_322 N_A_30_131#_c_332_n N_A_340_593#_c_562_n 0.0137879f $X=5.005 $Y=2.24
+ $X2=0 $Y2=0
cc_323 N_A_30_131#_c_333_n N_A_340_593#_c_562_n 0.00822643f $X=8.63 $Y=2.41
+ $X2=0 $Y2=0
cc_324 N_A_30_131#_c_303_n N_A_340_593#_c_562_n 0.0118943f $X=6.55 $Y=2.24 $X2=0
+ $Y2=0
cc_325 N_A_30_131#_c_340_n N_A_340_593#_c_562_n 0.00226556f $X=4.645 $Y=3.175
+ $X2=0 $Y2=0
cc_326 N_A_30_131#_c_333_n N_A_340_593#_c_581_n 0.0866481f $X=8.63 $Y=2.41 $X2=0
+ $Y2=0
cc_327 N_A_30_131#_c_333_n N_A_340_593#_c_563_n 0.0134853f $X=8.63 $Y=2.41 $X2=0
+ $Y2=0
cc_328 N_A_30_131#_c_338_n N_A_340_593#_c_563_n 0.0043185f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_329 N_A_30_131#_c_304_n N_A_340_593#_c_563_n 0.00640101f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_330 N_A_30_131#_c_310_n N_A_340_593#_c_639_n 0.0351446f $X=8.725 $Y=2.465
+ $X2=0 $Y2=0
cc_331 N_A_30_131#_M1018_g N_A_340_593#_c_564_n 9.05131e-19 $X=9.695 $Y=1.225
+ $X2=0 $Y2=0
cc_332 N_A_30_131#_c_304_n N_A_340_593#_c_564_n 0.0184206f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_333 N_A_30_131#_c_310_n N_A_340_593#_c_642_n 0.00879802f $X=8.725 $Y=2.465
+ $X2=0 $Y2=0
cc_334 N_A_30_131#_c_338_n N_A_340_593#_c_642_n 0.00652509f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_335 N_A_30_131#_c_304_n N_A_340_593#_c_642_n 0.00550126f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_336 N_A_30_131#_c_310_n N_A_340_593#_c_645_n 0.0085211f $X=8.725 $Y=2.465
+ $X2=0 $Y2=0
cc_337 N_A_30_131#_c_338_n N_A_340_593#_c_645_n 0.0132293f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_338 N_A_30_131#_c_310_n N_A_340_593#_c_583_n 0.00613383f $X=8.725 $Y=2.465
+ $X2=0 $Y2=0
cc_339 N_A_30_131#_c_310_n N_A_340_593#_c_586_n 0.00738825f $X=8.725 $Y=2.465
+ $X2=0 $Y2=0
cc_340 N_A_30_131#_c_310_n N_A_340_593#_c_589_n 0.00464054f $X=8.725 $Y=2.465
+ $X2=0 $Y2=0
cc_341 N_A_30_131#_c_338_n N_A_340_593#_c_589_n 0.0280448f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_342 N_A_30_131#_c_304_n N_A_340_593#_c_589_n 0.0332235f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_343 N_A_30_131#_M1028_g N_A_340_593#_c_590_n 0.0321616f $X=1.45 $Y=3.34 $X2=0
+ $Y2=0
cc_344 N_A_30_131#_M1028_g N_A_340_593#_c_591_n 0.0126755f $X=1.45 $Y=3.34 $X2=0
+ $Y2=0
cc_345 N_A_30_131#_c_333_n N_A_340_593#_c_565_n 0.0119737f $X=8.63 $Y=2.41 $X2=0
+ $Y2=0
cc_346 N_A_30_131#_c_333_n N_A_340_593#_c_655_n 0.00591703f $X=8.63 $Y=2.41
+ $X2=0 $Y2=0
cc_347 N_A_30_131#_c_304_n N_A_340_593#_c_655_n 7.26304e-19 $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_348 N_A_30_131#_M1018_g N_A_340_593#_c_566_n 8.96711e-19 $X=9.695 $Y=1.225
+ $X2=0 $Y2=0
cc_349 N_A_30_131#_c_338_n N_A_340_593#_c_566_n 0.0213244f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_350 N_A_30_131#_c_310_n N_A_340_593#_M1030_g 0.0278142f $X=8.725 $Y=2.465
+ $X2=0 $Y2=0
cc_351 N_A_30_131#_c_304_n N_A_340_593#_M1030_g 0.0349466f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_352 N_A_30_131#_c_300_n N_A_1000_81#_c_769_n 0.0156766f $X=6.465 $Y=2.24
+ $X2=0 $Y2=0
cc_353 N_A_30_131#_c_324_n N_A_1000_81#_c_775_n 0.0198784f $X=4.835 $Y=3.45
+ $X2=0 $Y2=0
cc_354 N_A_30_131#_c_330_n N_A_1000_81#_c_775_n 0.0422754f $X=4.92 $Y=3.285
+ $X2=0 $Y2=0
cc_355 N_A_30_131#_c_340_n N_A_1000_81#_c_775_n 8.80594e-19 $X=4.645 $Y=3.175
+ $X2=0 $Y2=0
cc_356 N_A_30_131#_c_300_n N_A_1000_81#_c_777_n 0.0463093f $X=6.465 $Y=2.24
+ $X2=0 $Y2=0
cc_357 N_A_30_131#_c_330_n N_A_1000_81#_c_787_n 0.0129663f $X=4.92 $Y=3.285
+ $X2=0 $Y2=0
cc_358 N_A_30_131#_c_300_n N_A_1000_81#_c_787_n 0.0174582f $X=6.465 $Y=2.24
+ $X2=0 $Y2=0
cc_359 N_A_30_131#_c_300_n N_A_1000_81#_c_789_n 0.00683636f $X=6.465 $Y=2.24
+ $X2=0 $Y2=0
cc_360 N_A_30_131#_c_303_n N_A_1000_81#_c_789_n 0.00680285f $X=6.55 $Y=2.24
+ $X2=0 $Y2=0
cc_361 N_A_30_131#_c_300_n N_A_1000_81#_c_791_n 0.0115442f $X=6.465 $Y=2.24
+ $X2=0 $Y2=0
cc_362 N_A_30_131#_c_333_n N_A_1000_81#_c_778_n 0.0168446f $X=8.63 $Y=2.41 $X2=0
+ $Y2=0
cc_363 N_A_30_131#_c_303_n N_A_1000_81#_c_778_n 0.00352253f $X=6.55 $Y=2.24
+ $X2=0 $Y2=0
cc_364 N_A_30_131#_c_324_n N_A_1000_81#_M1000_g 0.00235202f $X=4.835 $Y=3.45
+ $X2=0 $Y2=0
cc_365 N_A_30_131#_c_330_n N_A_1000_81#_M1000_g 0.0127016f $X=4.92 $Y=3.285
+ $X2=0 $Y2=0
cc_366 N_A_30_131#_c_300_n N_A_1000_81#_M1000_g 0.0119053f $X=6.465 $Y=2.24
+ $X2=0 $Y2=0
cc_367 N_A_30_131#_c_340_n N_A_1000_81#_M1000_g 0.0755629f $X=4.645 $Y=3.175
+ $X2=0 $Y2=0
cc_368 N_A_30_131#_c_333_n N_SET_B_M1026_g 0.0314141f $X=8.63 $Y=2.41 $X2=0
+ $Y2=0
cc_369 N_A_30_131#_c_303_n N_SET_B_M1026_g 0.00355449f $X=6.55 $Y=2.24 $X2=0
+ $Y2=0
cc_370 N_A_30_131#_c_333_n N_SET_B_c_845_n 8.8855e-19 $X=8.63 $Y=2.41 $X2=0
+ $Y2=0
cc_371 N_A_30_131#_M1018_g SET_B 0.0367756f $X=9.695 $Y=1.225 $X2=0 $Y2=0
cc_372 N_A_30_131#_c_300_n N_A_798_107#_c_940_n 0.030712f $X=6.465 $Y=2.24 $X2=0
+ $Y2=0
cc_373 N_A_30_131#_c_333_n N_A_798_107#_c_940_n 3.60328e-19 $X=8.63 $Y=2.41
+ $X2=0 $Y2=0
cc_374 N_A_30_131#_c_303_n N_A_798_107#_c_940_n 0.0168489f $X=6.55 $Y=2.24 $X2=0
+ $Y2=0
cc_375 N_A_30_131#_c_310_n N_A_798_107#_c_951_n 0.0579483f $X=8.725 $Y=2.465
+ $X2=0 $Y2=0
cc_376 N_A_30_131#_c_333_n N_A_798_107#_c_951_n 0.0348328f $X=8.63 $Y=2.41 $X2=0
+ $Y2=0
cc_377 N_A_30_131#_c_338_n N_A_798_107#_c_951_n 0.00102997f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_378 N_A_30_131#_c_304_n N_A_798_107#_c_951_n 0.0579483f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_379 N_A_30_131#_M1006_g N_A_798_107#_c_941_n 0.00381874f $X=3.74 $Y=0.745
+ $X2=0 $Y2=0
cc_380 N_A_30_131#_c_330_n N_A_798_107#_c_954_n 0.00951973f $X=4.92 $Y=3.285
+ $X2=0 $Y2=0
cc_381 N_A_30_131#_c_340_n N_A_798_107#_c_954_n 0.0013713f $X=4.645 $Y=3.175
+ $X2=0 $Y2=0
cc_382 N_A_30_131#_c_324_n N_A_798_107#_c_955_n 0.02534f $X=4.835 $Y=3.45 $X2=0
+ $Y2=0
cc_383 N_A_30_131#_c_327_n N_A_798_107#_c_955_n 3.98316e-19 $X=4.565 $Y=3.45
+ $X2=0 $Y2=0
cc_384 N_A_30_131#_c_299_n N_A_798_107#_c_946_n 0.00386412f $X=3.8 $Y=1.25 $X2=0
+ $Y2=0
cc_385 N_A_30_131#_M1006_g N_A_798_107#_c_946_n 0.00234597f $X=3.74 $Y=0.745
+ $X2=0 $Y2=0
cc_386 N_A_30_131#_c_299_n N_A_798_107#_c_947_n 0.13349f $X=3.8 $Y=1.25 $X2=0
+ $Y2=0
cc_387 N_A_30_131#_c_330_n N_A_798_107#_c_947_n 0.00838803f $X=4.92 $Y=3.285
+ $X2=0 $Y2=0
cc_388 N_A_30_131#_c_332_n N_A_798_107#_c_947_n 0.00532449f $X=5.005 $Y=2.24
+ $X2=0 $Y2=0
cc_389 N_A_30_131#_M1006_g N_A_798_107#_c_947_n 0.00494535f $X=3.74 $Y=0.745
+ $X2=0 $Y2=0
cc_390 N_A_30_131#_c_340_n N_A_798_107#_c_947_n 9.86757e-19 $X=4.645 $Y=3.175
+ $X2=0 $Y2=0
cc_391 N_A_30_131#_M1018_g N_A_2031_177#_c_1067_n 0.00207779f $X=9.695 $Y=1.225
+ $X2=0 $Y2=0
cc_392 N_A_30_131#_M1018_g N_A_2031_177#_M1019_g 0.0989115f $X=9.695 $Y=1.225
+ $X2=0 $Y2=0
cc_393 N_A_30_131#_M1018_g N_A_1787_137#_c_1131_n 0.0211334f $X=9.695 $Y=1.225
+ $X2=0 $Y2=0
cc_394 N_A_30_131#_c_304_n N_A_1787_137#_c_1131_n 0.00654989f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_395 N_A_30_131#_c_310_n N_A_1787_137#_c_1143_n 0.00471572f $X=8.725 $Y=2.465
+ $X2=0 $Y2=0
cc_396 N_A_30_131#_c_304_n N_A_1787_137#_c_1143_n 4.66604e-19 $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_397 N_A_30_131#_M1018_g N_A_1787_137#_c_1144_n 0.0176441f $X=9.695 $Y=1.225
+ $X2=0 $Y2=0
cc_398 N_A_30_131#_c_304_n N_A_1787_137#_c_1144_n 0.0247524f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_399 N_A_30_131#_c_310_n N_A_1787_137#_c_1155_n 9.7708e-19 $X=8.725 $Y=2.465
+ $X2=0 $Y2=0
cc_400 N_A_30_131#_c_304_n N_A_1787_137#_c_1145_n 0.00668953f $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_401 N_A_30_131#_c_304_n N_A_1787_137#_c_1146_n 8.57804e-19 $X=8.795 $Y=2.25
+ $X2=0 $Y2=0
cc_402 N_A_30_131#_M1028_g N_VPWR_c_1317_n 0.0522661f $X=1.45 $Y=3.34 $X2=0
+ $Y2=0
cc_403 N_A_30_131#_c_288_n N_VPWR_c_1317_n 0.0364612f $X=0.28 $Y=3.11 $X2=0
+ $Y2=0
cc_404 N_A_30_131#_M1028_g N_VPWR_c_1320_n 0.0024653f $X=1.45 $Y=3.34 $X2=0
+ $Y2=0
cc_405 N_A_30_131#_c_324_n N_VPWR_c_1323_n 8.63964e-19 $X=4.835 $Y=3.45 $X2=0
+ $Y2=0
cc_406 N_A_30_131#_c_327_n N_VPWR_c_1323_n 4.617e-19 $X=4.565 $Y=3.45 $X2=0
+ $Y2=0
cc_407 N_A_30_131#_c_310_n N_VPWR_c_1326_n 0.00303846f $X=8.725 $Y=2.465 $X2=0
+ $Y2=0
cc_408 N_A_30_131#_c_333_n N_VPWR_c_1326_n 0.0666112f $X=8.63 $Y=2.41 $X2=0
+ $Y2=0
cc_409 N_A_30_131#_M1016_s N_VPWR_c_1338_n 0.00221032f $X=0.155 $Y=2.965 $X2=0
+ $Y2=0
cc_410 N_A_30_131#_M1028_g N_VPWR_c_1338_n 0.0110801f $X=1.45 $Y=3.34 $X2=0
+ $Y2=0
cc_411 N_A_30_131#_c_310_n N_VPWR_c_1338_n 0.0180453f $X=8.725 $Y=2.465 $X2=0
+ $Y2=0
cc_412 N_A_30_131#_c_288_n N_VPWR_c_1338_n 0.034265f $X=0.28 $Y=3.11 $X2=0 $Y2=0
cc_413 N_A_30_131#_c_317_n N_VPWR_c_1338_n 0.0337605f $X=3.715 $Y=3.45 $X2=0
+ $Y2=0
cc_414 N_A_30_131#_c_320_n N_VPWR_c_1338_n 0.0119633f $X=3.185 $Y=3.45 $X2=0
+ $Y2=0
cc_415 N_A_30_131#_c_324_n N_VPWR_c_1338_n 0.0832049f $X=4.835 $Y=3.45 $X2=0
+ $Y2=0
cc_416 N_A_30_131#_c_327_n N_VPWR_c_1338_n 0.00622526f $X=4.565 $Y=3.45 $X2=0
+ $Y2=0
cc_417 N_A_30_131#_c_335_n N_VPWR_c_1338_n 0.0152705f $X=3.8 $Y=3.45 $X2=0 $Y2=0
cc_418 N_A_30_131#_c_296_n N_A_642_107#_c_1438_n 0.0129669f $X=3.015 $Y=1.26
+ $X2=0 $Y2=0
cc_419 N_A_30_131#_c_298_n N_A_642_107#_c_1438_n 0.106103f $X=3.1 $Y=3.285 $X2=0
+ $Y2=0
cc_420 N_A_30_131#_c_317_n N_A_642_107#_c_1438_n 0.0132499f $X=3.715 $Y=3.45
+ $X2=0 $Y2=0
cc_421 N_A_30_131#_c_299_n N_A_642_107#_c_1438_n 0.121499f $X=3.8 $Y=1.25 $X2=0
+ $Y2=0
cc_422 N_A_30_131#_M1006_g N_A_642_107#_c_1438_n 0.0212432f $X=3.74 $Y=0.745
+ $X2=0 $Y2=0
cc_423 N_A_30_131#_M1006_g N_A_642_107#_c_1439_n 0.0143774f $X=3.74 $Y=0.745
+ $X2=0 $Y2=0
cc_424 N_A_30_131#_c_330_n A_982_529# 0.00353241f $X=4.92 $Y=3.285 $X2=0 $Y2=0
cc_425 N_A_30_131#_M1029_g N_VGND_c_1476_n 0.00152888f $X=1.465 $Y=0.865 $X2=0
+ $Y2=0
cc_426 N_A_30_131#_c_286_n N_VGND_c_1476_n 0.0215213f $X=0.295 $Y=0.865 $X2=0
+ $Y2=0
cc_427 N_A_30_131#_c_289_n N_VGND_c_1476_n 0.0446459f $X=1.18 $Y=1.38 $X2=0
+ $Y2=0
cc_428 N_A_30_131#_c_290_n N_VGND_c_1476_n 0.0314214f $X=1.425 $Y=1.295 $X2=0
+ $Y2=0
cc_429 N_A_30_131#_c_293_n N_VGND_c_1476_n 0.00488837f $X=1.51 $Y=0.35 $X2=0
+ $Y2=0
cc_430 N_A_30_131#_c_291_n N_VGND_c_1478_n 0.00488091f $X=2.12 $Y=0.35 $X2=0
+ $Y2=0
cc_431 N_A_30_131#_c_295_n N_VGND_c_1478_n 0.0414645f $X=2.205 $Y=1.175 $X2=0
+ $Y2=0
cc_432 N_A_30_131#_c_296_n N_VGND_c_1478_n 0.0392731f $X=3.015 $Y=1.26 $X2=0
+ $Y2=0
cc_433 N_A_30_131#_M1006_g N_VGND_c_1478_n 8.39755e-19 $X=3.74 $Y=0.745 $X2=0
+ $Y2=0
cc_434 N_A_30_131#_M1029_g N_VGND_c_1488_n 0.0199945f $X=1.465 $Y=0.865 $X2=0
+ $Y2=0
cc_435 N_A_30_131#_c_286_n N_VGND_c_1488_n 0.0210742f $X=0.295 $Y=0.865 $X2=0
+ $Y2=0
cc_436 N_A_30_131#_c_290_n N_VGND_c_1488_n 0.0195194f $X=1.425 $Y=1.295 $X2=0
+ $Y2=0
cc_437 N_A_30_131#_c_291_n N_VGND_c_1488_n 0.0329517f $X=2.12 $Y=0.35 $X2=0
+ $Y2=0
cc_438 N_A_30_131#_c_293_n N_VGND_c_1488_n 0.00777234f $X=1.51 $Y=0.35 $X2=0
+ $Y2=0
cc_439 N_A_30_131#_c_295_n N_VGND_c_1488_n 0.0198019f $X=2.205 $Y=1.175 $X2=0
+ $Y2=0
cc_440 N_A_30_131#_c_296_n N_VGND_c_1488_n 0.0138792f $X=3.015 $Y=1.26 $X2=0
+ $Y2=0
cc_441 N_A_30_131#_c_299_n N_VGND_c_1488_n 0.00597472f $X=3.8 $Y=1.25 $X2=0
+ $Y2=0
cc_442 N_A_30_131#_c_302_n N_VGND_c_1488_n 0.00136403f $X=1.345 $Y=1.425 $X2=0
+ $Y2=0
cc_443 N_A_30_131#_M1006_g N_VGND_c_1488_n 0.0253541f $X=3.74 $Y=0.745 $X2=0
+ $Y2=0
cc_444 N_D_M1002_g N_A_340_593#_M1024_g 0.0169185f $X=3.06 $Y=2.855 $X2=0.24
+ $Y2=0
cc_445 N_D_M1002_g N_A_340_593#_c_568_n 0.0353351f $X=3.06 $Y=2.855 $X2=0 $Y2=0
cc_446 N_D_c_525_n N_A_340_593#_c_560_n 0.0219567f $X=3.06 $Y=2.515 $X2=0 $Y2=0
cc_447 D N_A_340_593#_c_560_n 0.0178403f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_448 N_D_c_525_n N_A_340_593#_c_575_n 0.0246749f $X=3.06 $Y=2.515 $X2=0 $Y2=0
cc_449 D N_A_340_593#_c_575_n 0.0248407f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_450 N_D_c_525_n N_A_340_593#_c_576_n 0.00714658f $X=3.06 $Y=2.515 $X2=0 $Y2=0
cc_451 N_D_M1002_g N_A_340_593#_c_576_n 0.0230283f $X=3.06 $Y=2.855 $X2=0 $Y2=0
cc_452 N_D_c_525_n N_A_340_593#_c_561_n 0.0169185f $X=3.06 $Y=2.515 $X2=0 $Y2=0
cc_453 N_D_c_525_n N_A_340_593#_c_590_n 0.0015494f $X=3.06 $Y=2.515 $X2=0 $Y2=0
cc_454 N_D_M1002_g N_VPWR_c_1320_n 0.00287869f $X=3.06 $Y=2.855 $X2=0 $Y2=0
cc_455 N_D_M1002_g N_VPWR_c_1338_n 0.00108457f $X=3.06 $Y=2.855 $X2=0 $Y2=0
cc_456 N_D_M1027_g N_A_642_107#_c_1438_n 0.00883576f $X=2.96 $Y=0.745 $X2=0
+ $Y2=0
cc_457 N_D_c_525_n N_A_642_107#_c_1438_n 0.00649497f $X=3.06 $Y=2.515 $X2=0
+ $Y2=0
cc_458 N_D_M1027_g N_A_642_107#_c_1439_n 0.0102143f $X=2.96 $Y=0.745 $X2=0 $Y2=0
cc_459 N_D_M1027_g N_VGND_c_1478_n 0.0369275f $X=2.96 $Y=0.745 $X2=0 $Y2=0
cc_460 N_D_c_525_n N_VGND_c_1478_n 0.00129608f $X=3.06 $Y=2.515 $X2=0 $Y2=0
cc_461 N_D_M1027_g N_VGND_c_1488_n 0.00553004f $X=2.96 $Y=0.745 $X2=0 $Y2=0
cc_462 N_A_340_593#_M1023_g N_A_1000_81#_M1003_g 0.0444555f $X=4.54 $Y=0.745
+ $X2=0 $Y2=0
cc_463 N_A_340_593#_c_562_n N_A_1000_81#_c_769_n 0.00361709f $X=6.815 $Y=1.89
+ $X2=0 $Y2=0
cc_464 N_A_340_593#_c_623_n N_A_1000_81#_c_770_n 0.00105158f $X=4.535 $Y=1.805
+ $X2=0 $Y2=0
cc_465 N_A_340_593#_c_674_p N_A_1000_81#_c_770_n 7.80729e-19 $X=4.535 $Y=1.66
+ $X2=0 $Y2=0
cc_466 N_A_340_593#_c_561_n N_A_1000_81#_c_770_n 0.0224949f $X=4.535 $Y=1.66
+ $X2=0 $Y2=0
cc_467 N_A_340_593#_c_562_n N_A_1000_81#_c_770_n 0.0215411f $X=6.815 $Y=1.89
+ $X2=0 $Y2=0
cc_468 N_A_340_593#_c_674_p N_A_1000_81#_c_771_n 5.94638e-19 $X=4.535 $Y=1.66
+ $X2=14.64 $Y2=0
cc_469 N_A_340_593#_c_561_n N_A_1000_81#_c_771_n 0.0444555f $X=4.535 $Y=1.66
+ $X2=14.64 $Y2=0
cc_470 N_A_340_593#_c_562_n N_A_1000_81#_c_771_n 0.00384947f $X=6.815 $Y=1.89
+ $X2=14.64 $Y2=0
cc_471 N_A_340_593#_M1023_g N_A_1000_81#_c_772_n 0.00140515f $X=4.54 $Y=0.745
+ $X2=0 $Y2=0
cc_472 N_A_340_593#_c_674_p N_A_1000_81#_c_772_n 0.00431324f $X=4.535 $Y=1.66
+ $X2=0 $Y2=0
cc_473 N_A_340_593#_c_562_n N_A_1000_81#_c_772_n 0.0496217f $X=6.815 $Y=1.89
+ $X2=0 $Y2=0
cc_474 N_A_340_593#_c_581_n N_SET_B_M1026_g 0.010681f $X=8.28 $Y=2.06 $X2=0
+ $Y2=0
cc_475 N_A_340_593#_c_565_n N_SET_B_M1026_g 0.00348933f $X=6.9 $Y=1.89 $X2=0
+ $Y2=0
cc_476 N_A_340_593#_c_581_n N_SET_B_c_844_n 0.06484f $X=8.28 $Y=2.06 $X2=14.64
+ $Y2=0
cc_477 N_A_340_593#_c_563_n N_SET_B_c_844_n 0.0183608f $X=8.45 $Y=1.71 $X2=14.64
+ $Y2=0
cc_478 N_A_340_593#_c_562_n N_SET_B_c_845_n 3.8428e-19 $X=6.815 $Y=1.89 $X2=0
+ $Y2=0
cc_479 N_A_340_593#_c_581_n N_SET_B_c_845_n 0.0164783f $X=8.28 $Y=2.06 $X2=0
+ $Y2=0
cc_480 N_A_340_593#_c_565_n N_SET_B_c_845_n 0.0147455f $X=6.9 $Y=1.89 $X2=0
+ $Y2=0
cc_481 N_A_340_593#_c_558_n N_SET_B_c_868_n 0.00303124f $X=8.685 $Y=1.315
+ $X2=7.44 $Y2=0.057
cc_482 N_A_340_593#_c_563_n N_SET_B_c_868_n 6.52697e-19 $X=8.45 $Y=1.71 $X2=7.44
+ $Y2=0.057
cc_483 N_A_340_593#_c_558_n SET_B 0.0455135f $X=8.685 $Y=1.315 $X2=0 $Y2=0
cc_484 N_A_340_593#_c_566_n SET_B 0.00502241f $X=8.785 $Y=1.71 $X2=0 $Y2=0
cc_485 N_A_340_593#_c_558_n N_SET_B_c_850_n 0.00897016f $X=8.685 $Y=1.315 $X2=0
+ $Y2=0
cc_486 N_A_340_593#_c_563_n N_SET_B_c_850_n 0.00529082f $X=8.45 $Y=1.71 $X2=0
+ $Y2=0
cc_487 N_A_340_593#_c_655_n N_SET_B_c_850_n 0.00502241f $X=8.62 $Y=1.71 $X2=0
+ $Y2=0
cc_488 N_A_340_593#_c_558_n N_A_798_107#_c_938_n 0.0898934f $X=8.685 $Y=1.315
+ $X2=0 $Y2=0
cc_489 N_A_340_593#_c_581_n N_A_798_107#_M1013_g 0.0187186f $X=8.28 $Y=2.06
+ $X2=0 $Y2=0
cc_490 N_A_340_593#_c_563_n N_A_798_107#_M1013_g 0.00918332f $X=8.45 $Y=1.71
+ $X2=0 $Y2=0
cc_491 N_A_340_593#_c_562_n N_A_798_107#_c_940_n 0.04982f $X=6.815 $Y=1.89 $X2=0
+ $Y2=0
cc_492 N_A_340_593#_c_565_n N_A_798_107#_c_940_n 0.003631f $X=6.9 $Y=1.89 $X2=0
+ $Y2=0
cc_493 N_A_340_593#_c_581_n N_A_798_107#_c_951_n 0.012213f $X=8.28 $Y=2.06 $X2=0
+ $Y2=0
cc_494 N_A_340_593#_c_639_n N_A_798_107#_c_951_n 0.00226459f $X=8.78 $Y=3.595
+ $X2=0 $Y2=0
cc_495 N_A_340_593#_c_645_n N_A_798_107#_c_951_n 5.0429e-19 $X=8.865 $Y=2.76
+ $X2=0 $Y2=0
cc_496 N_A_340_593#_c_583_n N_A_798_107#_c_951_n 3.77774e-19 $X=8.865 $Y=3.7
+ $X2=0 $Y2=0
cc_497 N_A_340_593#_M1023_g N_A_798_107#_c_941_n 0.0116057f $X=4.54 $Y=0.745
+ $X2=0 $Y2=0
cc_498 N_A_340_593#_M1024_g N_A_798_107#_c_954_n 0.00338232f $X=3.84 $Y=2.855
+ $X2=0 $Y2=0
cc_499 N_A_340_593#_c_561_n N_A_798_107#_c_954_n 0.00597303f $X=4.535 $Y=1.66
+ $X2=0 $Y2=0
cc_500 N_A_340_593#_M1024_g N_A_798_107#_c_955_n 0.00655295f $X=3.84 $Y=2.855
+ $X2=0 $Y2=0
cc_501 N_A_340_593#_M1023_g N_A_798_107#_c_943_n 0.0307297f $X=4.54 $Y=0.745
+ $X2=0 $Y2=0
cc_502 N_A_340_593#_c_674_p N_A_798_107#_c_943_n 0.00989034f $X=4.535 $Y=1.66
+ $X2=0 $Y2=0
cc_503 N_A_340_593#_c_562_n N_A_798_107#_c_943_n 0.0227902f $X=6.815 $Y=1.89
+ $X2=0 $Y2=0
cc_504 N_A_340_593#_M1023_g N_A_798_107#_c_946_n 0.00325849f $X=4.54 $Y=0.745
+ $X2=0 $Y2=0
cc_505 N_A_340_593#_c_561_n N_A_798_107#_c_946_n 0.00219114f $X=4.535 $Y=1.66
+ $X2=0 $Y2=0
cc_506 N_A_340_593#_M1024_g N_A_798_107#_c_947_n 0.00166784f $X=3.84 $Y=2.855
+ $X2=0 $Y2=0
cc_507 N_A_340_593#_M1023_g N_A_798_107#_c_947_n 0.00865842f $X=4.54 $Y=0.745
+ $X2=0 $Y2=0
cc_508 N_A_340_593#_c_623_n N_A_798_107#_c_947_n 0.0250672f $X=4.535 $Y=1.805
+ $X2=0 $Y2=0
cc_509 N_A_340_593#_c_674_p N_A_798_107#_c_947_n 0.0205827f $X=4.535 $Y=1.66
+ $X2=0 $Y2=0
cc_510 N_A_340_593#_c_561_n N_A_798_107#_c_947_n 0.0454985f $X=4.535 $Y=1.66
+ $X2=0 $Y2=0
cc_511 N_A_340_593#_M1030_g N_A_2031_177#_M1019_g 0.0455396f $X=9.695 $Y=2.785
+ $X2=0 $Y2=0
cc_512 N_A_340_593#_c_642_n N_A_1787_137#_M1014_d 0.00738526f $X=9.14 $Y=2.76
+ $X2=0 $Y2=0
cc_513 N_A_340_593#_c_589_n N_A_1787_137#_M1014_d 0.002229f $X=9.225 $Y=2.675
+ $X2=0 $Y2=0
cc_514 N_A_340_593#_c_558_n N_A_1787_137#_c_1131_n 0.00967637f $X=8.685 $Y=1.315
+ $X2=0 $Y2=0
cc_515 N_A_340_593#_c_564_n N_A_1787_137#_c_1131_n 0.0192994f $X=9.14 $Y=1.79
+ $X2=0 $Y2=0
cc_516 N_A_340_593#_c_639_n N_A_1787_137#_c_1143_n 0.0290535f $X=8.78 $Y=3.595
+ $X2=0 $Y2=0
cc_517 N_A_340_593#_c_642_n N_A_1787_137#_c_1143_n 0.0203672f $X=9.14 $Y=2.76
+ $X2=0 $Y2=0
cc_518 N_A_340_593#_c_586_n N_A_1787_137#_c_1143_n 0.0384071f $X=9.66 $Y=3.68
+ $X2=0 $Y2=0
cc_519 N_A_340_593#_M1030_g N_A_1787_137#_c_1143_n 0.0251331f $X=9.695 $Y=2.785
+ $X2=0 $Y2=0
cc_520 N_A_340_593#_c_558_n N_A_1787_137#_c_1144_n 5.26491e-19 $X=8.685 $Y=1.315
+ $X2=0 $Y2=0
cc_521 N_A_340_593#_c_564_n N_A_1787_137#_c_1144_n 0.012652f $X=9.14 $Y=1.79
+ $X2=0 $Y2=0
cc_522 N_A_340_593#_c_589_n N_A_1787_137#_c_1144_n 0.0290247f $X=9.225 $Y=2.675
+ $X2=0 $Y2=0
cc_523 N_A_340_593#_c_639_n N_A_1787_137#_c_1155_n 0.00411546f $X=8.78 $Y=3.595
+ $X2=0 $Y2=0
cc_524 N_A_340_593#_c_642_n N_A_1787_137#_c_1155_n 0.0127298f $X=9.14 $Y=2.76
+ $X2=0 $Y2=0
cc_525 N_A_340_593#_c_589_n N_A_1787_137#_c_1155_n 0.0128166f $X=9.225 $Y=2.675
+ $X2=0 $Y2=0
cc_526 N_A_340_593#_M1030_g N_A_1787_137#_c_1155_n 0.0220158f $X=9.695 $Y=2.785
+ $X2=0 $Y2=0
cc_527 N_A_340_593#_M1030_g N_A_1787_137#_c_1145_n 0.015417f $X=9.695 $Y=2.785
+ $X2=0 $Y2=0
cc_528 N_A_340_593#_c_589_n N_A_1787_137#_c_1146_n 0.0136026f $X=9.225 $Y=2.675
+ $X2=0 $Y2=0
cc_529 N_A_340_593#_M1030_g N_A_1787_137#_c_1146_n 0.00243934f $X=9.695 $Y=2.785
+ $X2=0 $Y2=0
cc_530 N_A_340_593#_c_576_n N_VPWR_M1002_s 0.00458388f $X=2.75 $Y=3.59 $X2=0
+ $Y2=0
cc_531 N_A_340_593#_c_571_n N_VPWR_c_1317_n 0.055719f $X=1.84 $Y=3.11 $X2=0
+ $Y2=0
cc_532 N_A_340_593#_c_590_n N_VPWR_c_1317_n 0.00138547f $X=1.84 $Y=2.945 $X2=0
+ $Y2=0
cc_533 N_A_340_593#_c_568_n N_VPWR_c_1320_n 0.00679253f $X=3.59 $Y=3.655 $X2=0
+ $Y2=0
cc_534 N_A_340_593#_c_575_n N_VPWR_c_1320_n 0.0201141f $X=2.665 $Y=2.36 $X2=0
+ $Y2=0
cc_535 N_A_340_593#_c_576_n N_VPWR_c_1320_n 0.0764407f $X=2.75 $Y=3.59 $X2=0
+ $Y2=0
cc_536 N_A_340_593#_c_590_n N_VPWR_c_1320_n 0.0678671f $X=1.84 $Y=2.945 $X2=0
+ $Y2=0
cc_537 N_A_340_593#_c_639_n N_VPWR_c_1326_n 0.0156774f $X=8.78 $Y=3.595 $X2=0
+ $Y2=0
cc_538 N_A_340_593#_c_645_n N_VPWR_c_1326_n 0.00449661f $X=8.865 $Y=2.76 $X2=0
+ $Y2=0
cc_539 N_A_340_593#_c_583_n N_VPWR_c_1326_n 9.2789e-19 $X=8.865 $Y=3.7 $X2=0
+ $Y2=0
cc_540 N_A_340_593#_c_586_n N_VPWR_c_1329_n 0.00698841f $X=9.66 $Y=3.68 $X2=0
+ $Y2=0
cc_541 N_A_340_593#_M1030_g N_VPWR_c_1329_n 0.0242748f $X=9.695 $Y=2.785 $X2=0
+ $Y2=0
cc_542 N_A_340_593#_c_568_n N_VPWR_c_1338_n 0.0251964f $X=3.59 $Y=3.655 $X2=0
+ $Y2=0
cc_543 N_A_340_593#_c_571_n N_VPWR_c_1338_n 0.038667f $X=1.84 $Y=3.11 $X2=0
+ $Y2=0
cc_544 N_A_340_593#_c_576_n N_VPWR_c_1338_n 0.024823f $X=2.75 $Y=3.59 $X2=0
+ $Y2=0
cc_545 N_A_340_593#_c_639_n N_VPWR_c_1338_n 0.0199241f $X=8.78 $Y=3.595 $X2=0
+ $Y2=0
cc_546 N_A_340_593#_c_642_n N_VPWR_c_1338_n 0.00536293f $X=9.14 $Y=2.76 $X2=0
+ $Y2=0
cc_547 N_A_340_593#_c_583_n N_VPWR_c_1338_n 0.0103651f $X=8.865 $Y=3.7 $X2=0
+ $Y2=0
cc_548 N_A_340_593#_c_586_n N_VPWR_c_1338_n 0.0385663f $X=9.66 $Y=3.68 $X2=0
+ $Y2=0
cc_549 N_A_340_593#_M1030_g N_VPWR_c_1338_n 0.0247621f $X=9.695 $Y=2.785 $X2=0
+ $Y2=0
cc_550 N_A_340_593#_c_568_n N_A_642_107#_c_1438_n 9.85483e-19 $X=3.59 $Y=3.655
+ $X2=0 $Y2=0
cc_551 N_A_340_593#_c_561_n N_A_642_107#_c_1438_n 0.00583109f $X=4.535 $Y=1.66
+ $X2=0 $Y2=0
cc_552 N_A_340_593#_M1023_g N_VGND_c_1480_n 0.00573023f $X=4.54 $Y=0.745 $X2=0
+ $Y2=0
cc_553 N_A_340_593#_c_558_n N_VGND_c_1482_n 3.17681e-19 $X=8.685 $Y=1.315 $X2=0
+ $Y2=0
cc_554 N_A_340_593#_c_581_n N_VGND_c_1482_n 0.00481635f $X=8.28 $Y=2.06 $X2=0
+ $Y2=0
cc_555 N_A_340_593#_c_565_n N_VGND_c_1482_n 0.00581331f $X=6.9 $Y=1.89 $X2=0
+ $Y2=0
cc_556 N_A_340_593#_M1023_g N_VGND_c_1488_n 0.0160574f $X=4.54 $Y=0.745 $X2=0
+ $Y2=0
cc_557 N_A_340_593#_c_558_n N_VGND_c_1488_n 0.00622132f $X=8.685 $Y=1.315 $X2=0
+ $Y2=0
cc_558 N_A_340_593#_c_560_n N_VGND_c_1488_n 0.0173761f $X=1.855 $Y=0.865 $X2=0
+ $Y2=0
cc_559 N_A_1000_81#_c_791_n N_SET_B_M1026_g 6.64176e-19 $X=6.2 $Y=2.59 $X2=0
+ $Y2=0
cc_560 N_A_1000_81#_c_778_n N_SET_B_M1026_g 0.00859337f $X=6.73 $Y=2.76 $X2=0
+ $Y2=0
cc_561 N_A_1000_81#_M1003_g N_A_798_107#_c_935_n 0.0175391f $X=5.25 $Y=0.745
+ $X2=0 $Y2=0
cc_562 N_A_1000_81#_c_771_n N_A_798_107#_M1025_g 0.0175391f $X=5.3 $Y=1.47
+ $X2=0.24 $Y2=0
cc_563 N_A_1000_81#_c_772_n N_A_798_107#_M1025_g 0.0163619f $X=5.7 $Y=1.465
+ $X2=0.24 $Y2=0
cc_564 N_A_1000_81#_c_775_n N_A_798_107#_M1009_g 8.98982e-19 $X=5.305 $Y=3.39
+ $X2=0 $Y2=0
cc_565 N_A_1000_81#_c_777_n N_A_798_107#_M1009_g 0.00512649f $X=6.115 $Y=2.59
+ $X2=0 $Y2=0
cc_566 N_A_1000_81#_c_789_n N_A_798_107#_M1009_g 0.0171568f $X=6.565 $Y=2.76
+ $X2=0 $Y2=0
cc_567 N_A_1000_81#_c_791_n N_A_798_107#_M1009_g 0.0158029f $X=6.2 $Y=2.59 $X2=0
+ $Y2=0
cc_568 N_A_1000_81#_c_778_n N_A_798_107#_M1009_g 0.0100447f $X=6.73 $Y=2.76
+ $X2=0 $Y2=0
cc_569 N_A_1000_81#_M1000_g N_A_798_107#_M1009_g 0.0115579f $X=5.37 $Y=2.855
+ $X2=0 $Y2=0
cc_570 N_A_1000_81#_c_769_n N_A_798_107#_c_940_n 0.0345076f $X=5.37 $Y=2.285
+ $X2=0 $Y2=0
cc_571 N_A_1000_81#_c_770_n N_A_798_107#_c_940_n 0.0175391f $X=5.37 $Y=2.035
+ $X2=0 $Y2=0
cc_572 N_A_1000_81#_c_777_n N_A_798_107#_c_940_n 0.00864026f $X=6.115 $Y=2.59
+ $X2=0 $Y2=0
cc_573 N_A_1000_81#_c_791_n N_A_798_107#_c_940_n 0.00280332f $X=6.2 $Y=2.59
+ $X2=0 $Y2=0
cc_574 N_A_1000_81#_M1003_g N_A_798_107#_c_941_n 7.89449e-19 $X=5.25 $Y=0.745
+ $X2=0 $Y2=0
cc_575 N_A_1000_81#_M1003_g N_A_798_107#_c_943_n 0.0274141f $X=5.25 $Y=0.745
+ $X2=0 $Y2=0
cc_576 N_A_1000_81#_c_772_n N_A_798_107#_c_943_n 0.0496218f $X=5.7 $Y=1.465
+ $X2=0 $Y2=0
cc_577 N_A_1000_81#_M1003_g N_A_798_107#_c_944_n 8.74964e-19 $X=5.25 $Y=0.745
+ $X2=0 $Y2=0
cc_578 N_A_1000_81#_c_777_n N_VPWR_M1000_d 0.00657569f $X=6.115 $Y=2.59 $X2=0
+ $Y2=0
cc_579 N_A_1000_81#_c_775_n N_VPWR_c_1323_n 0.0480121f $X=5.305 $Y=3.39 $X2=0
+ $Y2=0
cc_580 N_A_1000_81#_c_777_n N_VPWR_c_1323_n 0.0210122f $X=6.115 $Y=2.59 $X2=0
+ $Y2=0
cc_581 N_A_1000_81#_c_778_n N_VPWR_c_1323_n 0.00694629f $X=6.73 $Y=2.76 $X2=0
+ $Y2=0
cc_582 N_A_1000_81#_M1000_g N_VPWR_c_1323_n 0.0247787f $X=5.37 $Y=2.855 $X2=0
+ $Y2=0
cc_583 N_A_1000_81#_c_778_n N_VPWR_c_1326_n 0.0326319f $X=6.73 $Y=2.76 $X2=0
+ $Y2=0
cc_584 N_A_1000_81#_c_775_n N_VPWR_c_1338_n 0.0224424f $X=5.305 $Y=3.39 $X2=0
+ $Y2=0
cc_585 N_A_1000_81#_c_789_n N_VPWR_c_1338_n 0.00840658f $X=6.565 $Y=2.76 $X2=0
+ $Y2=0
cc_586 N_A_1000_81#_c_791_n N_VPWR_c_1338_n 0.00538432f $X=6.2 $Y=2.59 $X2=0
+ $Y2=0
cc_587 N_A_1000_81#_c_778_n N_VPWR_c_1338_n 0.0150071f $X=6.73 $Y=2.76 $X2=0
+ $Y2=0
cc_588 N_A_1000_81#_M1000_g N_VPWR_c_1338_n 0.0177082f $X=5.37 $Y=2.855 $X2=0
+ $Y2=0
cc_589 N_A_1000_81#_M1003_g N_VGND_c_1480_n 0.0361332f $X=5.25 $Y=0.745 $X2=0
+ $Y2=0
cc_590 N_SET_B_c_849_n N_A_798_107#_M1025_g 0.0212192f $X=7.182 $Y=1.545
+ $X2=0.24 $Y2=0
cc_591 N_SET_B_c_849_n N_A_798_107#_c_938_n 0.0200157f $X=7.182 $Y=1.545 $X2=0
+ $Y2=0
cc_592 N_SET_B_c_850_n N_A_798_107#_c_938_n 0.00385884f $X=8.512 $Y=0.782 $X2=0
+ $Y2=0
cc_593 N_SET_B_M1026_g N_A_798_107#_M1013_g 0.0168954f $X=7.12 $Y=2.855 $X2=0
+ $Y2=0
cc_594 N_SET_B_c_844_n N_A_798_107#_M1013_g 0.0265885f $X=7.93 $Y=1.675 $X2=0
+ $Y2=0
cc_595 N_SET_B_c_845_n N_A_798_107#_M1013_g 0.0355939f $X=7.33 $Y=1.71 $X2=0
+ $Y2=0
cc_596 N_SET_B_c_868_n N_A_798_107#_M1013_g 0.0242312f $X=8.015 $Y=1.555 $X2=0
+ $Y2=0
cc_597 N_SET_B_c_884_p N_A_798_107#_M1013_g 0.00844857f $X=8.1 $Y=0.925 $X2=0
+ $Y2=0
cc_598 N_SET_B_c_849_n N_A_798_107#_M1013_g 0.0142232f $X=7.182 $Y=1.545 $X2=0
+ $Y2=0
cc_599 N_SET_B_c_886_p N_A_798_107#_M1013_g 0.0110049f $X=8.285 $Y=0.782 $X2=0
+ $Y2=0
cc_600 N_SET_B_M1026_g N_A_798_107#_c_940_n 0.0375841f $X=7.12 $Y=2.855 $X2=0
+ $Y2=0
cc_601 N_SET_B_c_845_n N_A_798_107#_c_940_n 0.0134475f $X=7.33 $Y=1.71 $X2=0
+ $Y2=0
cc_602 N_SET_B_M1026_g N_A_798_107#_c_951_n 0.0140794f $X=7.12 $Y=2.855 $X2=0
+ $Y2=0
cc_603 N_SET_B_c_842_n N_A_2031_177#_c_1055_n 0.0431068f $X=11.15 $Y=1.85 $X2=0
+ $Y2=0
cc_604 SET_B N_A_2031_177#_c_1055_n 0.0076953f $X=10.715 $Y=0.84 $X2=0 $Y2=0
cc_605 N_SET_B_c_892_p N_A_2031_177#_c_1055_n 0.00697984f $X=11.05 $Y=0.72 $X2=0
+ $Y2=0
cc_606 N_SET_B_M1010_g N_A_2031_177#_c_1060_n 0.0114543f $X=11.185 $Y=2.785
+ $X2=0 $Y2=0
cc_607 N_SET_B_c_842_n N_A_2031_177#_c_1056_n 2.76638e-19 $X=11.15 $Y=1.85
+ $X2=14.64 $Y2=0
cc_608 N_SET_B_c_842_n N_A_2031_177#_c_1067_n 0.00231906f $X=11.15 $Y=1.85 $X2=0
+ $Y2=0
cc_609 SET_B N_A_2031_177#_c_1067_n 0.0103312f $X=10.715 $Y=0.84 $X2=0 $Y2=0
cc_610 N_SET_B_c_847_n N_A_2031_177#_c_1067_n 7.89191e-19 $X=11.05 $Y=0.72 $X2=0
+ $Y2=0
cc_611 N_SET_B_M1010_g N_A_2031_177#_M1019_g 0.015664f $X=11.185 $Y=2.785 $X2=0
+ $Y2=0
cc_612 SET_B N_A_2031_177#_M1019_g 0.0352632f $X=10.715 $Y=0.84 $X2=0 $Y2=0
cc_613 N_SET_B_c_847_n N_A_2031_177#_M1019_g 0.113812f $X=11.05 $Y=0.72 $X2=0
+ $Y2=0
cc_614 N_SET_B_c_892_p N_A_2031_177#_M1019_g 2.05814e-19 $X=11.05 $Y=0.72 $X2=0
+ $Y2=0
cc_615 SET_B N_A_1787_137#_M1015_d 0.00447341f $X=10.715 $Y=0.84 $X2=0 $Y2=0
cc_616 N_SET_B_c_842_n N_A_1787_137#_M1007_g 0.0337995f $X=11.15 $Y=1.85 $X2=0
+ $Y2=0
cc_617 N_SET_B_c_847_n N_A_1787_137#_M1007_g 0.0145705f $X=11.05 $Y=0.72 $X2=0
+ $Y2=0
cc_618 N_SET_B_M1010_g N_A_1787_137#_c_1138_n 0.0110694f $X=11.185 $Y=2.785
+ $X2=0 $Y2=0
cc_619 N_SET_B_M1010_g N_A_1787_137#_c_1139_n 0.0069264f $X=11.185 $Y=2.785
+ $X2=0 $Y2=0
cc_620 SET_B N_A_1787_137#_c_1131_n 0.046087f $X=10.715 $Y=0.84 $X2=0 $Y2=0
cc_621 N_SET_B_M1010_g N_A_1787_137#_c_1145_n 0.0212002f $X=11.185 $Y=2.785
+ $X2=0 $Y2=0
cc_622 N_SET_B_c_855_n N_A_1787_137#_c_1145_n 0.022144f $X=11.15 $Y=2.445 $X2=0
+ $Y2=0
cc_623 N_SET_B_c_855_n N_A_1787_137#_c_1147_n 0.0337995f $X=11.15 $Y=2.445 $X2=0
+ $Y2=0
cc_624 N_SET_B_c_843_n N_A_1787_137#_c_1148_n 0.00142931f $X=11.15 $Y=2.16 $X2=0
+ $Y2=0
cc_625 N_SET_B_M1010_g N_A_1787_137#_c_1148_n 0.0154736f $X=11.185 $Y=2.785
+ $X2=0 $Y2=0
cc_626 N_SET_B_c_855_n N_A_1787_137#_c_1148_n 0.0021381f $X=11.15 $Y=2.445 $X2=0
+ $Y2=0
cc_627 N_SET_B_M1026_g N_VPWR_c_1326_n 0.0413075f $X=7.12 $Y=2.855 $X2=0 $Y2=0
cc_628 N_SET_B_M1010_g N_VPWR_c_1329_n 0.0190393f $X=11.185 $Y=2.785 $X2=0 $Y2=0
cc_629 N_SET_B_c_855_n N_VPWR_c_1329_n 3.24599e-19 $X=11.15 $Y=2.445 $X2=0 $Y2=0
cc_630 N_SET_B_M1026_g N_VPWR_c_1338_n 0.00619492f $X=7.12 $Y=2.855 $X2=0 $Y2=0
cc_631 N_SET_B_M1010_g N_VPWR_c_1338_n 0.0098543f $X=11.185 $Y=2.785 $X2=0 $Y2=0
cc_632 N_SET_B_c_844_n N_VGND_c_1482_n 0.040448f $X=7.93 $Y=1.675 $X2=0 $Y2=0
cc_633 N_SET_B_c_845_n N_VGND_c_1482_n 0.0040588f $X=7.33 $Y=1.71 $X2=0 $Y2=0
cc_634 N_SET_B_c_868_n N_VGND_c_1482_n 0.0264004f $X=8.015 $Y=1.555 $X2=0 $Y2=0
cc_635 N_SET_B_c_884_p N_VGND_c_1482_n 0.0136768f $X=8.1 $Y=0.925 $X2=0 $Y2=0
cc_636 N_SET_B_c_849_n N_VGND_c_1482_n 0.052403f $X=7.182 $Y=1.545 $X2=0 $Y2=0
cc_637 N_SET_B_c_850_n N_VGND_c_1482_n 0.00893287f $X=8.512 $Y=0.782 $X2=0 $Y2=0
cc_638 N_SET_B_c_842_n N_VGND_c_1484_n 0.00211209f $X=11.15 $Y=1.85 $X2=0 $Y2=0
cc_639 N_SET_B_c_847_n N_VGND_c_1484_n 0.0368875f $X=11.05 $Y=0.72 $X2=0 $Y2=0
cc_640 N_SET_B_c_892_p N_VGND_c_1484_n 0.0370668f $X=11.05 $Y=0.72 $X2=0 $Y2=0
cc_641 N_SET_B_c_884_p N_VGND_c_1488_n 0.00795539f $X=8.1 $Y=0.925 $X2=0 $Y2=0
cc_642 SET_B N_VGND_c_1488_n 0.142368f $X=10.715 $Y=0.84 $X2=0 $Y2=0
cc_643 N_SET_B_c_847_n N_VGND_c_1488_n 0.016533f $X=11.05 $Y=0.72 $X2=0 $Y2=0
cc_644 N_SET_B_c_892_p N_VGND_c_1488_n 0.0217237f $X=11.05 $Y=0.72 $X2=0 $Y2=0
cc_645 N_SET_B_c_850_n N_VGND_c_1488_n 0.019044f $X=8.512 $Y=0.782 $X2=0 $Y2=0
cc_646 N_SET_B_c_886_p N_VGND_c_1488_n 0.00781261f $X=8.285 $Y=0.782 $X2=0 $Y2=0
cc_647 N_SET_B_c_850_n A_1645_137# 0.00392649f $X=8.512 $Y=0.782 $X2=0 $Y2=0
cc_648 N_A_798_107#_M1009_g N_VPWR_c_1323_n 0.00628462f $X=6.34 $Y=2.855 $X2=0
+ $Y2=0
cc_649 N_A_798_107#_c_940_n N_VPWR_c_1323_n 5.04822e-19 $X=6.215 $Y=2.515 $X2=0
+ $Y2=0
cc_650 N_A_798_107#_M1009_g N_VPWR_c_1326_n 5.51358e-19 $X=6.34 $Y=2.855 $X2=0
+ $Y2=0
cc_651 N_A_798_107#_c_951_n N_VPWR_c_1326_n 0.0516689f $X=7.995 $Y=2.465 $X2=0
+ $Y2=0
cc_652 N_A_798_107#_M1009_g N_VPWR_c_1338_n 0.0150362f $X=6.34 $Y=2.855 $X2=0
+ $Y2=0
cc_653 N_A_798_107#_c_951_n N_VPWR_c_1338_n 0.0187368f $X=7.995 $Y=2.465 $X2=0
+ $Y2=0
cc_654 N_A_798_107#_c_955_n N_VPWR_c_1338_n 0.00186757f $X=4.23 $Y=2.855 $X2=0
+ $Y2=0
cc_655 N_A_798_107#_c_941_n N_A_642_107#_c_1439_n 0.0127967f $X=4.15 $Y=0.745
+ $X2=0 $Y2=0
cc_656 N_A_798_107#_c_946_n N_A_642_107#_c_1439_n 0.00414964f $X=4.19 $Y=1.05
+ $X2=0 $Y2=0
cc_657 N_A_798_107#_c_935_n N_VGND_c_1480_n 0.00461416f $X=6.09 $Y=0.575 $X2=0
+ $Y2=0
cc_658 N_A_798_107#_c_941_n N_VGND_c_1480_n 0.00731308f $X=4.15 $Y=0.745 $X2=0
+ $Y2=0
cc_659 N_A_798_107#_c_943_n N_VGND_c_1480_n 0.0600343f $X=5.985 $Y=1.05 $X2=0
+ $Y2=0
cc_660 N_A_798_107#_c_944_n N_VGND_c_1480_n 0.0298877f $X=6.15 $Y=0.43 $X2=0
+ $Y2=0
cc_661 N_A_798_107#_M1025_g N_VGND_c_1482_n 0.00736387f $X=6.09 $Y=1.465 $X2=0
+ $Y2=0
cc_662 N_A_798_107#_c_938_n N_VGND_c_1482_n 0.0507198f $X=7.725 $Y=0.357 $X2=0
+ $Y2=0
cc_663 N_A_798_107#_M1013_g N_VGND_c_1482_n 0.0191693f $X=7.975 $Y=1.06 $X2=0
+ $Y2=0
cc_664 N_A_798_107#_c_943_n N_VGND_c_1482_n 0.00414505f $X=5.985 $Y=1.05 $X2=0
+ $Y2=0
cc_665 N_A_798_107#_c_944_n N_VGND_c_1482_n 0.0175474f $X=6.15 $Y=0.43 $X2=0
+ $Y2=0
cc_666 N_A_798_107#_M1006_d N_VGND_c_1488_n 0.00312781f $X=3.99 $Y=0.535 $X2=0
+ $Y2=0
cc_667 N_A_798_107#_c_935_n N_VGND_c_1488_n 0.00524234f $X=6.09 $Y=0.575 $X2=0
+ $Y2=0
cc_668 N_A_798_107#_M1025_g N_VGND_c_1488_n 0.00327716f $X=6.09 $Y=1.465 $X2=0
+ $Y2=0
cc_669 N_A_798_107#_c_938_n N_VGND_c_1488_n 0.0235916f $X=7.725 $Y=0.357 $X2=0
+ $Y2=0
cc_670 N_A_798_107#_M1013_g N_VGND_c_1488_n 0.0121523f $X=7.975 $Y=1.06 $X2=0
+ $Y2=0
cc_671 N_A_798_107#_c_941_n N_VGND_c_1488_n 0.0269684f $X=4.15 $Y=0.745 $X2=0
+ $Y2=0
cc_672 N_A_798_107#_c_943_n N_VGND_c_1488_n 0.0304736f $X=5.985 $Y=1.05 $X2=0
+ $Y2=0
cc_673 N_A_798_107#_c_944_n N_VGND_c_1488_n 0.0443781f $X=6.15 $Y=0.43 $X2=0
+ $Y2=0
cc_674 N_A_2031_177#_c_1055_n N_A_1787_137#_M1007_g 0.0305362f $X=12.12 $Y=1.74
+ $X2=0 $Y2=0
cc_675 N_A_2031_177#_c_1056_n N_A_1787_137#_M1007_g 0.0212471f $X=12.285
+ $Y=1.225 $X2=0 $Y2=0
cc_676 N_A_2031_177#_c_1057_n N_A_1787_137#_M1007_g 0.00580595f $X=12.475
+ $Y=3.005 $X2=0 $Y2=0
cc_677 N_A_2031_177#_c_1058_n N_A_1787_137#_M1007_g 0.00445567f $X=12.34 $Y=1.74
+ $X2=0 $Y2=0
cc_678 N_A_2031_177#_c_1057_n N_A_1787_137#_c_1133_n 0.0326321f $X=12.475
+ $Y=3.005 $X2=0 $Y2=0
cc_679 N_A_2031_177#_c_1056_n N_A_1787_137#_M1004_g 0.00202292f $X=12.285
+ $Y=1.225 $X2=7.44 $Y2=0.057
cc_680 N_A_2031_177#_c_1057_n N_A_1787_137#_M1004_g 6.9601e-19 $X=12.475
+ $Y=3.005 $X2=7.44 $Y2=0.057
cc_681 N_A_2031_177#_c_1058_n N_A_1787_137#_M1004_g 8.83584e-19 $X=12.34 $Y=1.74
+ $X2=7.44 $Y2=0.057
cc_682 N_A_2031_177#_c_1057_n N_A_1787_137#_c_1135_n 0.00139367f $X=12.475
+ $Y=3.005 $X2=0 $Y2=0
cc_683 N_A_2031_177#_c_1057_n N_A_1787_137#_c_1138_n 0.0175889f $X=12.475
+ $Y=3.005 $X2=0 $Y2=0
cc_684 N_A_2031_177#_c_1060_n N_A_1787_137#_c_1139_n 0.00701383f $X=11.425
+ $Y=3.38 $X2=0 $Y2=0
cc_685 N_A_2031_177#_c_1061_n N_A_1787_137#_c_1139_n 0.00272991f $X=11.465
+ $Y=3.505 $X2=0 $Y2=0
cc_686 N_A_2031_177#_c_1064_n N_A_1787_137#_c_1139_n 0.0336813f $X=12.39 $Y=3.09
+ $X2=0 $Y2=0
cc_687 N_A_2031_177#_M1019_g N_A_1787_137#_c_1131_n 0.00117754f $X=10.405
+ $Y=1.225 $X2=0 $Y2=0
cc_688 N_A_2031_177#_c_1067_n N_A_1787_137#_c_1144_n 0.013853f $X=10.47 $Y=1.71
+ $X2=0 $Y2=0
cc_689 N_A_2031_177#_M1019_g N_A_1787_137#_c_1144_n 0.00449134f $X=10.405
+ $Y=1.225 $X2=0 $Y2=0
cc_690 N_A_2031_177#_M1019_g N_A_1787_137#_c_1155_n 0.00100943f $X=10.405
+ $Y=1.225 $X2=0 $Y2=0
cc_691 N_A_2031_177#_c_1055_n N_A_1787_137#_c_1145_n 0.0237627f $X=12.12 $Y=1.74
+ $X2=0 $Y2=0
cc_692 N_A_2031_177#_c_1060_n N_A_1787_137#_c_1145_n 8.99742e-19 $X=11.425
+ $Y=3.38 $X2=0 $Y2=0
cc_693 N_A_2031_177#_c_1067_n N_A_1787_137#_c_1145_n 0.0235776f $X=10.47 $Y=1.71
+ $X2=0 $Y2=0
cc_694 N_A_2031_177#_M1019_g N_A_1787_137#_c_1145_n 0.0317626f $X=10.405
+ $Y=1.225 $X2=0 $Y2=0
cc_695 N_A_2031_177#_c_1064_n N_A_1787_137#_c_1147_n 4.3776e-19 $X=12.39 $Y=3.09
+ $X2=0 $Y2=0
cc_696 N_A_2031_177#_c_1058_n N_A_1787_137#_c_1147_n 0.00754709f $X=12.34
+ $Y=1.74 $X2=0 $Y2=0
cc_697 N_A_2031_177#_c_1055_n N_A_1787_137#_c_1148_n 0.03373f $X=12.12 $Y=1.74
+ $X2=0 $Y2=0
cc_698 N_A_2031_177#_c_1060_n N_A_1787_137#_c_1148_n 0.00933737f $X=11.425
+ $Y=3.38 $X2=0 $Y2=0
cc_699 N_A_2031_177#_c_1064_n N_A_1787_137#_c_1148_n 0.0352834f $X=12.39 $Y=3.09
+ $X2=0 $Y2=0
cc_700 N_A_2031_177#_c_1057_n N_A_1787_137#_c_1148_n 0.052697f $X=12.475
+ $Y=3.005 $X2=0 $Y2=0
cc_701 N_A_2031_177#_c_1058_n N_A_1787_137#_c_1148_n 0.00756206f $X=12.34
+ $Y=1.74 $X2=0 $Y2=0
cc_702 N_A_2031_177#_c_1056_n N_A_2553_203#_c_1257_n 0.0283781f $X=12.285
+ $Y=1.225 $X2=7.44 $Y2=0
cc_703 N_A_2031_177#_c_1056_n N_A_2553_203#_c_1258_n 0.00777948f $X=12.285
+ $Y=1.225 $X2=0 $Y2=0
cc_704 N_A_2031_177#_c_1057_n N_A_2553_203#_c_1258_n 0.018479f $X=12.475
+ $Y=3.005 $X2=0 $Y2=0
cc_705 N_A_2031_177#_c_1058_n N_A_2553_203#_c_1258_n 0.00969603f $X=12.34
+ $Y=1.74 $X2=0 $Y2=0
cc_706 N_A_2031_177#_c_1064_n N_A_2553_203#_c_1266_n 0.00954499f $X=12.39
+ $Y=3.09 $X2=0 $Y2=0
cc_707 N_A_2031_177#_c_1057_n N_A_2553_203#_c_1266_n 0.0301401f $X=12.475
+ $Y=3.005 $X2=0 $Y2=0
cc_708 N_A_2031_177#_c_1057_n N_A_2553_203#_c_1276_n 0.00809674f $X=12.475
+ $Y=3.005 $X2=0 $Y2=0
cc_709 N_A_2031_177#_c_1060_n N_VPWR_c_1329_n 0.0176622f $X=11.425 $Y=3.38 $X2=0
+ $Y2=0
cc_710 N_A_2031_177#_c_1061_n N_VPWR_c_1329_n 0.0129151f $X=11.465 $Y=3.505
+ $X2=0 $Y2=0
cc_711 N_A_2031_177#_M1019_g N_VPWR_c_1329_n 0.044716f $X=10.405 $Y=1.225 $X2=0
+ $Y2=0
cc_712 N_A_2031_177#_c_1061_n N_VPWR_c_1332_n 0.0172607f $X=11.465 $Y=3.505
+ $X2=0 $Y2=0
cc_713 N_A_2031_177#_c_1064_n N_VPWR_c_1332_n 0.0523742f $X=12.39 $Y=3.09 $X2=0
+ $Y2=0
cc_714 N_A_2031_177#_M1012_s N_VPWR_c_1338_n 0.00174254f $X=11.32 $Y=3.295 $X2=0
+ $Y2=0
cc_715 N_A_2031_177#_c_1061_n N_VPWR_c_1338_n 0.0255076f $X=11.465 $Y=3.505
+ $X2=0 $Y2=0
cc_716 N_A_2031_177#_c_1064_n N_VPWR_c_1338_n 0.0129125f $X=12.39 $Y=3.09 $X2=0
+ $Y2=0
cc_717 N_A_2031_177#_c_1055_n N_VGND_c_1484_n 0.0448467f $X=12.12 $Y=1.74 $X2=0
+ $Y2=0
cc_718 N_A_2031_177#_c_1056_n N_VGND_c_1484_n 0.0359178f $X=12.285 $Y=1.225
+ $X2=0 $Y2=0
cc_719 N_A_2031_177#_M1019_g N_VGND_c_1484_n 0.00136572f $X=10.405 $Y=1.225
+ $X2=0 $Y2=0
cc_720 N_A_2031_177#_c_1056_n N_VGND_c_1488_n 0.0156654f $X=12.285 $Y=1.225
+ $X2=0 $Y2=0
cc_721 N_A_1787_137#_M1004_g N_A_2553_203#_M1008_g 0.0145528f $X=13.3 $Y=1.225
+ $X2=0 $Y2=0
cc_722 N_A_1787_137#_c_1142_n N_A_2553_203#_M1001_g 0.0192935f $X=13.32 $Y=2.235
+ $X2=0 $Y2=0
cc_723 N_A_1787_137#_M1004_g N_A_2553_203#_c_1256_n 0.0197432f $X=13.3 $Y=1.225
+ $X2=0 $Y2=0
cc_724 N_A_1787_137#_M1007_g N_A_2553_203#_c_1257_n 0.0011881f $X=11.895
+ $Y=1.225 $X2=7.44 $Y2=0
cc_725 N_A_1787_137#_M1004_g N_A_2553_203#_c_1257_n 0.00714064f $X=13.3 $Y=1.225
+ $X2=7.44 $Y2=0
cc_726 N_A_1787_137#_c_1133_n N_A_2553_203#_c_1258_n 0.0109915f $X=13.05
+ $Y=2.235 $X2=0 $Y2=0
cc_727 N_A_1787_137#_M1004_g N_A_2553_203#_c_1258_n 0.0319553f $X=13.3 $Y=1.225
+ $X2=0 $Y2=0
cc_728 N_A_1787_137#_c_1142_n N_A_2553_203#_c_1258_n 0.0107883f $X=13.32
+ $Y=2.235 $X2=0 $Y2=0
cc_729 N_A_1787_137#_c_1133_n N_A_2553_203#_c_1266_n 0.00658014f $X=13.05
+ $Y=2.235 $X2=0 $Y2=0
cc_730 N_A_1787_137#_c_1135_n N_A_2553_203#_c_1266_n 0.0212129f $X=13.34
+ $Y=2.485 $X2=0 $Y2=0
cc_731 N_A_1787_137#_c_1139_n N_A_2553_203#_c_1266_n 0.00583206f $X=12.027
+ $Y=3.185 $X2=0 $Y2=0
cc_732 N_A_1787_137#_c_1142_n N_A_2553_203#_c_1266_n 0.00440038f $X=13.32
+ $Y=2.235 $X2=0 $Y2=0
cc_733 N_A_1787_137#_c_1142_n N_A_2553_203#_c_1268_n 0.0424926f $X=13.32
+ $Y=2.235 $X2=0 $Y2=0
cc_734 N_A_1787_137#_M1004_g N_A_2553_203#_c_1290_n 0.00172049f $X=13.3 $Y=1.225
+ $X2=0 $Y2=0
cc_735 N_A_1787_137#_c_1142_n N_A_2553_203#_c_1290_n 0.00169086f $X=13.32
+ $Y=2.235 $X2=0 $Y2=0
cc_736 N_A_1787_137#_c_1142_n N_A_2553_203#_c_1259_n 0.0236716f $X=13.32
+ $Y=2.235 $X2=0 $Y2=0
cc_737 N_A_1787_137#_c_1133_n N_A_2553_203#_c_1260_n 0.00371049f $X=13.05
+ $Y=2.235 $X2=0 $Y2=0
cc_738 N_A_1787_137#_M1004_g N_A_2553_203#_c_1260_n 0.00386717f $X=13.3 $Y=1.225
+ $X2=0 $Y2=0
cc_739 N_A_1787_137#_c_1133_n N_A_2553_203#_c_1276_n 0.00633656f $X=13.05
+ $Y=2.235 $X2=0 $Y2=0
cc_740 N_A_1787_137#_c_1142_n N_A_2553_203#_c_1276_n 0.00311713f $X=13.32
+ $Y=2.235 $X2=0 $Y2=0
cc_741 N_A_1787_137#_c_1143_n N_VPWR_c_1329_n 0.0200192f $X=9.49 $Y=3.22 $X2=0
+ $Y2=0
cc_742 N_A_1787_137#_c_1155_n N_VPWR_c_1329_n 0.0163218f $X=9.575 $Y=3.025 $X2=0
+ $Y2=0
cc_743 N_A_1787_137#_c_1145_n N_VPWR_c_1329_n 0.0643102f $X=11.41 $Y=2.4 $X2=0
+ $Y2=0
cc_744 N_A_1787_137#_c_1148_n N_VPWR_c_1329_n 0.00581004f $X=11.81 $Y=2.4 $X2=0
+ $Y2=0
cc_745 N_A_1787_137#_c_1135_n N_VPWR_c_1332_n 0.00232371f $X=13.34 $Y=2.485
+ $X2=0 $Y2=0
cc_746 N_A_1787_137#_c_1139_n N_VPWR_c_1332_n 0.0340593f $X=12.027 $Y=3.185
+ $X2=0 $Y2=0
cc_747 N_A_1787_137#_c_1135_n N_VPWR_c_1335_n 0.0622105f $X=13.34 $Y=2.485 $X2=0
+ $Y2=0
cc_748 N_A_1787_137#_M1014_d N_VPWR_c_1338_n 0.00347236f $X=8.975 $Y=2.575 $X2=0
+ $Y2=0
cc_749 N_A_1787_137#_c_1135_n N_VPWR_c_1338_n 0.0116796f $X=13.34 $Y=2.485 $X2=0
+ $Y2=0
cc_750 N_A_1787_137#_c_1139_n N_VPWR_c_1338_n 0.00387056f $X=12.027 $Y=3.185
+ $X2=0 $Y2=0
cc_751 N_A_1787_137#_c_1143_n N_VPWR_c_1338_n 0.0211883f $X=9.49 $Y=3.22 $X2=0
+ $Y2=0
cc_752 N_A_1787_137#_c_1148_n N_VPWR_c_1338_n 8.18759e-19 $X=11.81 $Y=2.4 $X2=0
+ $Y2=0
cc_753 N_A_1787_137#_M1007_g N_VGND_c_1484_n 0.0405294f $X=11.895 $Y=1.225 $X2=0
+ $Y2=0
cc_754 N_A_1787_137#_M1004_g N_VGND_c_1486_n 0.0590094f $X=13.3 $Y=1.225 $X2=0
+ $Y2=0
cc_755 N_A_1787_137#_c_1142_n N_VGND_c_1486_n 0.00135541f $X=13.32 $Y=2.235
+ $X2=0 $Y2=0
cc_756 N_A_1787_137#_M1007_g N_VGND_c_1488_n 0.00645752f $X=11.895 $Y=1.225
+ $X2=0 $Y2=0
cc_757 N_A_1787_137#_M1004_g N_VGND_c_1488_n 0.00615856f $X=13.3 $Y=1.225 $X2=0
+ $Y2=0
cc_758 N_A_1787_137#_c_1131_n N_VGND_c_1488_n 0.00228656f $X=9.49 $Y=1.332 $X2=0
+ $Y2=0
cc_759 N_A_2553_203#_c_1266_n N_VPWR_c_1332_n 7.35252e-19 $X=12.95 $Y=2.74 $X2=0
+ $Y2=0
cc_760 N_A_2553_203#_M1001_g N_VPWR_c_1335_n 0.0530997f $X=14.215 $Y=3.095 $X2=0
+ $Y2=0
cc_761 N_A_2553_203#_c_1264_n N_VPWR_c_1335_n 0.00220765f $X=14.177 $Y=2.465
+ $X2=0 $Y2=0
cc_762 N_A_2553_203#_c_1266_n N_VPWR_c_1335_n 0.0587722f $X=12.95 $Y=2.74 $X2=0
+ $Y2=0
cc_763 N_A_2553_203#_c_1268_n N_VPWR_c_1335_n 0.0739983f $X=13.91 $Y=2.31 $X2=0
+ $Y2=0
cc_764 N_A_2553_203#_M1001_g N_VPWR_c_1338_n 0.0148289f $X=14.215 $Y=3.095 $X2=0
+ $Y2=0
cc_765 N_A_2553_203#_c_1266_n N_VPWR_c_1338_n 0.0106225f $X=12.95 $Y=2.74 $X2=0
+ $Y2=0
cc_766 N_A_2553_203#_M1008_g N_Q_c_1461_n 0.0253281f $X=14.195 $Y=1.06 $X2=0
+ $Y2=0
cc_767 N_A_2553_203#_M1001_g N_Q_c_1461_n 0.0268854f $X=14.215 $Y=3.095 $X2=0
+ $Y2=0
cc_768 N_A_2553_203#_c_1256_n N_Q_c_1461_n 0.0166146f $X=14.177 $Y=1.852 $X2=0
+ $Y2=0
cc_769 N_A_2553_203#_c_1264_n N_Q_c_1461_n 0.0132894f $X=14.177 $Y=2.465 $X2=0
+ $Y2=0
cc_770 N_A_2553_203#_c_1268_n N_Q_c_1461_n 0.0130141f $X=13.91 $Y=2.31 $X2=0
+ $Y2=0
cc_771 N_A_2553_203#_c_1290_n N_Q_c_1461_n 0.0358236f $X=14.075 $Y=1.89 $X2=0
+ $Y2=0
cc_772 N_A_2553_203#_c_1259_n N_Q_c_1461_n 0.0125969f $X=14.075 $Y=1.89 $X2=0
+ $Y2=0
cc_773 N_A_2553_203#_M1008_g N_VGND_c_1486_n 0.053118f $X=14.195 $Y=1.06 $X2=0
+ $Y2=0
cc_774 N_A_2553_203#_c_1256_n N_VGND_c_1486_n 0.00217835f $X=14.177 $Y=1.852
+ $X2=0 $Y2=0
cc_775 N_A_2553_203#_c_1257_n N_VGND_c_1486_n 0.0379082f $X=12.91 $Y=1.225 $X2=0
+ $Y2=0
cc_776 N_A_2553_203#_c_1290_n N_VGND_c_1486_n 0.0183072f $X=14.075 $Y=1.89 $X2=0
+ $Y2=0
cc_777 N_A_2553_203#_M1008_g N_VGND_c_1488_n 0.0143581f $X=14.195 $Y=1.06 $X2=0
+ $Y2=0
cc_778 N_A_2553_203#_c_1257_n N_VGND_c_1488_n 0.0154896f $X=12.91 $Y=1.225 $X2=0
+ $Y2=0
cc_779 N_VPWR_c_1338_n N_A_642_107#_c_1438_n 9.76264e-19 $X=14.125 $Y=3.59
+ $X2=0.24 $Y2=4.07
cc_780 N_VPWR_c_1338_n A_1653_515# 0.00875788f $X=14.125 $Y=3.59 $X2=0 $Y2=3.985
cc_781 N_VPWR_c_1329_n A_1989_515# 0.00476837f $X=10.795 $Y=2.81 $X2=0 $Y2=3.985
cc_782 N_VPWR_c_1335_n N_Q_c_1461_n 0.0767481f $X=13.825 $Y=2.74 $X2=7.44
+ $Y2=4.07
cc_783 N_VPWR_c_1338_n N_Q_c_1461_n 0.037159f $X=14.125 $Y=3.59 $X2=7.44
+ $Y2=4.07
cc_784 N_A_642_107#_c_1439_n N_VGND_c_1478_n 0.0356375f $X=3.35 $Y=0.745 $X2=0
+ $Y2=0
cc_785 N_A_642_107#_c_1439_n N_VGND_c_1488_n 0.0332933f $X=3.35 $Y=0.745 $X2=0
+ $Y2=0
cc_786 N_Q_c_1461_n N_VGND_c_1486_n 0.0548845f $X=14.585 $Y=0.81 $X2=0 $Y2=0
cc_787 N_Q_c_1461_n N_VGND_c_1488_n 0.0158019f $X=14.585 $Y=0.81 $X2=0 $Y2=0
cc_788 N_VGND_c_1480_n A_958_107# 0.00424569f $X=5.69 $Y=0.48 $X2=0 $Y2=0
cc_789 N_VGND_c_1488_n A_958_107# 6.9132e-19 $X=14.09 $Y=0.48 $X2=0 $Y2=0
