* File: sky130_fd_sc_hvl__nor3_1.spice
* Created: Wed Sep  2 09:08:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__nor3_1.pex.spice"
.subckt sky130_fd_sc_hvl__nor3_1  VNB VPB A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_A_M1003_g N_VGND_M1003_s N_VNB_M1003_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000 SB=250002
+ A=0.375 P=2.5 MULT=1
MM1005 N_VGND_M1005_d N_B_M1005_g N_Y_M1003_d N_VNB_M1003_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250001 SB=250001
+ A=0.375 P=2.5 MULT=1
MM1004 N_Y_M1004_d N_C_M1004_g N_VGND_M1005_d N_VNB_M1003_b NHV L=0.5 W=0.75
+ AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250002 SB=250000
+ A=0.375 P=2.5 MULT=1
MM1000 A_205_443# N_A_M1000_g N_VPWR_M1000_s N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.1575 AS=0.4275 PD=1.71 PS=3.57 NRD=6.3603 NRS=0 M=1 R=3 SA=250000
+ SB=250001 A=0.75 P=4 MULT=1
MM1001 A_347_443# N_B_M1001_g A_205_443# N_VPB_M1000_b PHV L=0.5 W=1.5 AD=0.1575
+ AS=0.1575 PD=1.71 PS=1.71 NRD=6.3603 NRS=6.3603 M=1 R=3 SA=250001 SB=250001
+ A=0.75 P=4 MULT=1
MM1002 N_Y_M1002_d N_C_M1002_g A_347_443# N_VPB_M1000_b PHV L=0.5 W=1.5
+ AD=0.4275 AS=0.1575 PD=3.57 PS=1.71 NRD=0 NRS=6.3603 M=1 R=3 SA=250001
+ SB=250000 A=0.75 P=4 MULT=1
DX6_noxref N_VNB_M1003_b N_VPB_M1000_b NWDIODE A=10.452 P=13.24
*
.include "sky130_fd_sc_hvl__nor3_1.pxi.spice"
*
.ends
*
*
