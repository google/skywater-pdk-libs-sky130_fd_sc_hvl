* File: sky130_fd_sc_hvl__o22ai_1.pex.spice
* Created: Wed Sep  2 09:09:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__O22AI_1%VNB 5 7 11 25
c28 5 0 9.86576e-20 $X=-0.33 $Y=-0.265
r29 7 25 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=0.057
+ $X2=1.92 $Y2=0.058
r30 7 11 0.00185547 $w=3.84e-06 $l=5.7e-08 $layer=MET1_cond $X=1.92 $Y=0.057
+ $X2=1.92 $Y2=0
r31 5 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r32 5 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__O22AI_1%VPB 4 6 14 21
r31 10 21 0.00185547 $w=3.84e-06 $l=5.7e-08 $layer=MET1_cond $X=1.92 $Y=4.07
+ $X2=1.92 $Y2=4.013
r32 10 14 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=4.07
+ $X2=3.6 $Y2=4.07
r33 9 14 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=3.6
+ $Y2=4.07
r34 9 10 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r35 6 21 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=4.012
+ $X2=1.92 $Y2=4.013
r36 4 14 45.5 $w=1.7e-07 $l=3.64225e-06 $layer=licon1_NTAP_notbjt $count=4 $X=0
+ $Y=3.985 $X2=3.6 $Y2=4.07
r37 4 9 45.5 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=4 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__O22AI_1%B1 1 3 6 8 12 15
c29 6 0 4.74589e-20 $X=0.785 $Y=2.965
c30 1 0 9.86576e-20 $X=0.715 $Y=1.425
r31 14 15 7.49041 $w=5e-07 $l=7e-08 $layer=POLY_cond $X=0.715 $Y=1.675 $X2=0.785
+ $Y2=1.675
r32 11 14 35.3119 $w=5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.385 $Y=1.675
+ $X2=0.715 $Y2=1.675
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.7 $X2=0.385 $Y2=1.7
r34 8 12 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.7
+ $X2=0.385 $Y2=1.7
r35 4 15 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.785 $Y=1.925
+ $X2=0.785 $Y2=1.675
r36 4 6 111.286 $w=5e-07 $l=1.04e-06 $layer=POLY_cond $X=0.785 $Y=1.925
+ $X2=0.785 $Y2=2.965
r37 1 14 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.715 $Y=1.425
+ $X2=0.715 $Y2=1.675
r38 1 3 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.715 $Y=1.425 $X2=0.715
+ $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_HVL__O22AI_1%B2 1 4 8 10
c31 8 0 6.31983e-20 $X=1.43 $Y=1.645
r32 7 10 141.248 $w=5e-07 $l=1.32e-06 $layer=POLY_cond $X=1.495 $Y=1.645
+ $X2=1.495 $Y2=2.965
r33 7 8 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.43
+ $Y=1.645 $X2=1.43 $Y2=1.645
r34 4 7 75.4392 $w=5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.495 $Y=0.94 $X2=1.495
+ $Y2=1.645
r35 1 8 12.3285 $w=2.13e-07 $l=2.3e-07 $layer=LI1_cond $X=1.2 $Y=1.642 $X2=1.43
+ $Y2=1.642
.ends

.subckt PM_SKY130_FD_SC_HVL__O22AI_1%A2 3 7 8 11 14
c34 3 0 6.31983e-20 $X=2.275 $Y=0.94
r35 11 14 21.0588 $w=5.75e-07 $l=2.15e-07 $layer=POLY_cond $X=2.312 $Y=1.89
+ $X2=2.312 $Y2=2.105
r36 11 13 27.5722 $w=5.75e-07 $l=2.85e-07 $layer=POLY_cond $X=2.312 $Y=1.89
+ $X2=2.312 $Y2=1.605
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.89 $X2=2.415 $Y2=1.89
r38 8 12 8.23174 $w=3.13e-07 $l=2.25e-07 $layer=LI1_cond $X=2.64 $Y=1.962
+ $X2=2.415 $Y2=1.962
r39 7 14 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.35 $Y=2.965 $X2=2.35
+ $Y2=2.105
r40 3 13 71.1589 $w=5e-07 $l=6.65e-07 $layer=POLY_cond $X=2.275 $Y=0.94
+ $X2=2.275 $Y2=1.605
.ends

.subckt PM_SKY130_FD_SC_HVL__O22AI_1%A1 3 7 9 10 14
r26 14 17 19.0549 $w=5.95e-07 $l=1.95e-07 $layer=POLY_cond $X=3.107 $Y=1.89
+ $X2=3.107 $Y2=2.085
r27 14 16 41.5351 $w=5.95e-07 $l=4.45e-07 $layer=POLY_cond $X=3.107 $Y=1.89
+ $X2=3.107 $Y2=1.445
r28 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.21
+ $Y=1.89 $X2=3.21 $Y2=1.89
r29 10 15 14.2683 $w=3.13e-07 $l=3.9e-07 $layer=LI1_cond $X=3.6 $Y=1.962
+ $X2=3.21 $Y2=1.962
r30 9 15 3.29269 $w=3.13e-07 $l=9e-08 $layer=LI1_cond $X=3.12 $Y=1.962 $X2=3.21
+ $Y2=1.962
r31 7 16 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.155 $Y=0.94 $X2=3.155
+ $Y2=1.445
r32 3 17 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.06 $Y=2.965 $X2=3.06
+ $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_HVL__O22AI_1%VPWR 1 2 7 10 20 27
r35 24 27 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=2.42 $Y=3.63
+ $X2=3.5 $Y2=3.63
r36 23 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.5 $Y=3.59 $X2=3.5
+ $Y2=3.59
r37 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.42 $Y=3.59
+ $X2=2.42 $Y2=3.59
r38 20 23 11.2221 $w=1.308e-06 $l=1.205e-06 $layer=LI1_cond $X=2.96 $Y=2.385
+ $X2=2.96 $Y2=3.59
r39 14 17 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=0.18 $Y=3.63
+ $X2=1.26 $Y2=3.63
r40 13 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.26 $Y=3.59
+ $X2=1.26 $Y2=3.59
r41 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.18 $Y=3.59
+ $X2=0.18 $Y2=3.59
r42 10 13 11.9084 $w=1.253e-06 $l=1.225e-06 $layer=LI1_cond $X=0.717 $Y=2.365
+ $X2=0.717 $Y2=3.59
r43 7 24 0.191953 $w=3.7e-07 $l=5e-07 $layer=MET1_cond $X=1.92 $Y=3.63 $X2=2.42
+ $Y2=3.63
r44 7 17 0.253378 $w=3.7e-07 $l=6.6e-07 $layer=MET1_cond $X=1.92 $Y=3.63
+ $X2=1.26 $Y2=3.63
r45 2 23 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=3.31
+ $Y=2.215 $X2=3.45 $Y2=3.59
r46 2 20 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=3.31
+ $Y=2.215 $X2=3.45 $Y2=2.385
r47 1 13 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.25
+ $Y=2.215 $X2=0.395 $Y2=3.59
r48 1 10 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.25
+ $Y=2.215 $X2=0.395 $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_HVL__O22AI_1%Y 1 2 8 9 10 13 16 19 20 21 22 28 40
c45 8 0 4.74589e-20 $X=0.82 $Y=1.93
r46 44 45 7.80118 $w=5.18e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=3.175
+ $X2=1.785 $Y2=3.26
r47 28 40 1.40589 $w=5.2e-07 $l=3e-08 $layer=LI1_cond $X=1.785 $Y=2.435
+ $X2=1.785 $Y2=2.405
r48 22 44 0.690045 $w=5.18e-07 $l=3e-08 $layer=LI1_cond $X=1.785 $Y=3.145
+ $X2=1.785 $Y2=3.175
r49 22 29 3.33522 $w=5.18e-07 $l=1.45e-07 $layer=LI1_cond $X=1.785 $Y=3.145
+ $X2=1.785 $Y2=3
r50 21 29 5.17534 $w=5.18e-07 $l=2.25e-07 $layer=LI1_cond $X=1.785 $Y=2.775
+ $X2=1.785 $Y2=3
r51 20 40 0.858291 $w=3.98e-07 $l=2.8e-08 $layer=LI1_cond $X=1.785 $Y=2.377
+ $X2=1.785 $Y2=2.405
r52 20 37 1.13417 $w=3.98e-07 $l=3.7e-08 $layer=LI1_cond $X=1.785 $Y=2.377
+ $X2=1.785 $Y2=2.34
r53 20 21 7.19947 $w=5.18e-07 $l=3.13e-07 $layer=LI1_cond $X=1.785 $Y=2.462
+ $X2=1.785 $Y2=2.775
r54 20 28 0.621041 $w=5.18e-07 $l=2.7e-08 $layer=LI1_cond $X=1.785 $Y=2.462
+ $X2=1.785 $Y2=2.435
r55 19 37 9.34925 $w=3.98e-07 $l=3.05e-07 $layer=LI1_cond $X=1.785 $Y=2.035
+ $X2=1.785 $Y2=2.34
r56 19 33 0.613065 $w=3.98e-07 $l=2e-08 $layer=LI1_cond $X=1.785 $Y=2.035
+ $X2=1.785 $Y2=2.015
r57 16 18 20.6908 $w=5.33e-07 $l=6.55e-07 $layer=LI1_cond $X=1.002 $Y=0.7
+ $X2=1.002 $Y2=1.355
r58 13 45 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.96 $Y=3.59
+ $X2=1.96 $Y2=3.26
r59 9 33 5.74796 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=1.525 $Y=2.015
+ $X2=1.785 $Y2=2.015
r60 9 10 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.525 $Y=2.015
+ $X2=0.905 $Y2=2.015
r61 8 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.82 $Y=1.93
+ $X2=0.905 $Y2=2.015
r62 8 18 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.82 $Y=1.93
+ $X2=0.82 $Y2=1.355
r63 2 44 400 $w=1.7e-07 $l=1.06207e-06 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=2.215 $X2=1.96 $Y2=3.175
r64 2 37 400 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=2.215 $X2=1.96 $Y2=2.34
r65 2 13 600 $w=1.7e-07 $l=1.4786e-06 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=2.215 $X2=1.96 $Y2=3.59
r66 1 16 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=0.565 $X2=1.105 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__O22AI_1%A_36_113# 1 2 3 12 14 15 19 20 21 24
r43 22 24 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=3.545 $Y=1.455
+ $X2=3.545 $Y2=0.69
r44 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.42 $Y=1.54
+ $X2=3.545 $Y2=1.455
r45 20 21 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=3.42 $Y=1.54
+ $X2=1.97 $Y2=1.54
r46 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.885 $Y=1.455
+ $X2=1.97 $Y2=1.54
r47 17 19 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.885 $Y=1.455
+ $X2=1.885 $Y2=0.69
r48 16 19 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.885 $Y=0.435
+ $X2=1.885 $Y2=0.69
r49 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.8 $Y=0.35
+ $X2=1.885 $Y2=0.435
r50 14 15 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=1.8 $Y=0.35
+ $X2=0.49 $Y2=0.35
r51 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.325 $Y=0.435
+ $X2=0.49 $Y2=0.35
r52 10 12 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.325 $Y=0.435
+ $X2=0.325 $Y2=0.69
r53 3 24 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.565 $X2=3.545 $Y2=0.69
r54 2 19 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.745
+ $Y=0.565 $X2=1.885 $Y2=0.69
r55 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.18
+ $Y=0.565 $X2=0.325 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HVL__O22AI_1%VGND 1 4 7 11
r24 8 11 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.285 $Y=0.44
+ $X2=3.005 $Y2=0.44
r25 7 13 2.32909 $w=1.098e-06 $l=2.1e-07 $layer=LI1_cond $X=2.7 $Y=0.48 $X2=2.7
+ $Y2=0.69
r26 7 11 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.005 $Y=0.48
+ $X2=3.005 $Y2=0.48
r27 7 8 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.285 $Y=0.48
+ $X2=2.285 $Y2=0.48
r28 4 8 0.140125 $w=3.7e-07 $l=3.65e-07 $layer=MET1_cond $X=1.92 $Y=0.44
+ $X2=2.285 $Y2=0.44
r29 1 13 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.525
+ $Y=0.565 $X2=2.665 $Y2=0.69
.ends

