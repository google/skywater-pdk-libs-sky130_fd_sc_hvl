* File: sky130_fd_sc_hvl__decap_8.spice
* Created: Fri Aug 28 09:33:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__decap_8.pex.spice"
.subckt sky130_fd_sc_hvl__decap_8  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_s N_VPWR_M1001_g N_VGND_M1001_s N_VNB_M1001_b NHV L=1 W=0.75
+ AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=0.75 SA=500000 SB=500001
+ A=0.75 P=3.5 MULT=1
MM1003 N_VGND_M1001_s N_VPWR_M1003_g N_VGND_M1001_s N_VNB_M1001_b NHV L=1 W=0.75
+ AD=0.21375 AS=0.105 PD=2.07 PS=1.03 NRD=0 NRS=0 M=1 R=0.75 SA=500001 SB=500000
+ A=0.75 P=3.5 MULT=1
MM1000 N_VPWR_M1000_s N_VGND_M1000_g N_VPWR_M1000_s N_VPB_M1000_b PHV L=1 W=1
+ AD=0.14 AS=0.275 PD=1.28 PS=2.55 NRD=0 NRS=1.8909 M=1 R=1 SA=500000 SB=500001
+ A=1 P=4 MULT=1
MM1002 N_VPWR_M1000_s N_VGND_M1002_g N_VPWR_M1000_s N_VPB_M1000_b PHV L=1 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=1 SA=500001 SB=500000 A=1
+ P=4 MULT=1
DX4_noxref N_VNB_M1001_b N_VPB_M1000_b NWDIODE A=11.7 P=14.2
*
.include "sky130_fd_sc_hvl__decap_8.pxi.spice"
*
.ends
*
*
