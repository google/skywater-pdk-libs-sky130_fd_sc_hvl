# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hvl__buf_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  17.76000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  6.750000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.220000 1.580000 4.630000 1.815000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  5.040000 ;
    ANTENNAGATEAREA  6.750000 ;
    ANTENNAPARTIALMETALSIDEAREA  0.336000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  5.590000 2.290000  5.880000 2.320000 ;
        RECT  5.590000 2.320000 16.800000 2.490000 ;
        RECT  5.590000 2.490000  5.880000 2.520000 ;
        RECT  7.150000 2.290000  7.440000 2.320000 ;
        RECT  7.150000 2.490000  7.440000 2.520000 ;
        RECT  8.710000 2.290000  9.000000 2.320000 ;
        RECT  8.710000 2.490000  9.000000 2.520000 ;
        RECT 10.270000 2.290000 10.560000 2.320000 ;
        RECT 10.270000 2.490000 10.560000 2.520000 ;
        RECT 11.830000 2.290000 12.120000 2.320000 ;
        RECT 11.830000 2.490000 12.120000 2.520000 ;
        RECT 13.390000 2.290000 13.680000 2.320000 ;
        RECT 13.390000 2.490000 13.680000 2.520000 ;
        RECT 14.950000 2.290000 15.240000 2.320000 ;
        RECT 14.950000 2.490000 15.240000 2.520000 ;
        RECT 16.510000 2.290000 16.800000 2.320000 ;
        RECT 16.510000 2.490000 16.800000 2.520000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 17.760000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 17.760000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 17.760000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 17.760000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 17.760000 0.085000 ;
      RECT  0.000000  3.985000 17.760000 4.155000 ;
      RECT  0.110000  0.425000  0.645000 1.410000 ;
      RECT  0.110000  2.175000  0.680000 3.755000 ;
      RECT  0.815000  0.755000  1.170000 1.195000 ;
      RECT  0.815000  1.195000  5.350000 1.410000 ;
      RECT  0.850000  1.985000  5.350000 2.265000 ;
      RECT  0.850000  2.265000  1.160000 3.755000 ;
      RECT  1.340000  0.415000  2.230000 1.025000 ;
      RECT  1.340000  2.445000  2.230000 3.675000 ;
      RECT  2.400000  0.730000  2.790000 1.195000 ;
      RECT  2.400000  2.265000  2.710000 3.755000 ;
      RECT  2.880000  2.445000  3.770000 3.675000 ;
      RECT  2.960000  0.425000  3.855000 1.025000 ;
      RECT  3.940000  2.265000  4.290000 3.755000 ;
      RECT  4.025000  0.730000  4.270000 1.195000 ;
      RECT  4.440000  0.425000  5.330000 1.025000 ;
      RECT  4.460000  2.445000  5.350000 3.675000 ;
      RECT  4.800000  1.410000  5.350000 1.985000 ;
      RECT  5.570000  0.790000  5.900000 3.755000 ;
      RECT  6.070000  0.425000  6.960000 1.395000 ;
      RECT  6.070000  2.175000  6.960000 3.755000 ;
      RECT  6.160000  1.565000  6.830000 1.895000 ;
      RECT  7.130000  0.790000  7.460000 3.755000 ;
      RECT  7.630000  0.425000  8.520000 1.395000 ;
      RECT  7.630000  2.175000  8.520000 3.755000 ;
      RECT  7.720000  1.565000  8.390000 1.895000 ;
      RECT  8.690000  0.790000  9.020000 3.755000 ;
      RECT  9.190000  0.425000 10.080000 1.395000 ;
      RECT  9.190000  2.175000 10.080000 3.755000 ;
      RECT  9.280000  1.565000  9.950000 1.895000 ;
      RECT 10.250000  0.790000 10.580000 3.755000 ;
      RECT 10.750000  0.425000 11.640000 1.395000 ;
      RECT 10.750000  2.175000 11.640000 3.755000 ;
      RECT 10.840000  1.565000 11.510000 1.895000 ;
      RECT 11.810000  0.790000 12.140000 3.755000 ;
      RECT 12.310000  0.425000 13.200000 1.395000 ;
      RECT 12.310000  2.175000 13.200000 3.755000 ;
      RECT 12.400000  1.565000 13.070000 1.895000 ;
      RECT 13.370000  0.790000 13.700000 3.755000 ;
      RECT 13.870000  0.425000 14.760000 1.395000 ;
      RECT 13.870000  2.175000 14.760000 3.755000 ;
      RECT 13.960000  1.565000 14.630000 1.895000 ;
      RECT 14.930000  0.790000 15.260000 3.755000 ;
      RECT 15.430000  0.425000 16.320000 1.395000 ;
      RECT 15.430000  2.175000 16.320000 3.755000 ;
      RECT 15.520000  1.565000 16.190000 1.895000 ;
      RECT 16.490000  0.790000 16.900000 3.755000 ;
      RECT 17.070000  0.425000 17.600000 1.495000 ;
      RECT 17.070000  2.175000 17.600000 3.755000 ;
    LAYER mcon ;
      RECT  0.115000  0.425000  0.285000 0.595000 ;
      RECT  0.150000  3.475000  0.320000 3.645000 ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.475000  0.425000  0.645000 0.595000 ;
      RECT  0.510000  3.475000  0.680000 3.645000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.340000  0.425000  1.510000 0.595000 ;
      RECT  1.340000  3.475000  1.510000 3.645000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  1.700000  0.425000  1.870000 0.595000 ;
      RECT  1.700000  3.475000  1.870000 3.645000 ;
      RECT  2.060000  0.425000  2.230000 0.595000 ;
      RECT  2.060000  3.475000  2.230000 3.645000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.880000  3.475000  3.050000 3.645000 ;
      RECT  2.960000  0.425000  3.130000 0.595000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.240000  3.475000  3.410000 3.645000 ;
      RECT  3.320000  0.425000  3.490000 0.595000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.600000  3.475000  3.770000 3.645000 ;
      RECT  3.680000  0.425000  3.850000 0.595000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.440000  0.425000  4.610000 0.595000 ;
      RECT  4.460000  3.475000  4.630000 3.645000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.800000  0.425000  4.970000 0.595000 ;
      RECT  4.800000  1.580000  4.970000 1.750000 ;
      RECT  4.820000  3.475000  4.990000 3.645000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.160000  0.425000  5.330000 0.595000 ;
      RECT  5.160000  1.580000  5.330000 1.750000 ;
      RECT  5.180000  3.475000  5.350000 3.645000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.650000  2.320000  5.820000 2.490000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.070000  0.425000  6.240000 0.595000 ;
      RECT  6.070000  3.475000  6.240000 3.645000 ;
      RECT  6.230000  1.580000  6.400000 1.750000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.430000  0.425000  6.600000 0.595000 ;
      RECT  6.430000  3.475000  6.600000 3.645000 ;
      RECT  6.590000  1.580000  6.760000 1.750000 ;
      RECT  6.790000  0.425000  6.960000 0.595000 ;
      RECT  6.790000  3.475000  6.960000 3.645000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.210000  2.320000  7.380000 2.490000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.630000  0.425000  7.800000 0.595000 ;
      RECT  7.630000  3.475000  7.800000 3.645000 ;
      RECT  7.790000  1.580000  7.960000 1.750000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  7.990000  0.425000  8.160000 0.595000 ;
      RECT  7.990000  3.475000  8.160000 3.645000 ;
      RECT  8.150000  1.580000  8.320000 1.750000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.350000  0.425000  8.520000 0.595000 ;
      RECT  8.350000  3.475000  8.520000 3.645000 ;
      RECT  8.770000  2.320000  8.940000 2.490000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.190000  0.425000  9.360000 0.595000 ;
      RECT  9.190000  3.475000  9.360000 3.645000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.350000  1.580000  9.520000 1.750000 ;
      RECT  9.550000  0.425000  9.720000 0.595000 ;
      RECT  9.550000  3.475000  9.720000 3.645000 ;
      RECT  9.710000  1.580000  9.880000 1.750000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.910000  0.425000 10.080000 0.595000 ;
      RECT  9.910000  3.475000 10.080000 3.645000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.330000  2.320000 10.500000 2.490000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.750000  0.425000 10.920000 0.595000 ;
      RECT 10.750000  3.475000 10.920000 3.645000 ;
      RECT 10.910000  1.580000 11.080000 1.750000 ;
      RECT 11.110000  0.425000 11.280000 0.595000 ;
      RECT 11.110000  3.475000 11.280000 3.645000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.270000  1.580000 11.440000 1.750000 ;
      RECT 11.470000  0.425000 11.640000 0.595000 ;
      RECT 11.470000  3.475000 11.640000 3.645000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 11.890000  2.320000 12.060000 2.490000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.310000  0.425000 12.480000 0.595000 ;
      RECT 12.310000  3.475000 12.480000 3.645000 ;
      RECT 12.470000  1.580000 12.640000 1.750000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 12.670000  0.425000 12.840000 0.595000 ;
      RECT 12.670000  3.475000 12.840000 3.645000 ;
      RECT 12.830000  1.580000 13.000000 1.750000 ;
      RECT 13.030000  0.425000 13.200000 0.595000 ;
      RECT 13.030000  3.475000 13.200000 3.645000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.450000  2.320000 13.620000 2.490000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.870000  0.425000 14.040000 0.595000 ;
      RECT 13.870000  3.475000 14.040000 3.645000 ;
      RECT 14.030000  1.580000 14.200000 1.750000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.230000  0.425000 14.400000 0.595000 ;
      RECT 14.230000  3.475000 14.400000 3.645000 ;
      RECT 14.390000  1.580000 14.560000 1.750000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.590000  0.425000 14.760000 0.595000 ;
      RECT 14.590000  3.475000 14.760000 3.645000 ;
      RECT 15.010000  2.320000 15.180000 2.490000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.430000  0.425000 15.600000 0.595000 ;
      RECT 15.430000  3.475000 15.600000 3.645000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.590000  1.580000 15.760000 1.750000 ;
      RECT 15.790000  0.425000 15.960000 0.595000 ;
      RECT 15.790000  3.475000 15.960000 3.645000 ;
      RECT 15.950000  1.580000 16.120000 1.750000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.150000  0.425000 16.320000 0.595000 ;
      RECT 16.150000  3.475000 16.320000 3.645000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.570000  2.320000 16.740000 2.490000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 17.070000  0.425000 17.240000 0.595000 ;
      RECT 17.070000  3.475000 17.240000 3.645000 ;
      RECT 17.430000  0.425000 17.600000 0.595000 ;
      RECT 17.430000  3.475000 17.600000 3.645000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
    LAYER met1 ;
      RECT  4.740000 1.550000  5.360000 1.580000 ;
      RECT  4.740000 1.580000 16.250000 1.750000 ;
      RECT  4.740000 1.750000  5.360000 1.780000 ;
      RECT  6.170000 1.550000  6.820000 1.580000 ;
      RECT  6.170000 1.750000  6.820000 1.780000 ;
      RECT  7.730000 1.550000  8.380000 1.580000 ;
      RECT  7.730000 1.750000  8.380000 1.780000 ;
      RECT  9.290000 1.550000  9.940000 1.580000 ;
      RECT  9.290000 1.750000  9.940000 1.780000 ;
      RECT 10.850000 1.550000 11.500000 1.580000 ;
      RECT 10.850000 1.750000 11.500000 1.780000 ;
      RECT 12.410000 1.550000 13.060000 1.580000 ;
      RECT 12.410000 1.750000 13.060000 1.780000 ;
      RECT 13.970000 1.550000 14.620000 1.580000 ;
      RECT 13.970000 1.750000 14.620000 1.780000 ;
      RECT 15.530000 1.550000 16.180000 1.580000 ;
      RECT 15.530000 1.750000 16.180000 1.780000 ;
  END
END sky130_fd_sc_hvl__buf_16
