* File: sky130_fd_sc_hvl__sdfstp_1.pxi.spice
* Created: Wed Sep  2 09:10:18 2020
* 
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%VNB N_VNB_M1031_b VNB N_VNB_c_3_p
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%VNB
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%VPB N_VPB_M1012_b VPB N_VPB_c_124_p
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%VPB
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%SCE N_SCE_c_292_n N_SCE_M1012_g N_SCE_c_294_n
+ N_SCE_M1029_g N_SCE_M1039_g N_SCE_c_296_n N_SCE_c_285_n N_SCE_c_301_p SCE SCE
+ N_SCE_M1031_g N_SCE_c_288_n N_SCE_c_289_n N_SCE_c_290_n
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%SCE
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%A_30_107# N_A_30_107#_M1031_s
+ N_A_30_107#_M1012_s N_A_30_107#_c_357_n N_A_30_107#_M1017_g
+ N_A_30_107#_c_350_n N_A_30_107#_c_352_n N_A_30_107#_c_361_n
+ N_A_30_107#_c_353_n N_A_30_107#_c_362_n N_A_30_107#_c_377_n
+ N_A_30_107#_c_354_n N_A_30_107#_c_363_n N_A_30_107#_M1007_g
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%A_30_107#
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%D N_D_M1006_g N_D_M1030_g D N_D_c_425_n
+ N_D_c_436_n PM_SKY130_FD_SC_HVL__SDFSTP_1%D
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%SCD SCD SCD SCD N_SCD_M1001_g N_SCD_M1021_g
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%SCD
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%CLK N_CLK_M1028_g N_CLK_c_484_n N_CLK_M1008_g
+ N_CLK_c_488_n CLK CLK CLK N_CLK_c_486_n PM_SKY130_FD_SC_HVL__SDFSTP_1%CLK
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%A_935_107# N_A_935_107#_M1028_d
+ N_A_935_107#_M1008_d N_A_935_107#_c_542_n N_A_935_107#_M1037_g
+ N_A_935_107#_c_545_n N_A_935_107#_M1019_g N_A_935_107#_c_521_n
+ N_A_935_107#_M1036_g N_A_935_107#_M1026_g N_A_935_107#_c_522_n
+ N_A_935_107#_c_551_n N_A_935_107#_c_523_n N_A_935_107#_c_608_p
+ N_A_935_107#_c_613_p N_A_935_107#_c_524_n N_A_935_107#_c_526_n
+ N_A_935_107#_c_586_p N_A_935_107#_c_528_n N_A_935_107#_c_554_n
+ N_A_935_107#_c_557_n N_A_935_107#_c_600_p N_A_935_107#_c_560_n
+ N_A_935_107#_c_561_n N_A_935_107#_c_562_n N_A_935_107#_c_649_p
+ N_A_935_107#_c_563_n N_A_935_107#_c_564_n N_A_935_107#_c_654_p
+ N_A_935_107#_c_565_n N_A_935_107#_c_628_p N_A_935_107#_c_589_p
+ N_A_935_107#_c_566_n N_A_935_107#_c_529_n N_A_935_107#_c_591_p
+ N_A_935_107#_c_530_n N_A_935_107#_c_531_n N_A_935_107#_c_532_n
+ N_A_935_107#_c_534_n N_A_935_107#_c_535_n N_A_935_107#_c_536_n
+ N_A_935_107#_c_665_p N_A_935_107#_c_569_n N_A_935_107#_c_537_n
+ N_A_935_107#_M1002_g N_A_935_107#_M1034_g
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%A_935_107#
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%A_1201_123# N_A_1201_123#_M1002_d
+ N_A_1201_123#_M1037_d N_A_1201_123#_M1004_g N_A_1201_123#_M1024_g
+ N_A_1201_123#_M1013_g N_A_1201_123#_c_801_n N_A_1201_123#_M1005_g
+ N_A_1201_123#_c_792_n N_A_1201_123#_c_802_n N_A_1201_123#_c_793_n
+ N_A_1201_123#_c_794_n N_A_1201_123#_c_795_n N_A_1201_123#_c_796_n
+ N_A_1201_123#_c_797_n N_A_1201_123#_c_805_n N_A_1201_123#_c_806_n
+ N_A_1201_123#_c_807_n N_A_1201_123#_c_798_n N_A_1201_123#_c_799_n
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%A_1201_123#
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%A_1669_87# N_A_1669_87#_M1022_s
+ N_A_1669_87#_M1018_d N_A_1669_87#_c_948_n N_A_1669_87#_M1025_g
+ N_A_1669_87#_c_954_n N_A_1669_87#_c_949_n N_A_1669_87#_c_950_n
+ N_A_1669_87#_c_951_n N_A_1669_87#_c_965_n N_A_1669_87#_c_973_n
+ N_A_1669_87#_c_953_n N_A_1669_87#_M1000_g
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%A_1669_87#
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%A_1471_113# N_A_1471_113#_M1034_d
+ N_A_1471_113#_M1004_d N_A_1471_113#_M1022_g N_A_1471_113#_M1016_g
+ N_A_1471_113#_M1011_g N_A_1471_113#_c_1011_n N_A_1471_113#_c_1013_n
+ N_A_1471_113#_c_1014_n N_A_1471_113#_c_1026_n N_A_1471_113#_c_1027_n
+ N_A_1471_113#_c_1015_n N_A_1471_113#_c_1016_n N_A_1471_113#_c_1017_n
+ N_A_1471_113#_c_1018_n N_A_1471_113#_c_1050_n N_A_1471_113#_c_1029_n
+ N_A_1471_113#_c_1020_n N_A_1471_113#_c_1021_n N_A_1471_113#_c_1022_n
+ N_A_1471_113#_c_1110_n N_A_1471_113#_M1018_g
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%A_1471_113#
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%SET_B N_SET_B_M1027_g N_SET_B_c_1156_n
+ N_SET_B_c_1146_n N_SET_B_c_1165_n N_SET_B_c_1147_n N_SET_B_c_1149_n SET_B
+ SET_B SET_B N_SET_B_M1010_g N_SET_B_M1015_g N_SET_B_M1038_g N_SET_B_c_1155_n
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%SET_B
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%A_2698_421# N_A_2698_421#_M1023_d
+ N_A_2698_421#_M1020_s N_A_2698_421#_M1009_g N_A_2698_421#_M1014_g
+ N_A_2698_421#_c_1237_n N_A_2698_421#_c_1238_n N_A_2698_421#_c_1239_n
+ N_A_2698_421#_c_1240_n N_A_2698_421#_c_1243_n N_A_2698_421#_c_1246_n
+ N_A_2698_421#_c_1247_n N_A_2698_421#_c_1235_n N_A_2698_421#_c_1248_n
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%A_2698_421#
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%A_2477_543# N_A_2477_543#_M1013_d
+ N_A_2477_543#_M1019_d N_A_2477_543#_M1038_d N_A_2477_543#_M1023_g
+ N_A_2477_543#_M1020_g N_A_2477_543#_c_1307_n N_A_2477_543#_M1032_g
+ N_A_2477_543#_M1033_g N_A_2477_543#_c_1309_n N_A_2477_543#_c_1318_n
+ N_A_2477_543#_c_1332_n N_A_2477_543#_c_1310_n N_A_2477_543#_c_1322_n
+ N_A_2477_543#_c_1323_n N_A_2477_543#_c_1324_n N_A_2477_543#_c_1370_n
+ N_A_2477_543#_c_1325_n N_A_2477_543#_c_1350_n N_A_2477_543#_c_1326_n
+ N_A_2477_543#_c_1311_n PM_SKY130_FD_SC_HVL__SDFSTP_1%A_2477_543#
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%A_3321_173# N_A_3321_173#_M1032_s
+ N_A_3321_173#_M1033_s N_A_3321_173#_M1003_g N_A_3321_173#_M1035_g
+ N_A_3321_173#_c_1432_n N_A_3321_173#_c_1433_n N_A_3321_173#_c_1442_n
+ N_A_3321_173#_c_1438_n N_A_3321_173#_c_1439_n N_A_3321_173#_c_1459_n
+ N_A_3321_173#_c_1434_n PM_SKY130_FD_SC_HVL__SDFSTP_1%A_3321_173#
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%VPWR N_VPWR_M1012_d N_VPWR_M1021_d
+ N_VPWR_M1037_s N_VPWR_M1000_d N_VPWR_M1027_d N_VPWR_M1009_d N_VPWR_M1020_d
+ N_VPWR_M1033_d VPWR N_VPWR_c_1479_n N_VPWR_c_1482_n N_VPWR_c_1485_n
+ N_VPWR_c_1488_n N_VPWR_c_1491_n N_VPWR_c_1494_n N_VPWR_c_1497_n
+ N_VPWR_c_1500_n N_VPWR_c_1503_n PM_SKY130_FD_SC_HVL__SDFSTP_1%VPWR
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%A_481_107# N_A_481_107#_M1007_d
+ N_A_481_107#_M1034_s N_A_481_107#_M1030_d N_A_481_107#_M1004_s
+ N_A_481_107#_c_1610_n N_A_481_107#_c_1649_n N_A_481_107#_c_1611_n
+ N_A_481_107#_c_1617_n N_A_481_107#_c_1618_n N_A_481_107#_c_1673_n
+ N_A_481_107#_c_1619_n N_A_481_107#_c_1622_n N_A_481_107#_c_1625_n
+ N_A_481_107#_c_1626_n N_A_481_107#_c_1627_n N_A_481_107#_c_1628_n
+ N_A_481_107#_c_1629_n N_A_481_107#_c_1632_n N_A_481_107#_c_1635_n
+ N_A_481_107#_c_1636_n N_A_481_107#_c_1612_n N_A_481_107#_c_1637_n
+ N_A_481_107#_c_1661_n N_A_481_107#_c_1614_n N_A_481_107#_c_1615_n
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%A_481_107#
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%Q N_Q_M1003_d N_Q_M1035_d Q Q Q Q Q Q Q
+ N_Q_c_1748_n PM_SKY130_FD_SC_HVL__SDFSTP_1%Q
x_PM_SKY130_FD_SC_HVL__SDFSTP_1%VGND N_VGND_M1031_d N_VGND_M1001_d
+ N_VGND_M1002_s N_VGND_M1025_d N_VGND_M1010_d N_VGND_M1015_d N_VGND_M1032_d
+ VGND N_VGND_c_1760_n N_VGND_c_1762_n N_VGND_c_1764_n N_VGND_c_1766_n
+ N_VGND_c_1768_n N_VGND_c_1770_n N_VGND_c_1772_n N_VGND_c_1774_n
+ PM_SKY130_FD_SC_HVL__SDFSTP_1%VGND
cc_1 N_VNB_M1031_b N_SCE_c_285_n 0.0325683f $X=-0.33 $Y=-0.265 $X2=2.525
+ $Y2=1.58
cc_2 N_VNB_M1031_b N_SCE_M1031_g 0.125326f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=0.745
cc_3 N_VNB_c_3_p N_SCE_M1031_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=0.745
cc_4 N_VNB_M1031_b N_SCE_c_288_n 0.0726615f $X=-0.33 $Y=-0.265 $X2=2.8 $Y2=1.26
cc_5 N_VNB_M1031_b N_SCE_c_289_n 0.00493464f $X=-0.33 $Y=-0.265 $X2=2.8 $Y2=1.26
cc_6 N_VNB_M1031_b N_SCE_c_290_n 0.045087f $X=-0.33 $Y=-0.265 $X2=2.9 $Y2=1.075
cc_7 N_VNB_c_3_p N_SCE_c_290_n 0.0023273f $X=0.24 $Y=0 $X2=2.9 $Y2=1.075
cc_8 N_VNB_M1031_b N_A_30_107#_c_350_n 0.0310029f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_c_3_p N_A_30_107#_c_350_n 7.98897e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_10 N_VNB_M1031_b N_A_30_107#_c_352_n 0.0270621f $X=-0.33 $Y=-0.265 $X2=0.895
+ $Y2=1.58
cc_11 N_VNB_M1031_b N_A_30_107#_c_353_n 0.00980012f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1031_b N_A_30_107#_c_354_n 0.0154754f $X=-0.33 $Y=-0.265 $X2=2.707
+ $Y2=1.495
cc_13 N_VNB_M1031_b N_A_30_107#_M1007_g 0.0899623f $X=-0.33 $Y=-0.265 $X2=2.707
+ $Y2=1.295
cc_14 N_VNB_c_3_p N_A_30_107#_M1007_g 0.0023273f $X=0.24 $Y=0 $X2=2.707
+ $Y2=1.295
cc_15 N_VNB_M1031_b N_D_M1006_g 0.0937362f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=3.055
cc_16 N_VNB_c_3_p N_D_M1006_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=3.055
cc_17 N_VNB_M1031_b N_D_c_425_n 0.050044f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_18 N_VNB_M1031_b N_SCD_M1001_g 0.111002f $X=-0.33 $Y=-0.265 $X2=2.935
+ $Y2=0.745
cc_19 N_VNB_M1031_b N_CLK_M1028_g 0.0490406f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=3.055
cc_20 N_VNB_c_3_p N_CLK_M1028_g 0.00142431f $X=0.24 $Y=0 $X2=0.665 $Y2=3.055
cc_21 N_VNB_M1031_b N_CLK_c_484_n 0.0538882f $X=-0.33 $Y=-0.265 $X2=1.445
+ $Y2=3.055
cc_22 N_VNB_M1031_b CLK 0.00716946f $X=-0.33 $Y=-0.265 $X2=0.665 $Y2=2.235
cc_23 N_VNB_M1031_b N_CLK_c_486_n 0.0371453f $X=-0.33 $Y=-0.265 $X2=0.73
+ $Y2=1.66
cc_24 N_VNB_M1031_b N_A_935_107#_c_521_n 0.0776063f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_25 N_VNB_M1031_b N_A_935_107#_c_522_n 0.0175156f $X=-0.33 $Y=-0.265 $X2=2.9
+ $Y2=1.26
cc_26 N_VNB_M1031_b N_A_935_107#_c_523_n 0.0184674f $X=-0.33 $Y=-0.265 $X2=2.707
+ $Y2=1.495
cc_27 N_VNB_M1031_b N_A_935_107#_c_524_n 0.117892f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_28 N_VNB_c_3_p N_A_935_107#_c_524_n 0.00481902f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_29 N_VNB_M1031_b N_A_935_107#_c_526_n 0.0139086f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_30 N_VNB_c_3_p N_A_935_107#_c_526_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_31 N_VNB_M1031_b N_A_935_107#_c_528_n 0.00205295f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_32 N_VNB_M1031_b N_A_935_107#_c_529_n 0.00843232f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_33 N_VNB_M1031_b N_A_935_107#_c_530_n 0.00237288f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_M1031_b N_A_935_107#_c_531_n 0.00193739f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_35 N_VNB_M1031_b N_A_935_107#_c_532_n 0.019647f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_36 N_VNB_c_3_p N_A_935_107#_c_532_n 8.76825e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_37 N_VNB_M1031_b N_A_935_107#_c_534_n 0.00204459f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_38 N_VNB_M1031_b N_A_935_107#_c_535_n 8.03629e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_39 N_VNB_M1031_b N_A_935_107#_c_536_n 0.00363204f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_M1031_b N_A_935_107#_c_537_n 0.00224269f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_41 N_VNB_M1031_b N_A_935_107#_M1002_g 0.123567f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_42 N_VNB_c_3_p N_A_935_107#_M1002_g 5.37636e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_43 N_VNB_M1031_b N_A_935_107#_M1034_g 0.11061f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_44 N_VNB_c_3_p N_A_935_107#_M1034_g 5.61877e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_45 N_VNB_M1031_b N_A_1201_123#_M1024_g 0.0474885f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_c_3_p N_A_1201_123#_M1024_g 0.00224751f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_47 N_VNB_M1031_b N_A_1201_123#_M1013_g 0.0755963f $X=-0.33 $Y=-0.265 $X2=0.73
+ $Y2=1.58
cc_48 N_VNB_M1031_b N_A_1201_123#_c_792_n 0.00192959f $X=-0.33 $Y=-0.265
+ $X2=0.665 $Y2=0.745
cc_49 N_VNB_M1031_b N_A_1201_123#_c_793_n 0.0188958f $X=-0.33 $Y=-0.265 $X2=2.8
+ $Y2=1.26
cc_50 N_VNB_M1031_b N_A_1201_123#_c_794_n 0.00926345f $X=-0.33 $Y=-0.265
+ $X2=2.707 $Y2=1.495
cc_51 N_VNB_M1031_b N_A_1201_123#_c_795_n 0.00142625f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_52 N_VNB_M1031_b N_A_1201_123#_c_796_n 0.0544134f $X=-0.33 $Y=-0.265
+ $X2=2.707 $Y2=1.58
cc_53 N_VNB_M1031_b N_A_1201_123#_c_797_n 0.00696849f $X=-0.33 $Y=-0.265
+ $X2=2.707 $Y2=1.665
cc_54 N_VNB_M1031_b N_A_1201_123#_c_798_n 0.0190019f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_55 N_VNB_M1031_b N_A_1201_123#_c_799_n 0.0866134f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_56 N_VNB_M1031_b N_A_1669_87#_c_948_n 0.0395705f $X=-0.33 $Y=-0.265 $X2=2.935
+ $Y2=1.075
cc_57 N_VNB_M1031_b N_A_1669_87#_c_949_n 0.0268254f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_58 N_VNB_M1031_b N_A_1669_87#_c_950_n 0.00620141f $X=-0.33 $Y=-0.265
+ $X2=2.525 $Y2=1.58
cc_59 N_VNB_M1031_b N_A_1669_87#_c_951_n 0.0167518f $X=-0.33 $Y=-0.265 $X2=0.73
+ $Y2=1.66
cc_60 N_VNB_c_3_p N_A_1669_87#_c_951_n 7.98897e-19 $X=0.24 $Y=0 $X2=0.73
+ $Y2=1.66
cc_61 N_VNB_M1031_b N_A_1669_87#_c_953_n 0.0758152f $X=-0.33 $Y=-0.265 $X2=2.8
+ $Y2=1.26
cc_62 N_VNB_M1031_b N_A_1471_113#_M1011_g 0.0428346f $X=-0.33 $Y=-0.265
+ $X2=0.895 $Y2=1.58
cc_63 N_VNB_c_3_p N_A_1471_113#_M1011_g 8.58675e-19 $X=0.24 $Y=0 $X2=0.895
+ $Y2=1.58
cc_64 N_VNB_M1031_b N_A_1471_113#_c_1011_n 0.0516089f $X=-0.33 $Y=-0.265
+ $X2=0.73 $Y2=1.66
cc_65 N_VNB_c_3_p N_A_1471_113#_c_1011_n 0.0023273f $X=0.24 $Y=0 $X2=0.73
+ $Y2=1.66
cc_66 N_VNB_M1031_b N_A_1471_113#_c_1013_n 0.0633132f $X=-0.33 $Y=-0.265
+ $X2=2.555 $Y2=1.21
cc_67 N_VNB_M1031_b N_A_1471_113#_c_1014_n 7.89534e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_68 N_VNB_M1031_b N_A_1471_113#_c_1015_n 0.00727167f $X=-0.33 $Y=-0.265
+ $X2=2.8 $Y2=1.26
cc_69 N_VNB_M1031_b N_A_1471_113#_c_1016_n 0.0150463f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_70 N_VNB_M1031_b N_A_1471_113#_c_1017_n 0.0475753f $X=-0.33 $Y=-0.265
+ $X2=2.707 $Y2=1.295
cc_71 N_VNB_M1031_b N_A_1471_113#_c_1018_n 0.0173789f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_72 N_VNB_c_3_p N_A_1471_113#_c_1018_n 0.00118777f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_73 N_VNB_M1031_b N_A_1471_113#_c_1020_n 0.00348125f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_74 N_VNB_M1031_b N_A_1471_113#_c_1021_n 0.0299364f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_75 N_VNB_M1031_b N_A_1471_113#_c_1022_n 0.00670334f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_76 N_VNB_M1031_b N_SET_B_c_1146_n 0.00421789f $X=-0.33 $Y=-0.265 $X2=2.935
+ $Y2=1.075
cc_77 N_VNB_M1031_b N_SET_B_c_1147_n 0.205517f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_78 N_VNB_c_3_p N_SET_B_c_1147_n 0.00870408f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_79 N_VNB_M1031_b N_SET_B_c_1149_n 0.0135491f $X=-0.33 $Y=-0.265 $X2=2.525
+ $Y2=1.58
cc_80 N_VNB_c_3_p N_SET_B_c_1149_n 5.63772e-19 $X=0.24 $Y=0 $X2=2.525 $Y2=1.58
cc_81 N_VNB_M1031_b SET_B 7.27841e-19 $X=-0.33 $Y=-0.265 $X2=0.73 $Y2=1.66
cc_82 N_VNB_M1031_b SET_B 0.00201087f $X=-0.33 $Y=-0.265 $X2=0.73 $Y2=1.66
cc_83 N_VNB_M1031_b N_SET_B_M1010_g 0.110528f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=0.745
cc_84 N_VNB_M1031_b N_SET_B_M1015_g 0.0916883f $X=-0.33 $Y=-0.265 $X2=2.8
+ $Y2=1.26
cc_85 N_VNB_M1031_b N_SET_B_c_1155_n 0.0105949f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_86 N_VNB_M1031_b N_A_2698_421#_M1014_g 0.0738661f $X=-0.33 $Y=-0.265
+ $X2=1.445 $Y2=2.485
cc_87 N_VNB_M1031_b N_A_2698_421#_c_1235_n 0.0144478f $X=-0.33 $Y=-0.265 $X2=2.8
+ $Y2=1.26
cc_88 N_VNB_M1031_b N_A_2477_543#_M1023_g 0.0468003f $X=-0.33 $Y=-0.265
+ $X2=1.445 $Y2=2.485
cc_89 N_VNB_M1031_b N_A_2477_543#_c_1307_n 0.0714245f $X=-0.33 $Y=-0.265
+ $X2=0.73 $Y2=1.66
cc_90 N_VNB_M1031_b N_A_2477_543#_M1032_g 0.0492136f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_91 N_VNB_M1031_b N_A_2477_543#_c_1309_n 0.0365535f $X=-0.33 $Y=-0.265 $X2=2.9
+ $Y2=1.26
cc_92 N_VNB_M1031_b N_A_2477_543#_c_1310_n 0.00566183f $X=-0.33 $Y=-0.265
+ $X2=2.707 $Y2=1.58
cc_93 N_VNB_M1031_b N_A_2477_543#_c_1311_n 0.0669545f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_94 N_VNB_M1031_b N_A_3321_173#_M1003_g 0.0502601f $X=-0.33 $Y=-0.265
+ $X2=2.935 $Y2=0.745
cc_95 N_VNB_c_3_p N_A_3321_173#_M1003_g 0.00112176f $X=0.24 $Y=0 $X2=2.935
+ $Y2=0.745
cc_96 N_VNB_M1031_b N_A_3321_173#_c_1432_n 0.013755f $X=-0.33 $Y=-0.265 $X2=0.73
+ $Y2=1.58
cc_97 N_VNB_M1031_b N_A_3321_173#_c_1433_n 0.0131103f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_98 N_VNB_M1031_b N_A_3321_173#_c_1434_n 0.0526842f $X=-0.33 $Y=-0.265
+ $X2=2.707 $Y2=1.495
cc_99 N_VNB_M1031_b N_A_481_107#_c_1610_n 0.00506017f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_100 N_VNB_M1031_b N_A_481_107#_c_1611_n 0.00773422f $X=-0.33 $Y=-0.265
+ $X2=0.73 $Y2=1.66
cc_101 N_VNB_M1031_b N_A_481_107#_c_1612_n 0.0109104f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_102 N_VNB_c_3_p N_A_481_107#_c_1612_n 8.65969e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_103 N_VNB_M1031_b N_A_481_107#_c_1614_n 0.00796369f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_104 N_VNB_M1031_b N_A_481_107#_c_1615_n 0.00896739f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_105 N_VNB_M1031_b N_Q_c_1748_n 0.0649641f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_106 N_VNB_c_3_p N_Q_c_1748_n 8.66888e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_107 N_VNB_M1031_b N_VGND_c_1760_n 0.0468651f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=0.745
cc_108 N_VNB_c_3_p N_VGND_c_1760_n 0.00269953f $X=0.24 $Y=0 $X2=0.665 $Y2=0.745
cc_109 N_VNB_M1031_b N_VGND_c_1762_n 0.0518185f $X=-0.33 $Y=-0.265 $X2=2.707
+ $Y2=1.26
cc_110 N_VNB_c_3_p N_VGND_c_1762_n 0.00269373f $X=0.24 $Y=0 $X2=2.707 $Y2=1.26
cc_111 N_VNB_M1031_b N_VGND_c_1764_n 0.0317956f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_112 N_VNB_c_3_p N_VGND_c_1764_n 7.0368e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_113 N_VNB_M1031_b N_VGND_c_1766_n 0.0546544f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_114 N_VNB_c_3_p N_VGND_c_1766_n 0.00270051f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_115 N_VNB_M1031_b N_VGND_c_1768_n 0.0504695f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_116 N_VNB_c_3_p N_VGND_c_1768_n 0.00269373f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_117 N_VNB_M1031_b N_VGND_c_1770_n 0.069283f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_118 N_VNB_c_3_p N_VGND_c_1770_n 0.00252021f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_119 N_VNB_M1031_b N_VGND_c_1772_n 0.0613398f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_120 N_VNB_c_3_p N_VGND_c_1772_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_121 N_VNB_M1031_b N_VGND_c_1774_n 0.29611f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_122 N_VNB_c_3_p N_VGND_c_1774_n 2.00125f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_123 N_VPB_M1012_b N_SCE_c_292_n 0.0413919f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=2.735
cc_124 N_VPB_c_124_p N_SCE_c_292_n 0.00540119f $X=18.48 $Y=4.07 $X2=0.665
+ $Y2=2.735
cc_125 N_VPB_M1012_b N_SCE_c_294_n 0.0354165f $X=-0.33 $Y=1.885 $X2=1.445
+ $Y2=2.735
cc_126 N_VPB_c_124_p N_SCE_c_294_n 0.00386003f $X=18.48 $Y=4.07 $X2=1.445
+ $Y2=2.735
cc_127 N_VPB_M1012_b N_SCE_c_296_n 0.11064f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=2.485
cc_128 N_VPB_M1012_b N_SCE_M1031_g 0.0420682f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=0.745
cc_129 N_VPB_M1012_b N_A_30_107#_c_357_n 0.0722858f $X=-0.33 $Y=1.885 $X2=2.935
+ $Y2=1.075
cc_130 N_VPB_M1012_b N_A_30_107#_M1017_g 0.0396839f $X=-0.33 $Y=1.885 $X2=2.935
+ $Y2=0.745
cc_131 N_VPB_c_124_p N_A_30_107#_M1017_g 0.0110649f $X=18.48 $Y=4.07 $X2=2.935
+ $Y2=0.745
cc_132 N_VPB_M1012_b N_A_30_107#_c_352_n 0.0313207f $X=-0.33 $Y=1.885 $X2=0.895
+ $Y2=1.58
cc_133 N_VPB_M1012_b N_A_30_107#_c_361_n 0.0268401f $X=-0.33 $Y=1.885 $X2=0.73
+ $Y2=1.66
cc_134 N_VPB_M1012_b N_A_30_107#_c_362_n 0.0189891f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_135 N_VPB_M1012_b N_A_30_107#_c_363_n 0.0132078f $X=-0.33 $Y=1.885 $X2=2.707
+ $Y2=1.26
cc_136 N_VPB_M1012_b N_D_M1030_g 0.100451f $X=-0.33 $Y=1.885 $X2=2.935 $Y2=1.075
cc_137 N_VPB_c_124_p N_D_M1030_g 0.0110649f $X=18.48 $Y=4.07 $X2=2.935 $Y2=1.075
cc_138 N_VPB_M1012_b N_D_c_425_n 0.0487498f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_139 N_VPB_M1012_b N_SCD_M1001_g 0.111112f $X=-0.33 $Y=1.885 $X2=2.935
+ $Y2=0.745
cc_140 N_VPB_c_124_p N_SCD_M1001_g 0.00193359f $X=18.48 $Y=4.07 $X2=2.935
+ $Y2=0.745
cc_141 N_VPB_M1012_b N_CLK_c_484_n 0.061208f $X=-0.33 $Y=1.885 $X2=1.445
+ $Y2=3.055
cc_142 N_VPB_M1012_b N_CLK_c_488_n 0.0769451f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=2.485
cc_143 VPB N_CLK_c_488_n 0.00104305f $X=0 $Y=3.955 $X2=0.665 $Y2=2.485
cc_144 N_VPB_c_124_p N_CLK_c_488_n 0.00653579f $X=18.48 $Y=4.07 $X2=0.665
+ $Y2=2.485
cc_145 N_VPB_M1012_b CLK 0.00443942f $X=-0.33 $Y=1.885 $X2=0.665 $Y2=2.235
cc_146 N_VPB_M1012_b N_A_935_107#_c_542_n 0.081629f $X=-0.33 $Y=1.885 $X2=2.935
+ $Y2=1.075
cc_147 VPB N_A_935_107#_c_542_n 5.14587e-19 $X=0 $Y=3.955 $X2=2.935 $Y2=1.075
cc_148 N_VPB_c_124_p N_A_935_107#_c_542_n 0.00310579f $X=18.48 $Y=4.07 $X2=2.935
+ $Y2=1.075
cc_149 N_VPB_M1012_b N_A_935_107#_c_545_n 0.0352336f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=2.485
cc_150 N_VPB_M1012_b N_A_935_107#_M1019_g 0.0394981f $X=-0.33 $Y=1.885 $X2=1.445
+ $Y2=2.485
cc_151 VPB N_A_935_107#_M1019_g 0.00970178f $X=0 $Y=3.955 $X2=1.445 $Y2=2.485
cc_152 N_VPB_c_124_p N_A_935_107#_M1019_g 0.0193887f $X=18.48 $Y=4.07 $X2=1.445
+ $Y2=2.485
cc_153 N_VPB_M1012_b N_A_935_107#_c_521_n 0.00717334f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_154 N_VPB_M1012_b N_A_935_107#_M1026_g 0.0411776f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=0.745
cc_155 N_VPB_M1012_b N_A_935_107#_c_551_n 0.0220628f $X=-0.33 $Y=1.885 $X2=2.9
+ $Y2=1.075
cc_156 N_VPB_M1012_b N_A_935_107#_c_523_n 0.0102397f $X=-0.33 $Y=1.885 $X2=2.707
+ $Y2=1.495
cc_157 N_VPB_M1012_b N_A_935_107#_c_528_n 0.0055263f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_158 N_VPB_M1012_b N_A_935_107#_c_554_n 0.0174324f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_159 VPB N_A_935_107#_c_554_n 0.00191626f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_160 N_VPB_c_124_p N_A_935_107#_c_554_n 0.0203558f $X=18.48 $Y=4.07 $X2=0
+ $Y2=0
cc_161 N_VPB_M1012_b N_A_935_107#_c_557_n 0.002919f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_162 VPB N_A_935_107#_c_557_n 3.71311e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_163 N_VPB_c_124_p N_A_935_107#_c_557_n 0.00411424f $X=18.48 $Y=4.07 $X2=0
+ $Y2=0
cc_164 N_VPB_M1012_b N_A_935_107#_c_560_n 0.0348582f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_165 N_VPB_M1012_b N_A_935_107#_c_561_n 0.0039068f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_166 N_VPB_M1012_b N_A_935_107#_c_562_n 0.00650467f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_167 N_VPB_M1012_b N_A_935_107#_c_563_n 0.00760745f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_168 N_VPB_M1012_b N_A_935_107#_c_564_n 0.00232023f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_169 N_VPB_M1012_b N_A_935_107#_c_565_n 0.00195104f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_170 N_VPB_M1012_b N_A_935_107#_c_566_n 0.00454934f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_171 N_VPB_M1012_b N_A_935_107#_c_530_n 0.00711877f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_172 N_VPB_M1012_b N_A_935_107#_c_534_n 2.72612e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_173 N_VPB_M1012_b N_A_935_107#_c_569_n 0.00216962f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_174 N_VPB_M1012_b N_A_935_107#_M1002_g 0.0512353f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_175 N_VPB_M1012_b N_A_1201_123#_M1004_g 0.0390771f $X=-0.33 $Y=1.885
+ $X2=2.935 $Y2=0.745
cc_176 N_VPB_M1012_b N_A_1201_123#_c_801_n 0.0398688f $X=-0.33 $Y=1.885 $X2=0.73
+ $Y2=1.66
cc_177 N_VPB_M1012_b N_A_1201_123#_c_802_n 0.00372622f $X=-0.33 $Y=1.885 $X2=2.9
+ $Y2=1.26
cc_178 N_VPB_M1012_b N_A_1201_123#_c_793_n 0.0288896f $X=-0.33 $Y=1.885 $X2=2.8
+ $Y2=1.26
cc_179 N_VPB_M1012_b N_A_1201_123#_c_796_n 0.00786525f $X=-0.33 $Y=1.885
+ $X2=2.707 $Y2=1.58
cc_180 N_VPB_M1012_b N_A_1201_123#_c_805_n 0.00293847f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_181 N_VPB_M1012_b N_A_1201_123#_c_806_n 0.00348554f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_182 N_VPB_M1012_b N_A_1201_123#_c_807_n 0.0017887f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_183 N_VPB_M1012_b N_A_1201_123#_c_798_n 0.103499f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_184 N_VPB_M1012_b N_A_1201_123#_c_799_n 0.188649f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_185 N_VPB_M1012_b N_A_1669_87#_c_954_n 0.00907499f $X=-0.33 $Y=1.885
+ $X2=0.665 $Y2=2.485
cc_186 N_VPB_M1012_b N_A_1669_87#_c_949_n 0.103733f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_187 N_VPB_M1012_b N_A_1471_113#_M1016_g 0.104272f $X=-0.33 $Y=1.885 $X2=1.445
+ $Y2=2.485
cc_188 VPB N_A_1471_113#_M1016_g 0.00970178f $X=0 $Y=3.955 $X2=1.445 $Y2=2.485
cc_189 N_VPB_c_124_p N_A_1471_113#_M1016_g 0.013715f $X=18.48 $Y=4.07 $X2=1.445
+ $Y2=2.485
cc_190 N_VPB_M1012_b N_A_1471_113#_c_1026_n 0.00193084f $X=-0.33 $Y=1.885
+ $X2=0.665 $Y2=0.745
cc_191 N_VPB_M1012_b N_A_1471_113#_c_1027_n 0.00227208f $X=-0.33 $Y=1.885
+ $X2=0.665 $Y2=1.66
cc_192 N_VPB_M1012_b N_A_1471_113#_c_1017_n 0.00500453f $X=-0.33 $Y=1.885
+ $X2=2.707 $Y2=1.295
cc_193 N_VPB_M1012_b N_A_1471_113#_c_1029_n 0.00236711f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_194 N_VPB_M1012_b N_A_1471_113#_c_1021_n 0.0999848f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_195 N_VPB_M1012_b N_SET_B_c_1156_n 0.0925428f $X=-0.33 $Y=1.885 $X2=1.445
+ $Y2=3.055
cc_196 N_VPB_M1012_b N_SET_B_M1010_g 0.0191578f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=0.745
cc_197 N_VPB_M1012_b N_SET_B_M1015_g 0.105251f $X=-0.33 $Y=1.885 $X2=2.8
+ $Y2=1.26
cc_198 N_VPB_M1012_b N_A_2698_421#_M1014_g 0.020625f $X=-0.33 $Y=1.885 $X2=1.445
+ $Y2=2.485
cc_199 N_VPB_M1012_b N_A_2698_421#_c_1237_n 0.00538603f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_200 N_VPB_M1012_b N_A_2698_421#_c_1238_n 0.0493852f $X=-0.33 $Y=1.885
+ $X2=0.73 $Y2=1.58
cc_201 N_VPB_M1012_b N_A_2698_421#_c_1239_n 0.00301661f $X=-0.33 $Y=1.885
+ $X2=2.555 $Y2=1.21
cc_202 N_VPB_M1012_b N_A_2698_421#_c_1240_n 0.024262f $X=-0.33 $Y=1.885
+ $X2=2.555 $Y2=1.58
cc_203 VPB N_A_2698_421#_c_1240_n 0.00234622f $X=0 $Y=3.955 $X2=2.555 $Y2=1.58
cc_204 N_VPB_c_124_p N_A_2698_421#_c_1240_n 0.0236375f $X=18.48 $Y=4.07
+ $X2=2.555 $Y2=1.58
cc_205 N_VPB_M1012_b N_A_2698_421#_c_1243_n 0.00296331f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_206 VPB N_A_2698_421#_c_1243_n 3.61175e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_207 N_VPB_c_124_p N_A_2698_421#_c_1243_n 0.00388086f $X=18.48 $Y=4.07 $X2=0
+ $Y2=0
cc_208 N_VPB_M1012_b N_A_2698_421#_c_1246_n 0.00850178f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_209 N_VPB_M1012_b N_A_2698_421#_c_1247_n 0.00631733f $X=-0.33 $Y=1.885
+ $X2=0.665 $Y2=1.66
cc_210 N_VPB_M1012_b N_A_2698_421#_c_1248_n 0.0333105f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_211 N_VPB_M1012_b N_A_2477_543#_M1020_g 0.130455f $X=-0.33 $Y=1.885 $X2=0.895
+ $Y2=1.58
cc_212 VPB N_A_2477_543#_M1020_g 9.49031e-19 $X=0 $Y=3.955 $X2=0.895 $Y2=1.58
cc_213 N_VPB_c_124_p N_A_2477_543#_M1020_g 0.00564585f $X=18.48 $Y=4.07
+ $X2=0.895 $Y2=1.58
cc_214 N_VPB_M1012_b N_A_2477_543#_c_1307_n 0.0308499f $X=-0.33 $Y=1.885
+ $X2=0.73 $Y2=1.66
cc_215 N_VPB_M1012_b N_A_2477_543#_M1033_g 0.0746129f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_216 N_VPB_M1012_b N_A_2477_543#_c_1309_n 0.0023398f $X=-0.33 $Y=1.885 $X2=2.9
+ $Y2=1.26
cc_217 N_VPB_M1012_b N_A_2477_543#_c_1318_n 0.00886411f $X=-0.33 $Y=1.885
+ $X2=2.9 $Y2=1.075
cc_218 VPB N_A_2477_543#_c_1318_n 0.00104693f $X=0 $Y=3.955 $X2=2.9 $Y2=1.075
cc_219 N_VPB_c_124_p N_A_2477_543#_c_1318_n 0.0172373f $X=18.48 $Y=4.07 $X2=2.9
+ $Y2=1.075
cc_220 N_VPB_M1012_b N_A_2477_543#_c_1310_n 7.27999e-19 $X=-0.33 $Y=1.885
+ $X2=2.707 $Y2=1.58
cc_221 N_VPB_M1012_b N_A_2477_543#_c_1322_n 8.1348e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_222 N_VPB_M1012_b N_A_2477_543#_c_1323_n 0.0172685f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_223 N_VPB_M1012_b N_A_2477_543#_c_1324_n 0.0138448f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_224 N_VPB_M1012_b N_A_2477_543#_c_1325_n 0.00345197f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_225 N_VPB_M1012_b N_A_2477_543#_c_1326_n 0.0176571f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_226 N_VPB_M1012_b N_A_2477_543#_c_1311_n 0.0591383f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_227 N_VPB_M1012_b N_A_3321_173#_M1035_g 0.0446362f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_228 VPB N_A_3321_173#_M1035_g 8.8035e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_229 N_VPB_c_124_p N_A_3321_173#_M1035_g 0.00465039f $X=18.48 $Y=4.07 $X2=0
+ $Y2=0
cc_230 N_VPB_M1012_b N_A_3321_173#_c_1438_n 0.0172285f $X=-0.33 $Y=1.885 $X2=2.8
+ $Y2=1.26
cc_231 N_VPB_M1012_b N_A_3321_173#_c_1439_n 0.0113325f $X=-0.33 $Y=1.885 $X2=2.8
+ $Y2=1.26
cc_232 N_VPB_M1012_b N_A_3321_173#_c_1434_n 0.0416092f $X=-0.33 $Y=1.885
+ $X2=2.707 $Y2=1.495
cc_233 N_VPB_M1012_b N_VPWR_c_1479_n 0.0203426f $X=-0.33 $Y=1.885 $X2=2.9
+ $Y2=1.26
cc_234 VPB N_VPWR_c_1479_n 0.00269049f $X=0 $Y=3.955 $X2=2.9 $Y2=1.26
cc_235 N_VPB_c_124_p N_VPWR_c_1479_n 0.0409968f $X=18.48 $Y=4.07 $X2=2.9
+ $Y2=1.26
cc_236 N_VPB_M1012_b N_VPWR_c_1482_n 0.0166293f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1482_n 0.00258014f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_238 N_VPB_c_124_p N_VPWR_c_1482_n 0.0385227f $X=18.48 $Y=4.07 $X2=0 $Y2=0
cc_239 N_VPB_M1012_b N_VPWR_c_1485_n 0.00710721f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1485_n 5.05177e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_241 N_VPB_c_124_p N_VPWR_c_1485_n 0.00769771f $X=18.48 $Y=4.07 $X2=0 $Y2=0
cc_242 N_VPB_M1012_b N_VPWR_c_1488_n 0.0318697f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1488_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_244 N_VPB_c_124_p N_VPWR_c_1488_n 0.0409968f $X=18.48 $Y=4.07 $X2=0 $Y2=0
cc_245 N_VPB_M1012_b N_VPWR_c_1491_n 0.0143787f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1491_n 0.00370794f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_247 N_VPB_c_124_p N_VPWR_c_1491_n 0.0478243f $X=18.48 $Y=4.07 $X2=0 $Y2=0
cc_248 N_VPB_M1012_b N_VPWR_c_1494_n 0.0305748f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1494_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_250 N_VPB_c_124_p N_VPWR_c_1494_n 0.0409968f $X=18.48 $Y=4.07 $X2=0 $Y2=0
cc_251 N_VPB_M1012_b N_VPWR_c_1497_n 0.0316946f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1497_n 0.00166957f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_253 N_VPB_c_124_p N_VPWR_c_1497_n 0.025416f $X=18.48 $Y=4.07 $X2=0 $Y2=0
cc_254 N_VPB_M1012_b N_VPWR_c_1500_n 0.0366882f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1500_n 0.0026763f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_256 N_VPB_c_124_p N_VPWR_c_1500_n 0.0407806f $X=18.48 $Y=4.07 $X2=0 $Y2=0
cc_257 N_VPB_M1012_b N_VPWR_c_1503_n 0.265206f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1503_n 2.00034f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_259 N_VPB_c_124_p N_VPWR_c_1503_n 0.0994181f $X=18.48 $Y=4.07 $X2=0 $Y2=0
cc_260 N_VPB_M1012_b N_A_481_107#_c_1611_n 0.00612158f $X=-0.33 $Y=1.885
+ $X2=0.73 $Y2=1.66
cc_261 N_VPB_M1012_b N_A_481_107#_c_1617_n 0.00193804f $X=-0.33 $Y=1.885
+ $X2=2.555 $Y2=1.21
cc_262 N_VPB_M1012_b N_A_481_107#_c_1618_n 0.0180378f $X=-0.33 $Y=1.885
+ $X2=2.555 $Y2=1.58
cc_263 N_VPB_M1012_b N_A_481_107#_c_1619_n 0.00964404f $X=-0.33 $Y=1.885
+ $X2=0.665 $Y2=0.745
cc_264 VPB N_A_481_107#_c_1619_n 0.00235993f $X=0 $Y=3.955 $X2=0.665 $Y2=0.745
cc_265 N_VPB_c_124_p N_A_481_107#_c_1619_n 0.0462904f $X=18.48 $Y=4.07 $X2=0.665
+ $Y2=0.745
cc_266 N_VPB_M1012_b N_A_481_107#_c_1622_n 0.00164055f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_267 VPB N_A_481_107#_c_1622_n 5.70856e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_268 N_VPB_c_124_p N_A_481_107#_c_1622_n 0.0114989f $X=18.48 $Y=4.07 $X2=0
+ $Y2=0
cc_269 N_VPB_M1012_b N_A_481_107#_c_1625_n 0.0234622f $X=-0.33 $Y=1.885 $X2=2.9
+ $Y2=1.26
cc_270 N_VPB_M1012_b N_A_481_107#_c_1626_n 0.0101542f $X=-0.33 $Y=1.885 $X2=2.8
+ $Y2=1.26
cc_271 N_VPB_M1012_b N_A_481_107#_c_1627_n 0.00421263f $X=-0.33 $Y=1.885 $X2=2.8
+ $Y2=1.26
cc_272 N_VPB_M1012_b N_A_481_107#_c_1628_n 0.00112416f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_273 N_VPB_M1012_b N_A_481_107#_c_1629_n 0.0172109f $X=-0.33 $Y=1.885
+ $X2=2.707 $Y2=1.495
cc_274 VPB N_A_481_107#_c_1629_n 0.00342347f $X=0 $Y=3.955 $X2=2.707 $Y2=1.495
cc_275 N_VPB_c_124_p N_A_481_107#_c_1629_n 0.0677031f $X=18.48 $Y=4.07 $X2=2.707
+ $Y2=1.495
cc_276 N_VPB_M1012_b N_A_481_107#_c_1632_n 0.00218078f $X=-0.33 $Y=1.885
+ $X2=2.707 $Y2=1.26
cc_277 VPB N_A_481_107#_c_1632_n 5.70856e-19 $X=0 $Y=3.955 $X2=2.707 $Y2=1.26
cc_278 N_VPB_c_124_p N_A_481_107#_c_1632_n 0.0114989f $X=18.48 $Y=4.07 $X2=2.707
+ $Y2=1.26
cc_279 N_VPB_M1012_b N_A_481_107#_c_1635_n 0.00456559f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_280 N_VPB_M1012_b N_A_481_107#_c_1636_n 0.0185309f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_281 N_VPB_M1012_b N_A_481_107#_c_1637_n 0.00335007f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_282 N_VPB_M1012_b N_A_481_107#_c_1615_n 0.00303457f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_283 N_VPB_M1012_b N_Q_c_1748_n 0.0639382f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_284 N_VPB_c_124_p N_Q_c_1748_n 0.00495073f $X=18.48 $Y=4.07 $X2=0 $Y2=0
cc_285 N_SCE_c_285_n N_A_30_107#_c_357_n 0.00118322f $X=2.525 $Y=1.58 $X2=0
+ $Y2=0
cc_286 N_SCE_c_288_n N_A_30_107#_c_357_n 0.038867f $X=2.8 $Y=1.26 $X2=0 $Y2=0
cc_287 N_SCE_M1031_g N_A_30_107#_c_350_n 0.0184028f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_288 N_SCE_c_301_p N_A_30_107#_c_352_n 0.034719f $X=0.73 $Y=1.66 $X2=18.48
+ $Y2=0
cc_289 N_SCE_M1031_g N_A_30_107#_c_352_n 0.0369641f $X=0.665 $Y=0.745 $X2=18.48
+ $Y2=0
cc_290 N_SCE_c_292_n N_A_30_107#_c_361_n 0.0172661f $X=0.665 $Y=2.735 $X2=0
+ $Y2=0
cc_291 N_SCE_c_296_n N_A_30_107#_c_361_n 0.00203586f $X=0.665 $Y=2.485 $X2=0
+ $Y2=0
cc_292 N_SCE_c_285_n N_A_30_107#_c_353_n 0.0948981f $X=2.525 $Y=1.58 $X2=9.36
+ $Y2=0.057
cc_293 N_SCE_c_301_p N_A_30_107#_c_353_n 0.0244093f $X=0.73 $Y=1.66 $X2=9.36
+ $Y2=0.057
cc_294 N_SCE_M1031_g N_A_30_107#_c_353_n 0.0310813f $X=0.665 $Y=0.745 $X2=9.36
+ $Y2=0.057
cc_295 N_SCE_c_289_n N_A_30_107#_c_353_n 0.0130212f $X=2.8 $Y=1.26 $X2=9.36
+ $Y2=0.057
cc_296 N_SCE_c_296_n N_A_30_107#_c_362_n 0.0806618f $X=0.665 $Y=2.485 $X2=0
+ $Y2=0
cc_297 N_SCE_c_301_p N_A_30_107#_c_362_n 0.0133261f $X=0.73 $Y=1.66 $X2=0 $Y2=0
cc_298 N_SCE_c_285_n N_A_30_107#_c_377_n 0.0165171f $X=2.525 $Y=1.58 $X2=0 $Y2=0
cc_299 N_SCE_c_288_n N_A_30_107#_c_377_n 9.90829e-19 $X=2.8 $Y=1.26 $X2=0 $Y2=0
cc_300 N_SCE_M1031_g N_A_30_107#_c_354_n 0.00626054f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_301 N_SCE_c_296_n N_A_30_107#_c_363_n 0.00513266f $X=0.665 $Y=2.485 $X2=0
+ $Y2=0
cc_302 N_SCE_c_285_n N_A_30_107#_M1007_g 0.00627809f $X=2.525 $Y=1.58 $X2=0
+ $Y2=0
cc_303 N_SCE_c_288_n N_A_30_107#_M1007_g 0.025306f $X=2.8 $Y=1.26 $X2=0 $Y2=0
cc_304 N_SCE_c_289_n N_A_30_107#_M1007_g 0.00565697f $X=2.8 $Y=1.26 $X2=0 $Y2=0
cc_305 N_SCE_c_290_n N_A_30_107#_M1007_g 0.0149147f $X=2.9 $Y=1.075 $X2=0 $Y2=0
cc_306 N_SCE_c_285_n N_D_M1006_g 0.0306036f $X=2.525 $Y=1.58 $X2=0 $Y2=0
cc_307 N_SCE_c_301_p N_D_M1006_g 0.00234193f $X=0.73 $Y=1.66 $X2=0 $Y2=0
cc_308 N_SCE_M1031_g N_D_M1006_g 0.0629152f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_309 N_SCE_c_296_n N_D_M1030_g 0.0831523f $X=0.665 $Y=2.485 $X2=0 $Y2=0
cc_310 N_SCE_c_296_n N_D_c_425_n 0.0263993f $X=0.665 $Y=2.485 $X2=0 $Y2=0
cc_311 N_SCE_c_285_n N_D_c_425_n 0.0195091f $X=2.525 $Y=1.58 $X2=0 $Y2=0
cc_312 N_SCE_c_288_n N_D_c_425_n 0.00732748f $X=2.8 $Y=1.26 $X2=0 $Y2=0
cc_313 N_SCE_c_296_n N_D_c_436_n 4.89178e-19 $X=0.665 $Y=2.485 $X2=0 $Y2=0
cc_314 N_SCE_c_285_n N_D_c_436_n 0.0245274f $X=2.525 $Y=1.58 $X2=0 $Y2=0
cc_315 N_SCE_c_288_n SCD 6.52614e-19 $X=2.8 $Y=1.26 $X2=0 $Y2=0
cc_316 N_SCE_c_290_n N_SCD_M1001_g 0.0912486f $X=2.9 $Y=1.075 $X2=0 $Y2=0
cc_317 N_SCE_c_292_n N_VPWR_c_1479_n 0.0371899f $X=0.665 $Y=2.735 $X2=0 $Y2=0
cc_318 N_SCE_c_294_n N_VPWR_c_1479_n 0.0412105f $X=1.445 $Y=2.735 $X2=0 $Y2=0
cc_319 N_SCE_c_296_n N_VPWR_c_1479_n 0.00260931f $X=0.665 $Y=2.485 $X2=0 $Y2=0
cc_320 N_SCE_c_292_n N_VPWR_c_1503_n 0.00697248f $X=0.665 $Y=2.735 $X2=0 $Y2=0
cc_321 N_SCE_c_294_n N_VPWR_c_1503_n 0.00426472f $X=1.445 $Y=2.735 $X2=0 $Y2=0
cc_322 N_SCE_c_289_n N_A_481_107#_c_1610_n 0.0123821f $X=2.8 $Y=1.26 $X2=0 $Y2=0
cc_323 N_SCE_c_290_n N_A_481_107#_c_1610_n 0.0288031f $X=2.9 $Y=1.075 $X2=0
+ $Y2=0
cc_324 N_SCE_c_288_n N_A_481_107#_c_1611_n 0.0212587f $X=2.8 $Y=1.26 $X2=0 $Y2=0
cc_325 N_SCE_c_289_n N_A_481_107#_c_1611_n 0.0470714f $X=2.8 $Y=1.26 $X2=0 $Y2=0
cc_326 N_SCE_c_290_n N_A_481_107#_c_1611_n 0.00529711f $X=2.9 $Y=1.075 $X2=0
+ $Y2=0
cc_327 N_SCE_c_285_n N_A_481_107#_c_1612_n 0.0036861f $X=2.525 $Y=1.58 $X2=0
+ $Y2=0
cc_328 N_SCE_c_288_n N_A_481_107#_c_1612_n 0.00174394f $X=2.8 $Y=1.26 $X2=0
+ $Y2=0
cc_329 N_SCE_c_289_n N_A_481_107#_c_1612_n 0.0120828f $X=2.8 $Y=1.26 $X2=0 $Y2=0
cc_330 N_SCE_c_290_n N_A_481_107#_c_1612_n 0.00822988f $X=2.9 $Y=1.075 $X2=0
+ $Y2=0
cc_331 N_SCE_c_294_n N_A_481_107#_c_1637_n 0.0012815f $X=1.445 $Y=2.735 $X2=0
+ $Y2=0
cc_332 N_SCE_M1031_g N_VGND_c_1760_n 0.0319645f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_333 N_SCE_c_290_n N_VGND_c_1762_n 0.00356734f $X=2.9 $Y=1.075 $X2=0 $Y2=0
cc_334 N_SCE_M1031_g N_VGND_c_1774_n 0.00624345f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_335 N_SCE_c_289_n N_VGND_c_1774_n 0.0011881f $X=2.8 $Y=1.26 $X2=0 $Y2=0
cc_336 N_SCE_c_290_n N_VGND_c_1774_n 0.0151013f $X=2.9 $Y=1.075 $X2=0 $Y2=0
cc_337 N_A_30_107#_c_353_n N_D_M1006_g 0.0300401f $X=2.09 $Y=1.23 $X2=0 $Y2=0
cc_338 N_A_30_107#_M1007_g N_D_M1006_g 0.0769671f $X=2.155 $Y=0.745 $X2=0 $Y2=0
cc_339 N_A_30_107#_M1017_g N_D_M1030_g 0.0162736f $X=2.935 $Y=3.055 $X2=0 $Y2=0
cc_340 N_A_30_107#_c_362_n N_D_M1030_g 0.0445849f $X=2.635 $Y=2.62 $X2=0 $Y2=0
cc_341 N_A_30_107#_c_357_n N_D_c_425_n 0.0493438f $X=2.935 $Y=2.715 $X2=0 $Y2=0
cc_342 N_A_30_107#_c_362_n N_D_c_425_n 0.00830226f $X=2.635 $Y=2.62 $X2=0 $Y2=0
cc_343 N_A_30_107#_c_377_n N_D_c_425_n 0.00263469f $X=2.8 $Y=2.18 $X2=0 $Y2=0
cc_344 N_A_30_107#_M1007_g N_D_c_425_n 0.0328631f $X=2.155 $Y=0.745 $X2=0 $Y2=0
cc_345 N_A_30_107#_c_357_n N_D_c_436_n 0.0011825f $X=2.935 $Y=2.715 $X2=0 $Y2=0
cc_346 N_A_30_107#_c_362_n N_D_c_436_n 0.0232944f $X=2.635 $Y=2.62 $X2=0 $Y2=0
cc_347 N_A_30_107#_c_377_n N_D_c_436_n 0.0136779f $X=2.8 $Y=2.18 $X2=0 $Y2=0
cc_348 N_A_30_107#_c_357_n N_SCD_M1001_g 0.0880664f $X=2.935 $Y=2.715 $X2=0
+ $Y2=0
cc_349 N_A_30_107#_c_361_n N_VPWR_c_1479_n 0.0303552f $X=0.275 $Y=3.055 $X2=0
+ $Y2=0
cc_350 N_A_30_107#_c_362_n N_VPWR_c_1479_n 0.0647546f $X=2.635 $Y=2.62 $X2=0
+ $Y2=0
cc_351 N_A_30_107#_M1017_g N_VPWR_c_1482_n 0.00261351f $X=2.935 $Y=3.055 $X2=0
+ $Y2=0
cc_352 N_A_30_107#_M1017_g N_VPWR_c_1503_n 0.0169235f $X=2.935 $Y=3.055 $X2=0
+ $Y2=0
cc_353 N_A_30_107#_c_361_n N_VPWR_c_1503_n 0.018898f $X=0.275 $Y=3.055 $X2=0
+ $Y2=0
cc_354 N_A_30_107#_M1017_g N_A_481_107#_c_1649_n 0.0278784f $X=2.935 $Y=3.055
+ $X2=0 $Y2=0
cc_355 N_A_30_107#_c_362_n N_A_481_107#_c_1649_n 0.0131097f $X=2.635 $Y=2.62
+ $X2=0 $Y2=0
cc_356 N_A_30_107#_c_357_n N_A_481_107#_c_1611_n 0.013655f $X=2.935 $Y=2.715
+ $X2=0 $Y2=0
cc_357 N_A_30_107#_c_377_n N_A_481_107#_c_1611_n 0.0293705f $X=2.8 $Y=2.18 $X2=0
+ $Y2=0
cc_358 N_A_30_107#_M1007_g N_A_481_107#_c_1611_n 6.52142e-19 $X=2.155 $Y=0.745
+ $X2=0 $Y2=0
cc_359 N_A_30_107#_c_357_n N_A_481_107#_c_1617_n 0.00248729f $X=2.935 $Y=2.715
+ $X2=0 $Y2=0
cc_360 N_A_30_107#_M1017_g N_A_481_107#_c_1617_n 0.00563237f $X=2.935 $Y=3.055
+ $X2=0 $Y2=0
cc_361 N_A_30_107#_c_362_n N_A_481_107#_c_1617_n 0.00578689f $X=2.635 $Y=2.62
+ $X2=0 $Y2=0
cc_362 N_A_30_107#_M1007_g N_A_481_107#_c_1612_n 0.0116924f $X=2.155 $Y=0.745
+ $X2=0 $Y2=0
cc_363 N_A_30_107#_c_357_n N_A_481_107#_c_1637_n 0.00173043f $X=2.935 $Y=2.715
+ $X2=0 $Y2=0
cc_364 N_A_30_107#_M1017_g N_A_481_107#_c_1637_n 0.00829232f $X=2.935 $Y=3.055
+ $X2=0 $Y2=0
cc_365 N_A_30_107#_c_362_n N_A_481_107#_c_1637_n 0.0203888f $X=2.635 $Y=2.62
+ $X2=0 $Y2=0
cc_366 N_A_30_107#_c_357_n N_A_481_107#_c_1661_n 0.00584954f $X=2.935 $Y=2.715
+ $X2=0 $Y2=0
cc_367 N_A_30_107#_c_362_n N_A_481_107#_c_1661_n 0.00727324f $X=2.635 $Y=2.62
+ $X2=0 $Y2=0
cc_368 N_A_30_107#_c_377_n N_A_481_107#_c_1661_n 0.00595203f $X=2.8 $Y=2.18
+ $X2=0 $Y2=0
cc_369 N_A_30_107#_c_350_n N_VGND_c_1760_n 0.0287634f $X=0.275 $Y=0.745 $X2=0
+ $Y2=0
cc_370 N_A_30_107#_c_353_n N_VGND_c_1760_n 0.0630617f $X=2.09 $Y=1.23 $X2=0
+ $Y2=0
cc_371 N_A_30_107#_M1007_g N_VGND_c_1760_n 0.00362967f $X=2.155 $Y=0.745 $X2=0
+ $Y2=0
cc_372 N_A_30_107#_c_350_n N_VGND_c_1774_n 0.0319953f $X=0.275 $Y=0.745 $X2=0
+ $Y2=0
cc_373 N_A_30_107#_c_353_n N_VGND_c_1774_n 0.0321069f $X=2.09 $Y=1.23 $X2=0
+ $Y2=0
cc_374 N_A_30_107#_M1007_g N_VGND_c_1774_n 0.0212499f $X=2.155 $Y=0.745 $X2=0
+ $Y2=0
cc_375 N_D_M1030_g N_VPWR_c_1479_n 0.0028297f $X=2.155 $Y=3.055 $X2=0 $Y2=0
cc_376 N_D_M1030_g N_VPWR_c_1503_n 0.0169235f $X=2.155 $Y=3.055 $X2=0 $Y2=0
cc_377 N_D_c_425_n N_A_481_107#_c_1611_n 0.00540326f $X=2.11 $Y=1.93 $X2=0 $Y2=0
cc_378 N_D_M1030_g N_A_481_107#_c_1617_n 6.24781e-19 $X=2.155 $Y=3.055 $X2=0
+ $Y2=0
cc_379 N_D_M1006_g N_A_481_107#_c_1612_n 0.0014684f $X=1.445 $Y=0.745 $X2=0
+ $Y2=0
cc_380 N_D_M1030_g N_A_481_107#_c_1637_n 0.0115244f $X=2.155 $Y=3.055 $X2=0
+ $Y2=0
cc_381 N_D_M1006_g N_VGND_c_1760_n 0.0397166f $X=1.445 $Y=0.745 $X2=0 $Y2=0
cc_382 N_D_M1006_g N_VGND_c_1774_n 0.00445548f $X=1.445 $Y=0.745 $X2=0 $Y2=0
cc_383 N_SCD_M1001_g N_CLK_M1028_g 0.0958755f $X=3.645 $Y=0.745 $X2=0 $Y2=0
cc_384 N_SCD_M1001_g N_CLK_c_488_n 0.0132777f $X=3.645 $Y=0.745 $X2=0.24 $Y2=0
cc_385 SCD CLK 0.067581f $X=3.515 $Y=1.21 $X2=0.24 $Y2=0
cc_386 N_SCD_M1001_g CLK 0.00950814f $X=3.645 $Y=0.745 $X2=0.24 $Y2=0
cc_387 SCD N_CLK_c_486_n 7.30243e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_388 N_SCD_M1001_g N_VPWR_c_1482_n 0.0584291f $X=3.645 $Y=0.745 $X2=0 $Y2=0
cc_389 N_SCD_M1001_g N_VPWR_c_1503_n 8.80022e-19 $X=3.645 $Y=0.745 $X2=0 $Y2=0
cc_390 SCD N_A_481_107#_c_1611_n 0.070186f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_391 N_SCD_M1001_g N_A_481_107#_c_1611_n 0.0205596f $X=3.645 $Y=0.745 $X2=0
+ $Y2=0
cc_392 N_SCD_M1001_g N_A_481_107#_c_1617_n 0.00415436f $X=3.645 $Y=0.745 $X2=0
+ $Y2=0
cc_393 SCD N_A_481_107#_c_1618_n 0.015622f $X=3.515 $Y=1.21 $X2=9.36 $Y2=0
cc_394 N_SCD_M1001_g N_A_481_107#_c_1618_n 0.0330127f $X=3.645 $Y=0.745 $X2=9.36
+ $Y2=0
cc_395 N_SCD_M1001_g N_A_481_107#_c_1673_n 0.00110166f $X=3.645 $Y=0.745 $X2=0
+ $Y2=0
cc_396 N_SCD_M1001_g N_A_481_107#_c_1612_n 9.53229e-19 $X=3.645 $Y=0.745 $X2=0
+ $Y2=0
cc_397 N_SCD_M1001_g N_A_481_107#_c_1637_n 7.66324e-19 $X=3.645 $Y=0.745 $X2=0
+ $Y2=0
cc_398 SCD N_VGND_c_1762_n 0.0254652f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_399 N_SCD_M1001_g N_VGND_c_1762_n 0.05491f $X=3.645 $Y=0.745 $X2=0 $Y2=0
cc_400 SCD N_VGND_c_1774_n 0.00119919f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_401 N_SCD_M1001_g N_VGND_c_1774_n 0.00254032f $X=3.645 $Y=0.745 $X2=0 $Y2=0
cc_402 N_CLK_c_484_n N_A_935_107#_c_542_n 0.0078306f $X=4.482 $Y=2.428 $X2=0
+ $Y2=0
cc_403 N_CLK_M1028_g N_A_935_107#_c_522_n 0.00408753f $X=4.425 $Y=0.745 $X2=0
+ $Y2=0
cc_404 CLK N_A_935_107#_c_522_n 0.0272446f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_405 N_CLK_c_486_n N_A_935_107#_c_522_n 0.0125457f $X=4.36 $Y=1.34 $X2=0 $Y2=0
cc_406 N_CLK_c_484_n N_A_935_107#_c_551_n 0.0293737f $X=4.482 $Y=2.428 $X2=0
+ $Y2=0
cc_407 CLK N_A_935_107#_c_551_n 0.0119166f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_408 N_CLK_M1028_g N_A_935_107#_c_532_n 0.0116555f $X=4.425 $Y=0.745 $X2=0
+ $Y2=0
cc_409 N_CLK_c_486_n N_A_935_107#_c_532_n 0.00565049f $X=4.36 $Y=1.34 $X2=0
+ $Y2=0
cc_410 N_CLK_c_484_n N_A_935_107#_c_534_n 0.0032677f $X=4.482 $Y=2.428 $X2=0
+ $Y2=0
cc_411 CLK N_A_935_107#_c_534_n 0.00927024f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_412 N_CLK_c_486_n N_A_935_107#_M1002_g 0.0078306f $X=4.36 $Y=1.34 $X2=0 $Y2=0
cc_413 N_CLK_c_488_n N_VPWR_c_1482_n 0.0226259f $X=4.482 $Y=2.735 $X2=0 $Y2=0
cc_414 N_CLK_c_488_n N_VPWR_c_1503_n 0.0192867f $X=4.482 $Y=2.735 $X2=0 $Y2=0
cc_415 N_CLK_c_488_n N_A_481_107#_c_1618_n 0.0343869f $X=4.482 $Y=2.735 $X2=9.36
+ $Y2=0
cc_416 CLK N_A_481_107#_c_1618_n 0.028501f $X=3.995 $Y=1.21 $X2=9.36 $Y2=0
cc_417 N_CLK_c_488_n N_A_481_107#_c_1673_n 0.0386021f $X=4.482 $Y=2.735 $X2=0
+ $Y2=0
cc_418 N_CLK_c_488_n N_A_481_107#_c_1619_n 0.00802989f $X=4.482 $Y=2.735 $X2=0
+ $Y2=0
cc_419 N_CLK_c_488_n N_A_481_107#_c_1622_n 0.00508647f $X=4.482 $Y=2.735 $X2=0
+ $Y2=0
cc_420 N_CLK_c_488_n N_A_481_107#_c_1625_n 0.00381613f $X=4.482 $Y=2.735 $X2=0
+ $Y2=0
cc_421 N_CLK_M1028_g N_VGND_c_1762_n 0.0296175f $X=4.425 $Y=0.745 $X2=0 $Y2=0
cc_422 CLK N_VGND_c_1762_n 0.0331243f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_423 N_CLK_M1028_g N_VGND_c_1764_n 0.00247214f $X=4.425 $Y=0.745 $X2=0 $Y2=0
cc_424 N_CLK_M1028_g N_VGND_c_1774_n 0.0140086f $X=4.425 $Y=0.745 $X2=0 $Y2=0
cc_425 CLK N_VGND_c_1774_n 0.00656154f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_426 N_A_935_107#_M1026_g N_A_1201_123#_M1004_g 0.0134958f $X=8.18 $Y=2.925
+ $X2=0 $Y2=0
cc_427 N_A_935_107#_c_528_n N_A_1201_123#_M1004_g 0.0297975f $X=7.36 $Y=3.355
+ $X2=0 $Y2=0
cc_428 N_A_935_107#_c_554_n N_A_1201_123#_M1004_g 0.00887434f $X=8.135 $Y=3.44
+ $X2=0 $Y2=0
cc_429 N_A_935_107#_c_561_n N_A_1201_123#_M1004_g 5.62571e-19 $X=8.22 $Y=3.355
+ $X2=0 $Y2=0
cc_430 N_A_935_107#_c_586_p N_A_1201_123#_M1024_g 0.00101071f $X=7.145 $Y=1.27
+ $X2=0 $Y2=0
cc_431 N_A_935_107#_M1034_g N_A_1201_123#_M1024_g 0.0138865f $X=7.105 $Y=0.775
+ $X2=0 $Y2=0
cc_432 N_A_935_107#_c_521_n N_A_1201_123#_M1013_g 0.0246985f $X=13.095 $Y=1.395
+ $X2=18.48 $Y2=0
cc_433 N_A_935_107#_c_589_p N_A_1201_123#_M1013_g 0.025526f $X=12.18 $Y=1.335
+ $X2=18.48 $Y2=0
cc_434 N_A_935_107#_c_529_n N_A_1201_123#_M1013_g 0.013451f $X=13.1 $Y=0.7
+ $X2=18.48 $Y2=0
cc_435 N_A_935_107#_c_591_p N_A_1201_123#_M1013_g 0.00634335f $X=12.265 $Y=0.7
+ $X2=18.48 $Y2=0
cc_436 N_A_935_107#_c_530_n N_A_1201_123#_M1013_g 0.0104243f $X=12.485 $Y=2.225
+ $X2=18.48 $Y2=0
cc_437 N_A_935_107#_c_531_n N_A_1201_123#_M1013_g 5.35057e-19 $X=13.185 $Y=1.58
+ $X2=18.48 $Y2=0
cc_438 N_A_935_107#_c_537_n N_A_1201_123#_M1013_g 0.0249527f $X=12.485 $Y=1.42
+ $X2=18.48 $Y2=0
cc_439 N_A_935_107#_M1019_g N_A_1201_123#_c_801_n 0.0103425f $X=12.135 $Y=3.215
+ $X2=0 $Y2=0
cc_440 N_A_935_107#_c_523_n N_A_1201_123#_c_792_n 0.00928991f $X=5.505 $Y=1.82
+ $X2=0 $Y2=0
cc_441 N_A_935_107#_c_542_n N_A_1201_123#_c_802_n 0.0242094f $X=6.03 $Y=2.555
+ $X2=0 $Y2=0
cc_442 N_A_935_107#_M1002_g N_A_1201_123#_c_802_n 0.00328751f $X=5.755 $Y=0.825
+ $X2=0 $Y2=0
cc_443 N_A_935_107#_c_545_n N_A_1201_123#_c_793_n 0.00126784f $X=12.135 $Y=2.565
+ $X2=0 $Y2=0
cc_444 N_A_935_107#_c_600_p N_A_1201_123#_c_793_n 0.00779006f $X=8.245 $Y=2.39
+ $X2=0 $Y2=0
cc_445 N_A_935_107#_c_560_n N_A_1201_123#_c_793_n 0.00300435f $X=8.245 $Y=2.39
+ $X2=0 $Y2=0
cc_446 N_A_935_107#_c_562_n N_A_1201_123#_c_793_n 0.0117682f $X=9.625 $Y=2.66
+ $X2=0 $Y2=0
cc_447 N_A_935_107#_c_565_n N_A_1201_123#_c_793_n 0.00497349f $X=12.042 $Y=2.395
+ $X2=0 $Y2=0
cc_448 N_A_935_107#_c_524_n N_A_1201_123#_c_794_n 0.0142774f $X=7.06 $Y=0.35
+ $X2=0 $Y2=0
cc_449 N_A_935_107#_c_535_n N_A_1201_123#_c_794_n 0.025921f $X=5.67 $Y=1.235
+ $X2=0 $Y2=0
cc_450 N_A_935_107#_M1002_g N_A_1201_123#_c_794_n 0.00846629f $X=5.755 $Y=0.825
+ $X2=0 $Y2=0
cc_451 N_A_935_107#_M1034_g N_A_1201_123#_c_794_n 0.00246195f $X=7.105 $Y=0.775
+ $X2=0 $Y2=0
cc_452 N_A_935_107#_c_608_p N_A_1201_123#_c_795_n 0.0126109f $X=5.67 $Y=1.735
+ $X2=0 $Y2=0
cc_453 N_A_935_107#_M1034_g N_A_1201_123#_c_795_n 2.7862e-19 $X=7.105 $Y=0.775
+ $X2=0 $Y2=0
cc_454 N_A_935_107#_c_608_p N_A_1201_123#_c_796_n 2.93944e-19 $X=5.67 $Y=1.735
+ $X2=0 $Y2=0
cc_455 N_A_935_107#_M1002_g N_A_1201_123#_c_796_n 0.0502843f $X=5.755 $Y=0.825
+ $X2=0 $Y2=0
cc_456 N_A_935_107#_M1034_g N_A_1201_123#_c_796_n 0.0233509f $X=7.105 $Y=0.775
+ $X2=0 $Y2=0
cc_457 N_A_935_107#_c_613_p N_A_1201_123#_c_797_n 0.0126109f $X=5.67 $Y=1.4
+ $X2=0 $Y2=0
cc_458 N_A_935_107#_c_535_n N_A_1201_123#_c_797_n 0.0076403f $X=5.67 $Y=1.235
+ $X2=0 $Y2=0
cc_459 N_A_935_107#_M1002_g N_A_1201_123#_c_797_n 0.0185701f $X=5.755 $Y=0.825
+ $X2=0 $Y2=0
cc_460 N_A_935_107#_c_542_n N_A_1201_123#_c_805_n 0.00340288f $X=6.03 $Y=2.555
+ $X2=0 $Y2=0
cc_461 N_A_935_107#_M1026_g N_A_1201_123#_c_806_n 0.00192468f $X=8.18 $Y=2.925
+ $X2=0 $Y2=0
cc_462 N_A_935_107#_c_600_p N_A_1201_123#_c_806_n 0.0135931f $X=8.245 $Y=2.39
+ $X2=0 $Y2=0
cc_463 N_A_935_107#_c_560_n N_A_1201_123#_c_806_n 0.0024389f $X=8.245 $Y=2.39
+ $X2=0 $Y2=0
cc_464 N_A_935_107#_c_545_n N_A_1201_123#_c_807_n 9.51131e-19 $X=12.135 $Y=2.565
+ $X2=0 $Y2=0
cc_465 N_A_935_107#_c_565_n N_A_1201_123#_c_807_n 0.016984f $X=12.042 $Y=2.395
+ $X2=0 $Y2=0
cc_466 N_A_935_107#_c_566_n N_A_1201_123#_c_807_n 0.00282274f $X=12.4 $Y=2.31
+ $X2=0 $Y2=0
cc_467 N_A_935_107#_c_530_n N_A_1201_123#_c_807_n 0.0241859f $X=12.485 $Y=2.225
+ $X2=0 $Y2=0
cc_468 N_A_935_107#_c_537_n N_A_1201_123#_c_807_n 0.00855996f $X=12.485 $Y=1.42
+ $X2=0 $Y2=0
cc_469 N_A_935_107#_c_545_n N_A_1201_123#_c_798_n 0.0477133f $X=12.135 $Y=2.565
+ $X2=0 $Y2=0
cc_470 N_A_935_107#_c_521_n N_A_1201_123#_c_798_n 0.0267418f $X=13.095 $Y=1.395
+ $X2=0 $Y2=0
cc_471 N_A_935_107#_c_565_n N_A_1201_123#_c_798_n 2.41999e-19 $X=12.042 $Y=2.395
+ $X2=0 $Y2=0
cc_472 N_A_935_107#_c_628_p N_A_1201_123#_c_798_n 6.52562e-19 $X=12.042 $Y=2.935
+ $X2=0 $Y2=0
cc_473 N_A_935_107#_c_566_n N_A_1201_123#_c_798_n 0.00546778f $X=12.4 $Y=2.31
+ $X2=0 $Y2=0
cc_474 N_A_935_107#_c_530_n N_A_1201_123#_c_798_n 0.0215871f $X=12.485 $Y=2.225
+ $X2=0 $Y2=0
cc_475 N_A_935_107#_c_537_n N_A_1201_123#_c_798_n 3.33999e-19 $X=12.485 $Y=1.42
+ $X2=0 $Y2=0
cc_476 N_A_935_107#_c_542_n N_A_1201_123#_c_799_n 0.0177825f $X=6.03 $Y=2.555
+ $X2=0 $Y2=0
cc_477 N_A_935_107#_M1026_g N_A_1201_123#_c_799_n 0.00310683f $X=8.18 $Y=2.925
+ $X2=0 $Y2=0
cc_478 N_A_935_107#_c_586_p N_A_1201_123#_c_799_n 0.00162491f $X=7.145 $Y=1.27
+ $X2=0 $Y2=0
cc_479 N_A_935_107#_c_528_n N_A_1201_123#_c_799_n 0.039074f $X=7.36 $Y=3.355
+ $X2=0 $Y2=0
cc_480 N_A_935_107#_c_600_p N_A_1201_123#_c_799_n 9.79966e-19 $X=8.245 $Y=2.39
+ $X2=0 $Y2=0
cc_481 N_A_935_107#_c_560_n N_A_1201_123#_c_799_n 0.0324128f $X=8.245 $Y=2.39
+ $X2=0 $Y2=0
cc_482 N_A_935_107#_c_536_n N_A_1201_123#_c_799_n 0.00328815f $X=7.36 $Y=1.69
+ $X2=0 $Y2=0
cc_483 N_A_935_107#_M1002_g N_A_1201_123#_c_799_n 0.00427596f $X=5.755 $Y=0.825
+ $X2=0 $Y2=0
cc_484 N_A_935_107#_M1034_g N_A_1201_123#_c_799_n 0.081149f $X=7.105 $Y=0.775
+ $X2=0 $Y2=0
cc_485 N_A_935_107#_c_563_n N_A_1669_87#_M1018_d 0.00180746f $X=10.485 $Y=3.19
+ $X2=0 $Y2=0
cc_486 N_A_935_107#_c_600_p N_A_1669_87#_c_954_n 0.00691291f $X=8.245 $Y=2.39
+ $X2=0.24 $Y2=0
cc_487 N_A_935_107#_c_560_n N_A_1669_87#_c_954_n 4.76317e-19 $X=8.245 $Y=2.39
+ $X2=0.24 $Y2=0
cc_488 N_A_935_107#_c_562_n N_A_1669_87#_c_954_n 0.0691553f $X=9.625 $Y=2.66
+ $X2=0.24 $Y2=0
cc_489 N_A_935_107#_c_600_p N_A_1669_87#_c_949_n 0.00195909f $X=8.245 $Y=2.39
+ $X2=0 $Y2=0
cc_490 N_A_935_107#_c_560_n N_A_1669_87#_c_949_n 0.070866f $X=8.245 $Y=2.39
+ $X2=0 $Y2=0
cc_491 N_A_935_107#_c_561_n N_A_1669_87#_c_949_n 0.00128819f $X=8.22 $Y=3.355
+ $X2=0 $Y2=0
cc_492 N_A_935_107#_c_562_n N_A_1669_87#_c_949_n 0.0276333f $X=9.625 $Y=2.66
+ $X2=0 $Y2=0
cc_493 N_A_935_107#_c_649_p N_A_1669_87#_c_949_n 6.43668e-19 $X=9.71 $Y=3.105
+ $X2=0 $Y2=0
cc_494 N_A_935_107#_c_562_n N_A_1669_87#_c_965_n 0.0129587f $X=9.625 $Y=2.66
+ $X2=9.36 $Y2=0.057
cc_495 N_A_935_107#_c_649_p N_A_1669_87#_c_965_n 0.012246f $X=9.71 $Y=3.105
+ $X2=9.36 $Y2=0.057
cc_496 N_A_935_107#_c_563_n N_A_1669_87#_c_965_n 0.0157078f $X=10.485 $Y=3.19
+ $X2=9.36 $Y2=0.057
cc_497 N_A_935_107#_c_545_n N_A_1471_113#_M1016_g 0.114215f $X=12.135 $Y=2.565
+ $X2=0 $Y2=0
cc_498 N_A_935_107#_c_654_p N_A_1471_113#_M1016_g 0.0410852f $X=11.905 $Y=3.02
+ $X2=0 $Y2=0
cc_499 N_A_935_107#_c_565_n N_A_1471_113#_M1016_g 0.00119133f $X=12.042 $Y=2.395
+ $X2=0 $Y2=0
cc_500 N_A_935_107#_c_628_p N_A_1471_113#_M1016_g 0.00381137f $X=12.042 $Y=2.935
+ $X2=0 $Y2=0
cc_501 N_A_935_107#_c_569_n N_A_1471_113#_M1016_g 0.00122364f $X=10.57 $Y=3.02
+ $X2=0 $Y2=0
cc_502 N_A_935_107#_c_589_p N_A_1471_113#_M1011_g 0.00183039f $X=12.18 $Y=1.335
+ $X2=18.48 $Y2=0
cc_503 N_A_935_107#_c_591_p N_A_1471_113#_M1011_g 5.648e-19 $X=12.265 $Y=0.7
+ $X2=18.48 $Y2=0
cc_504 N_A_935_107#_c_537_n N_A_1471_113#_M1011_g 9.24487e-19 $X=12.485 $Y=1.42
+ $X2=18.48 $Y2=0
cc_505 N_A_935_107#_c_586_p N_A_1471_113#_c_1014_n 0.0116664f $X=7.145 $Y=1.27
+ $X2=0 $Y2=0
cc_506 N_A_935_107#_M1034_g N_A_1471_113#_c_1014_n 0.0015779f $X=7.105 $Y=0.775
+ $X2=0 $Y2=0
cc_507 N_A_935_107#_M1026_g N_A_1471_113#_c_1026_n 0.00383774f $X=8.18 $Y=2.925
+ $X2=0 $Y2=0
cc_508 N_A_935_107#_c_561_n N_A_1471_113#_c_1026_n 0.0292634f $X=8.22 $Y=3.355
+ $X2=0 $Y2=0
cc_509 N_A_935_107#_c_665_p N_A_1471_113#_c_1026_n 0.00533593f $X=8.272 $Y=2.66
+ $X2=0 $Y2=0
cc_510 N_A_935_107#_M1026_g N_A_1471_113#_c_1027_n 0.00629349f $X=8.18 $Y=2.925
+ $X2=0 $Y2=0
cc_511 N_A_935_107#_c_554_n N_A_1471_113#_c_1027_n 0.0237347f $X=8.135 $Y=3.44
+ $X2=0 $Y2=0
cc_512 N_A_935_107#_c_530_n N_A_1471_113#_c_1017_n 6.37081e-19 $X=12.485
+ $Y=2.225 $X2=0 $Y2=0
cc_513 N_A_935_107#_c_586_p N_A_1471_113#_c_1018_n 0.0199238f $X=7.145 $Y=1.27
+ $X2=0 $Y2=0
cc_514 N_A_935_107#_c_536_n N_A_1471_113#_c_1018_n 0.00122374f $X=7.36 $Y=1.69
+ $X2=0 $Y2=0
cc_515 N_A_935_107#_M1034_g N_A_1471_113#_c_1018_n 8.49365e-19 $X=7.105 $Y=0.775
+ $X2=0 $Y2=0
cc_516 N_A_935_107#_c_586_p N_A_1471_113#_c_1050_n 0.00654906f $X=7.145 $Y=1.27
+ $X2=0 $Y2=0
cc_517 N_A_935_107#_M1034_g N_A_1471_113#_c_1050_n 6.36459e-19 $X=7.105 $Y=0.775
+ $X2=0 $Y2=0
cc_518 N_A_935_107#_M1026_g N_A_1471_113#_c_1029_n 8.12473e-19 $X=8.18 $Y=2.925
+ $X2=0 $Y2=0
cc_519 N_A_935_107#_c_586_p N_A_1471_113#_c_1029_n 0.00273232f $X=7.145 $Y=1.27
+ $X2=0 $Y2=0
cc_520 N_A_935_107#_c_528_n N_A_1471_113#_c_1029_n 0.0930345f $X=7.36 $Y=3.355
+ $X2=0 $Y2=0
cc_521 N_A_935_107#_c_600_p N_A_1471_113#_c_1029_n 0.0148783f $X=8.245 $Y=2.39
+ $X2=0 $Y2=0
cc_522 N_A_935_107#_c_560_n N_A_1471_113#_c_1029_n 0.00226616f $X=8.245 $Y=2.39
+ $X2=0 $Y2=0
cc_523 N_A_935_107#_c_536_n N_A_1471_113#_c_1029_n 0.0123678f $X=7.36 $Y=1.69
+ $X2=0 $Y2=0
cc_524 N_A_935_107#_c_665_p N_A_1471_113#_c_1029_n 0.00469284f $X=8.272 $Y=2.66
+ $X2=0 $Y2=0
cc_525 N_A_935_107#_M1034_g N_A_1471_113#_c_1029_n 4.69619e-19 $X=7.105 $Y=0.775
+ $X2=0 $Y2=0
cc_526 N_A_935_107#_c_562_n N_A_1471_113#_c_1021_n 0.0190146f $X=9.625 $Y=2.66
+ $X2=0 $Y2=0
cc_527 N_A_935_107#_c_649_p N_A_1471_113#_c_1021_n 0.0153426f $X=9.71 $Y=3.105
+ $X2=0 $Y2=0
cc_528 N_A_935_107#_c_563_n N_A_1471_113#_c_1021_n 0.0160918f $X=10.485 $Y=3.19
+ $X2=0 $Y2=0
cc_529 N_A_935_107#_c_564_n N_A_1471_113#_c_1021_n 0.00626001f $X=9.795 $Y=3.19
+ $X2=0 $Y2=0
cc_530 N_A_935_107#_c_569_n N_A_1471_113#_c_1021_n 6.40009e-19 $X=10.57 $Y=3.02
+ $X2=0 $Y2=0
cc_531 N_A_935_107#_c_649_p N_SET_B_c_1156_n 5.99284e-19 $X=9.71 $Y=3.105 $X2=0
+ $Y2=0
cc_532 N_A_935_107#_c_563_n N_SET_B_c_1156_n 0.0171342f $X=10.485 $Y=3.19 $X2=0
+ $Y2=0
cc_533 N_A_935_107#_c_654_p N_SET_B_c_1156_n 0.0160081f $X=11.905 $Y=3.02 $X2=0
+ $Y2=0
cc_534 N_A_935_107#_c_569_n N_SET_B_c_1156_n 0.0220842f $X=10.57 $Y=3.02 $X2=0
+ $Y2=0
cc_535 N_A_935_107#_c_589_p N_SET_B_c_1146_n 0.00541825f $X=12.18 $Y=1.335 $X2=0
+ $Y2=0
cc_536 N_A_935_107#_c_537_n N_SET_B_c_1146_n 3.28736e-19 $X=12.485 $Y=1.42 $X2=0
+ $Y2=0
cc_537 N_A_935_107#_c_589_p N_SET_B_c_1165_n 0.0117551f $X=12.18 $Y=1.335 $X2=0
+ $Y2=0
cc_538 N_A_935_107#_c_591_p N_SET_B_c_1165_n 0.0055995f $X=12.265 $Y=0.7 $X2=0
+ $Y2=0
cc_539 N_A_935_107#_c_521_n N_SET_B_c_1147_n 0.00232685f $X=13.095 $Y=1.395
+ $X2=0 $Y2=0
cc_540 N_A_935_107#_c_529_n N_SET_B_c_1147_n 0.0703948f $X=13.1 $Y=0.7 $X2=0
+ $Y2=0
cc_541 N_A_935_107#_c_591_p N_SET_B_c_1147_n 0.0104792f $X=12.265 $Y=0.7 $X2=0
+ $Y2=0
cc_542 N_A_935_107#_c_521_n SET_B 0.00107495f $X=13.095 $Y=1.395 $X2=0 $Y2=0
cc_543 N_A_935_107#_c_521_n N_A_2698_421#_M1014_g 0.0769759f $X=13.095 $Y=1.395
+ $X2=0 $Y2=0
cc_544 N_A_935_107#_c_529_n N_A_2698_421#_M1014_g 0.00131888f $X=13.1 $Y=0.7
+ $X2=0 $Y2=0
cc_545 N_A_935_107#_c_531_n N_A_2698_421#_M1014_g 0.00795273f $X=13.185 $Y=1.58
+ $X2=0 $Y2=0
cc_546 N_A_935_107#_c_529_n N_A_2477_543#_M1013_d 0.00345369f $X=13.1 $Y=0.7
+ $X2=0 $Y2=0
cc_547 N_A_935_107#_M1019_g N_A_2477_543#_c_1318_n 0.0197231f $X=12.135 $Y=3.215
+ $X2=0 $Y2=0
cc_548 N_A_935_107#_c_654_p N_A_2477_543#_c_1318_n 0.0129587f $X=11.905 $Y=3.02
+ $X2=0 $Y2=0
cc_549 N_A_935_107#_c_628_p N_A_2477_543#_c_1318_n 0.00632773f $X=12.042
+ $Y=2.935 $X2=0 $Y2=0
cc_550 N_A_935_107#_c_521_n N_A_2477_543#_c_1332_n 0.00796177f $X=13.095
+ $Y=1.395 $X2=0 $Y2=0
cc_551 N_A_935_107#_c_589_p N_A_2477_543#_c_1332_n 0.0132738f $X=12.18 $Y=1.335
+ $X2=0 $Y2=0
cc_552 N_A_935_107#_c_529_n N_A_2477_543#_c_1332_n 0.0259654f $X=13.1 $Y=0.7
+ $X2=0 $Y2=0
cc_553 N_A_935_107#_c_531_n N_A_2477_543#_c_1332_n 0.0137965f $X=13.185 $Y=1.58
+ $X2=0 $Y2=0
cc_554 N_A_935_107#_c_537_n N_A_2477_543#_c_1332_n 0.00673784f $X=12.485 $Y=1.42
+ $X2=0 $Y2=0
cc_555 N_A_935_107#_c_521_n N_A_2477_543#_c_1310_n 0.0193287f $X=13.095 $Y=1.395
+ $X2=0 $Y2=0
cc_556 N_A_935_107#_c_589_p N_A_2477_543#_c_1310_n 0.00566112f $X=12.18 $Y=1.335
+ $X2=0 $Y2=0
cc_557 N_A_935_107#_c_530_n N_A_2477_543#_c_1310_n 0.0304408f $X=12.485 $Y=2.225
+ $X2=0 $Y2=0
cc_558 N_A_935_107#_c_531_n N_A_2477_543#_c_1310_n 0.0398118f $X=13.185 $Y=1.58
+ $X2=0 $Y2=0
cc_559 N_A_935_107#_c_537_n N_A_2477_543#_c_1310_n 0.0132276f $X=12.485 $Y=1.42
+ $X2=0 $Y2=0
cc_560 N_A_935_107#_c_545_n N_A_2477_543#_c_1322_n 8.05076e-19 $X=12.135
+ $Y=2.565 $X2=0 $Y2=0
cc_561 N_A_935_107#_M1019_g N_A_2477_543#_c_1322_n 6.01121e-19 $X=12.135
+ $Y=3.215 $X2=0 $Y2=0
cc_562 N_A_935_107#_c_628_p N_A_2477_543#_c_1322_n 0.00750395f $X=12.042
+ $Y=2.935 $X2=0 $Y2=0
cc_563 N_A_935_107#_c_566_n N_A_2477_543#_c_1322_n 0.013112f $X=12.4 $Y=2.31
+ $X2=0 $Y2=0
cc_564 N_A_935_107#_c_530_n N_A_2477_543#_c_1322_n 0.00780963f $X=12.485
+ $Y=2.225 $X2=0 $Y2=0
cc_565 N_A_935_107#_M1019_g N_A_2477_543#_c_1325_n 0.00390331f $X=12.135
+ $Y=3.215 $X2=0 $Y2=0
cc_566 N_A_935_107#_c_628_p N_A_2477_543#_c_1325_n 0.0124429f $X=12.042 $Y=2.935
+ $X2=0 $Y2=0
cc_567 N_A_935_107#_c_566_n N_A_2477_543#_c_1325_n 0.0120452f $X=12.4 $Y=2.31
+ $X2=0 $Y2=0
cc_568 N_A_935_107#_c_530_n N_A_2477_543#_c_1350_n 0.012385f $X=12.485 $Y=2.225
+ $X2=0 $Y2=0
cc_569 N_A_935_107#_c_521_n N_A_2477_543#_c_1326_n 0.00768775f $X=13.095
+ $Y=1.395 $X2=0 $Y2=0
cc_570 N_A_935_107#_c_531_n N_A_2477_543#_c_1326_n 0.0178555f $X=13.185 $Y=1.58
+ $X2=0 $Y2=0
cc_571 N_A_935_107#_c_562_n N_VPWR_M1000_d 0.00267852f $X=9.625 $Y=2.66 $X2=0
+ $Y2=0
cc_572 N_A_935_107#_c_654_p N_VPWR_M1027_d 0.0127626f $X=11.905 $Y=3.02
+ $X2=-0.33 $Y2=-0.265
cc_573 N_A_935_107#_c_542_n N_VPWR_c_1485_n 0.0124043f $X=6.03 $Y=2.555 $X2=0
+ $Y2=0
cc_574 N_A_935_107#_M1026_g N_VPWR_c_1488_n 0.00285189f $X=8.18 $Y=2.925 $X2=0
+ $Y2=0
cc_575 N_A_935_107#_c_554_n N_VPWR_c_1488_n 0.0130687f $X=8.135 $Y=3.44 $X2=0
+ $Y2=0
cc_576 N_A_935_107#_c_561_n N_VPWR_c_1488_n 0.0317254f $X=8.22 $Y=3.355 $X2=0
+ $Y2=0
cc_577 N_A_935_107#_c_562_n N_VPWR_c_1488_n 0.0622168f $X=9.625 $Y=2.66 $X2=0
+ $Y2=0
cc_578 N_A_935_107#_c_564_n N_VPWR_c_1488_n 0.0131067f $X=9.795 $Y=3.19 $X2=0
+ $Y2=0
cc_579 N_A_935_107#_M1019_g N_VPWR_c_1491_n 0.00531142f $X=12.135 $Y=3.215 $X2=0
+ $Y2=0
cc_580 N_A_935_107#_c_654_p N_VPWR_c_1491_n 0.0565954f $X=11.905 $Y=3.02 $X2=0
+ $Y2=0
cc_581 N_A_935_107#_M1008_d N_VPWR_c_1503_n 0.00479598f $X=4.79 $Y=2.845 $X2=0
+ $Y2=0
cc_582 N_A_935_107#_c_542_n N_VPWR_c_1503_n 0.0210103f $X=6.03 $Y=2.555 $X2=0
+ $Y2=0
cc_583 N_A_935_107#_M1019_g N_VPWR_c_1503_n 0.0219336f $X=12.135 $Y=3.215 $X2=0
+ $Y2=0
cc_584 N_A_935_107#_M1026_g N_VPWR_c_1503_n 0.00395199f $X=8.18 $Y=2.925 $X2=0
+ $Y2=0
cc_585 N_A_935_107#_c_551_n N_VPWR_c_1503_n 0.0117486f $X=4.93 $Y=3.13 $X2=0
+ $Y2=0
cc_586 N_A_935_107#_c_554_n N_VPWR_c_1503_n 0.0408621f $X=8.135 $Y=3.44 $X2=0
+ $Y2=0
cc_587 N_A_935_107#_c_557_n N_VPWR_c_1503_n 0.0100934f $X=7.445 $Y=3.44 $X2=0
+ $Y2=0
cc_588 N_A_935_107#_c_563_n N_VPWR_c_1503_n 0.0345138f $X=10.485 $Y=3.19 $X2=0
+ $Y2=0
cc_589 N_A_935_107#_c_564_n N_VPWR_c_1503_n 0.0097757f $X=9.795 $Y=3.19 $X2=0
+ $Y2=0
cc_590 N_A_935_107#_c_654_p N_VPWR_c_1503_n 0.0278549f $X=11.905 $Y=3.02 $X2=0
+ $Y2=0
cc_591 N_A_935_107#_c_569_n N_VPWR_c_1503_n 0.00898857f $X=10.57 $Y=3.02 $X2=0
+ $Y2=0
cc_592 N_A_935_107#_c_551_n N_A_481_107#_c_1618_n 0.0130055f $X=4.93 $Y=3.13
+ $X2=9.36 $Y2=0
cc_593 N_A_935_107#_c_551_n N_A_481_107#_c_1673_n 0.0348648f $X=4.93 $Y=3.13
+ $X2=0 $Y2=0
cc_594 N_A_935_107#_c_551_n N_A_481_107#_c_1619_n 0.0112524f $X=4.93 $Y=3.13
+ $X2=0 $Y2=0
cc_595 N_A_935_107#_c_542_n N_A_481_107#_c_1625_n 0.00465193f $X=6.03 $Y=2.555
+ $X2=0 $Y2=0
cc_596 N_A_935_107#_c_551_n N_A_481_107#_c_1625_n 0.0721322f $X=4.93 $Y=3.13
+ $X2=0 $Y2=0
cc_597 N_A_935_107#_c_542_n N_A_481_107#_c_1626_n 0.0168284f $X=6.03 $Y=2.555
+ $X2=0 $Y2=0
cc_598 N_A_935_107#_c_523_n N_A_481_107#_c_1626_n 0.0195311f $X=5.505 $Y=1.82
+ $X2=0 $Y2=0
cc_599 N_A_935_107#_M1002_g N_A_481_107#_c_1626_n 0.0230838f $X=5.755 $Y=0.825
+ $X2=0 $Y2=0
cc_600 N_A_935_107#_c_551_n N_A_481_107#_c_1627_n 0.0137873f $X=4.93 $Y=3.13
+ $X2=0 $Y2=0
cc_601 N_A_935_107#_c_523_n N_A_481_107#_c_1627_n 0.00836921f $X=5.505 $Y=1.82
+ $X2=0 $Y2=0
cc_602 N_A_935_107#_c_542_n N_A_481_107#_c_1628_n 0.0472342f $X=6.03 $Y=2.555
+ $X2=0 $Y2=0
cc_603 N_A_935_107#_c_542_n N_A_481_107#_c_1629_n 0.00673315f $X=6.03 $Y=2.555
+ $X2=0 $Y2=0
cc_604 N_A_935_107#_c_528_n N_A_481_107#_c_1635_n 0.0328735f $X=7.36 $Y=3.355
+ $X2=0 $Y2=0
cc_605 N_A_935_107#_c_542_n N_A_481_107#_c_1636_n 0.00117117f $X=6.03 $Y=2.555
+ $X2=0 $Y2=0
cc_606 N_A_935_107#_c_557_n N_A_481_107#_c_1636_n 0.0132801f $X=7.445 $Y=3.44
+ $X2=0 $Y2=0
cc_607 N_A_935_107#_c_524_n N_A_481_107#_c_1614_n 0.0209942f $X=7.06 $Y=0.35
+ $X2=0 $Y2=0
cc_608 N_A_935_107#_c_586_p N_A_481_107#_c_1614_n 0.0654149f $X=7.145 $Y=1.27
+ $X2=0 $Y2=0
cc_609 N_A_935_107#_M1002_g N_A_481_107#_c_1614_n 0.00154693f $X=5.755 $Y=0.825
+ $X2=0 $Y2=0
cc_610 N_A_935_107#_M1034_g N_A_481_107#_c_1614_n 0.00792265f $X=7.105 $Y=0.775
+ $X2=0 $Y2=0
cc_611 N_A_935_107#_c_542_n N_A_481_107#_c_1615_n 0.002045f $X=6.03 $Y=2.555
+ $X2=0 $Y2=0
cc_612 N_A_935_107#_c_528_n N_A_481_107#_c_1615_n 0.0328539f $X=7.36 $Y=3.355
+ $X2=0 $Y2=0
cc_613 N_A_935_107#_c_536_n N_A_481_107#_c_1615_n 0.0116604f $X=7.36 $Y=1.69
+ $X2=0 $Y2=0
cc_614 N_A_935_107#_M1034_g N_A_481_107#_c_1615_n 0.0207873f $X=7.105 $Y=0.775
+ $X2=0 $Y2=0
cc_615 N_A_935_107#_c_562_n A_1686_543# 0.00129068f $X=9.625 $Y=2.66 $X2=0 $Y2=0
cc_616 N_A_935_107#_c_654_p A_2335_543# 0.00488274f $X=11.905 $Y=3.02 $X2=0
+ $Y2=0
cc_617 N_A_935_107#_c_522_n N_VGND_c_1762_n 7.13035e-19 $X=4.93 $Y=1.735 $X2=0
+ $Y2=0
cc_618 N_A_935_107#_c_532_n N_VGND_c_1762_n 0.0228804f $X=4.815 $Y=0.745 $X2=0
+ $Y2=0
cc_619 N_A_935_107#_c_526_n N_VGND_c_1764_n 0.00482354f $X=5.8 $Y=0.35 $X2=0
+ $Y2=0
cc_620 N_A_935_107#_c_532_n N_VGND_c_1764_n 0.0401811f $X=4.815 $Y=0.745 $X2=0
+ $Y2=0
cc_621 N_A_935_107#_c_535_n N_VGND_c_1764_n 0.0267653f $X=5.67 $Y=1.235 $X2=0
+ $Y2=0
cc_622 N_A_935_107#_M1002_g N_VGND_c_1764_n 0.00409519f $X=5.755 $Y=0.825 $X2=0
+ $Y2=0
cc_623 N_A_935_107#_c_613_p N_VGND_c_1774_n 0.00478617f $X=5.67 $Y=1.4 $X2=0
+ $Y2=0
cc_624 N_A_935_107#_c_524_n N_VGND_c_1774_n 0.0589663f $X=7.06 $Y=0.35 $X2=0
+ $Y2=0
cc_625 N_A_935_107#_c_526_n N_VGND_c_1774_n 0.00777234f $X=5.8 $Y=0.35 $X2=0
+ $Y2=0
cc_626 N_A_935_107#_c_586_p N_VGND_c_1774_n 0.021482f $X=7.145 $Y=1.27 $X2=0
+ $Y2=0
cc_627 N_A_935_107#_c_529_n N_VGND_c_1774_n 0.0394975f $X=13.1 $Y=0.7 $X2=0
+ $Y2=0
cc_628 N_A_935_107#_c_591_p N_VGND_c_1774_n 0.0118098f $X=12.265 $Y=0.7 $X2=0
+ $Y2=0
cc_629 N_A_935_107#_c_532_n N_VGND_c_1774_n 0.0299488f $X=4.815 $Y=0.745 $X2=0
+ $Y2=0
cc_630 N_A_935_107#_c_535_n N_VGND_c_1774_n 0.0205364f $X=5.67 $Y=1.235 $X2=0
+ $Y2=0
cc_631 N_A_935_107#_M1002_g N_VGND_c_1774_n 0.0183322f $X=5.755 $Y=0.825 $X2=0
+ $Y2=0
cc_632 N_A_935_107#_M1034_g N_VGND_c_1774_n 0.0208516f $X=7.105 $Y=0.775 $X2=0
+ $Y2=0
cc_633 N_A_1201_123#_M1024_g N_A_1669_87#_c_948_n 0.0346001f $X=7.885 $Y=0.775
+ $X2=0 $Y2=0
cc_634 N_A_1201_123#_c_793_n N_A_1669_87#_c_954_n 0.105923f $X=11.97 $Y=1.96
+ $X2=0.24 $Y2=0
cc_635 N_A_1201_123#_c_793_n N_A_1669_87#_c_949_n 0.0286517f $X=11.97 $Y=1.96
+ $X2=0 $Y2=0
cc_636 N_A_1201_123#_c_806_n N_A_1669_87#_c_949_n 0.00136043f $X=8.14 $Y=1.815
+ $X2=0 $Y2=0
cc_637 N_A_1201_123#_c_799_n N_A_1669_87#_c_949_n 0.0163155f $X=7.885 $Y=1.985
+ $X2=0 $Y2=0
cc_638 N_A_1201_123#_M1024_g N_A_1669_87#_c_973_n 7.12507e-19 $X=7.885 $Y=0.775
+ $X2=0 $Y2=0
cc_639 N_A_1201_123#_c_793_n N_A_1669_87#_c_953_n 0.00151323f $X=11.97 $Y=1.96
+ $X2=0 $Y2=0
cc_640 N_A_1201_123#_c_799_n N_A_1669_87#_c_953_n 0.0386755f $X=7.885 $Y=1.985
+ $X2=0 $Y2=0
cc_641 N_A_1201_123#_c_793_n N_A_1471_113#_M1016_g 0.0315195f $X=11.97 $Y=1.96
+ $X2=0 $Y2=0
cc_642 N_A_1201_123#_c_798_n N_A_1471_113#_M1016_g 0.00425102f $X=12.135 $Y=1.85
+ $X2=0 $Y2=0
cc_643 N_A_1201_123#_M1013_g N_A_1471_113#_M1011_g 0.0530536f $X=12.22 $Y=0.91
+ $X2=18.48 $Y2=0
cc_644 N_A_1201_123#_c_793_n N_A_1471_113#_c_1013_n 8.78178e-19 $X=11.97 $Y=1.96
+ $X2=0 $Y2=0
cc_645 N_A_1201_123#_M1024_g N_A_1471_113#_c_1014_n 0.00418657f $X=7.885
+ $Y=0.775 $X2=0 $Y2=0
cc_646 N_A_1201_123#_c_799_n N_A_1471_113#_c_1014_n 0.0107611f $X=7.885 $Y=1.985
+ $X2=0 $Y2=0
cc_647 N_A_1201_123#_M1004_g N_A_1471_113#_c_1026_n 0.00341076f $X=7.4 $Y=2.925
+ $X2=0 $Y2=0
cc_648 N_A_1201_123#_c_799_n N_A_1471_113#_c_1026_n 0.00482128f $X=7.885
+ $Y=1.985 $X2=0 $Y2=0
cc_649 N_A_1201_123#_M1004_g N_A_1471_113#_c_1027_n 0.00641061f $X=7.4 $Y=2.925
+ $X2=0 $Y2=0
cc_650 N_A_1201_123#_c_793_n N_A_1471_113#_c_1015_n 0.00814632f $X=11.97 $Y=1.96
+ $X2=0 $Y2=0
cc_651 N_A_1201_123#_c_806_n N_A_1471_113#_c_1015_n 0.023175f $X=8.14 $Y=1.815
+ $X2=0 $Y2=0
cc_652 N_A_1201_123#_c_799_n N_A_1471_113#_c_1015_n 0.0372255f $X=7.885 $Y=1.985
+ $X2=0 $Y2=0
cc_653 N_A_1201_123#_M1013_g N_A_1471_113#_c_1016_n 7.40292e-19 $X=12.22 $Y=0.91
+ $X2=0 $Y2=0
cc_654 N_A_1201_123#_c_807_n N_A_1471_113#_c_1016_n 3.2208e-19 $X=12.135 $Y=1.85
+ $X2=0 $Y2=0
cc_655 N_A_1201_123#_c_793_n N_A_1471_113#_c_1017_n 0.0176918f $X=11.97 $Y=1.96
+ $X2=0 $Y2=0
cc_656 N_A_1201_123#_c_807_n N_A_1471_113#_c_1017_n 0.00143681f $X=12.135
+ $Y=1.85 $X2=0 $Y2=0
cc_657 N_A_1201_123#_c_798_n N_A_1471_113#_c_1017_n 0.0530536f $X=12.135 $Y=1.85
+ $X2=0 $Y2=0
cc_658 N_A_1201_123#_M1024_g N_A_1471_113#_c_1018_n 0.0188375f $X=7.885 $Y=0.775
+ $X2=0 $Y2=0
cc_659 N_A_1201_123#_c_799_n N_A_1471_113#_c_1018_n 0.00289451f $X=7.885
+ $Y=1.985 $X2=0 $Y2=0
cc_660 N_A_1201_123#_c_799_n N_A_1471_113#_c_1050_n 0.00452645f $X=7.885
+ $Y=1.985 $X2=0 $Y2=0
cc_661 N_A_1201_123#_M1004_g N_A_1471_113#_c_1029_n 0.00207946f $X=7.4 $Y=2.925
+ $X2=0 $Y2=0
cc_662 N_A_1201_123#_c_806_n N_A_1471_113#_c_1029_n 0.023378f $X=8.14 $Y=1.815
+ $X2=0 $Y2=0
cc_663 N_A_1201_123#_c_799_n N_A_1471_113#_c_1029_n 0.0511806f $X=7.885 $Y=1.985
+ $X2=0 $Y2=0
cc_664 N_A_1201_123#_c_793_n N_A_1471_113#_c_1020_n 0.0127692f $X=11.97 $Y=1.96
+ $X2=0 $Y2=0
cc_665 N_A_1201_123#_c_799_n N_A_1471_113#_c_1020_n 0.00369781f $X=7.885
+ $Y=1.985 $X2=0 $Y2=0
cc_666 N_A_1201_123#_c_793_n N_A_1471_113#_c_1021_n 0.0269928f $X=11.97 $Y=1.96
+ $X2=0 $Y2=0
cc_667 N_A_1201_123#_c_793_n N_A_1471_113#_c_1022_n 0.194179f $X=11.97 $Y=1.96
+ $X2=0 $Y2=0
cc_668 N_A_1201_123#_c_793_n N_SET_B_c_1156_n 0.00449676f $X=11.97 $Y=1.96 $X2=0
+ $Y2=0
cc_669 N_A_1201_123#_M1013_g N_SET_B_c_1146_n 5.64047e-19 $X=12.22 $Y=0.91 $X2=0
+ $Y2=0
cc_670 N_A_1201_123#_c_793_n N_SET_B_c_1146_n 0.00329288f $X=11.97 $Y=1.96 $X2=0
+ $Y2=0
cc_671 N_A_1201_123#_M1013_g N_SET_B_c_1165_n 0.00334078f $X=12.22 $Y=0.91 $X2=0
+ $Y2=0
cc_672 N_A_1201_123#_M1013_g N_SET_B_c_1147_n 0.0169208f $X=12.22 $Y=0.91 $X2=0
+ $Y2=0
cc_673 N_A_1201_123#_c_793_n N_SET_B_M1010_g 0.04147f $X=11.97 $Y=1.96 $X2=0
+ $Y2=0
cc_674 N_A_1201_123#_c_798_n N_A_2698_421#_c_1237_n 9.71813e-19 $X=12.135
+ $Y=1.85 $X2=0 $Y2=0
cc_675 N_A_1201_123#_c_798_n N_A_2698_421#_c_1238_n 0.0410273f $X=12.135 $Y=1.85
+ $X2=18.48 $Y2=0
cc_676 N_A_1201_123#_c_801_n N_A_2698_421#_c_1248_n 0.0410273f $X=13.03 $Y=2.605
+ $X2=0 $Y2=0
cc_677 N_A_1201_123#_c_801_n N_A_2477_543#_c_1318_n 0.00651293f $X=13.03
+ $Y=2.605 $X2=0 $Y2=0
cc_678 N_A_1201_123#_M1013_g N_A_2477_543#_c_1332_n 0.00379626f $X=12.22 $Y=0.91
+ $X2=0 $Y2=0
cc_679 N_A_1201_123#_c_798_n N_A_2477_543#_c_1332_n 0.00451279f $X=12.135
+ $Y=1.85 $X2=0 $Y2=0
cc_680 N_A_1201_123#_M1013_g N_A_2477_543#_c_1310_n 0.00252612f $X=12.22 $Y=0.91
+ $X2=0 $Y2=0
cc_681 N_A_1201_123#_c_798_n N_A_2477_543#_c_1310_n 0.00445246f $X=12.135
+ $Y=1.85 $X2=0 $Y2=0
cc_682 N_A_1201_123#_c_801_n N_A_2477_543#_c_1322_n 0.00345749f $X=13.03
+ $Y=2.605 $X2=0 $Y2=0
cc_683 N_A_1201_123#_c_798_n N_A_2477_543#_c_1322_n 0.0233112f $X=12.135 $Y=1.85
+ $X2=0 $Y2=0
cc_684 N_A_1201_123#_c_801_n N_A_2477_543#_c_1325_n 0.0117449f $X=13.03 $Y=2.605
+ $X2=0 $Y2=0
cc_685 N_A_1201_123#_c_798_n N_A_2477_543#_c_1325_n 0.00869441f $X=12.135
+ $Y=1.85 $X2=0 $Y2=0
cc_686 N_A_1201_123#_c_798_n N_A_2477_543#_c_1350_n 0.0100538f $X=12.135 $Y=1.85
+ $X2=0 $Y2=0
cc_687 N_A_1201_123#_c_798_n N_A_2477_543#_c_1326_n 0.0183868f $X=12.135 $Y=1.85
+ $X2=0 $Y2=0
cc_688 N_A_1201_123#_c_801_n N_VPWR_c_1494_n 0.02054f $X=13.03 $Y=2.605 $X2=0
+ $Y2=0
cc_689 N_A_1201_123#_M1004_g N_VPWR_c_1503_n 0.00395199f $X=7.4 $Y=2.925 $X2=0
+ $Y2=0
cc_690 N_A_1201_123#_c_801_n N_VPWR_c_1503_n 0.015231f $X=13.03 $Y=2.605 $X2=0
+ $Y2=0
cc_691 N_A_1201_123#_c_802_n N_VPWR_c_1503_n 0.0191099f $X=6.42 $Y=2.79 $X2=0
+ $Y2=0
cc_692 N_A_1201_123#_c_802_n N_A_481_107#_c_1626_n 0.0137367f $X=6.42 $Y=2.79
+ $X2=0 $Y2=0
cc_693 N_A_1201_123#_c_799_n N_A_481_107#_c_1626_n 3.35965e-19 $X=7.885 $Y=1.985
+ $X2=0 $Y2=0
cc_694 N_A_1201_123#_c_802_n N_A_481_107#_c_1628_n 0.0677365f $X=6.42 $Y=2.79
+ $X2=0 $Y2=0
cc_695 N_A_1201_123#_c_802_n N_A_481_107#_c_1629_n 0.0186039f $X=6.42 $Y=2.79
+ $X2=0 $Y2=0
cc_696 N_A_1201_123#_M1004_g N_A_481_107#_c_1635_n 0.0056354f $X=7.4 $Y=2.925
+ $X2=0 $Y2=0
cc_697 N_A_1201_123#_c_792_n N_A_481_107#_c_1635_n 0.0496454f $X=6.335 $Y=1.9
+ $X2=0 $Y2=0
cc_698 N_A_1201_123#_c_799_n N_A_481_107#_c_1635_n 0.0110659f $X=7.885 $Y=1.985
+ $X2=0 $Y2=0
cc_699 N_A_1201_123#_c_805_n N_A_481_107#_c_1636_n 0.0496454f $X=6.335 $Y=2.095
+ $X2=0 $Y2=0
cc_700 N_A_1201_123#_c_794_n N_A_481_107#_c_1614_n 0.0229129f $X=6.145 $Y=0.825
+ $X2=0 $Y2=0
cc_701 N_A_1201_123#_c_796_n N_A_481_107#_c_1614_n 0.00342053f $X=6.4 $Y=1.59
+ $X2=0 $Y2=0
cc_702 N_A_1201_123#_M1004_g N_A_481_107#_c_1615_n 0.00212133f $X=7.4 $Y=2.925
+ $X2=0 $Y2=0
cc_703 N_A_1201_123#_c_794_n N_A_481_107#_c_1615_n 0.0166048f $X=6.145 $Y=0.825
+ $X2=0 $Y2=0
cc_704 N_A_1201_123#_c_795_n N_A_481_107#_c_1615_n 0.0496454f $X=6.4 $Y=1.59
+ $X2=0 $Y2=0
cc_705 N_A_1201_123#_c_796_n N_A_481_107#_c_1615_n 0.00825389f $X=6.4 $Y=1.59
+ $X2=0 $Y2=0
cc_706 N_A_1201_123#_c_799_n N_A_481_107#_c_1615_n 0.0383529f $X=7.885 $Y=1.985
+ $X2=0 $Y2=0
cc_707 N_A_1201_123#_M1024_g N_VGND_c_1766_n 0.00665476f $X=7.885 $Y=0.775 $X2=0
+ $Y2=0
cc_708 N_A_1201_123#_M1002_d N_VGND_c_1774_n 0.00212289f $X=6.005 $Y=0.615 $X2=0
+ $Y2=0
cc_709 N_A_1201_123#_M1024_g N_VGND_c_1774_n 0.024072f $X=7.885 $Y=0.775 $X2=0
+ $Y2=0
cc_710 N_A_1201_123#_M1013_g N_VGND_c_1774_n 0.00964903f $X=12.22 $Y=0.91 $X2=0
+ $Y2=0
cc_711 N_A_1201_123#_c_794_n N_VGND_c_1774_n 0.0119459f $X=6.145 $Y=0.825 $X2=0
+ $Y2=0
cc_712 N_A_1669_87#_c_951_n N_A_1471_113#_c_1011_n 0.0168529f $X=9.535 $Y=0.745
+ $X2=0 $Y2=0
cc_713 N_A_1669_87#_c_948_n N_A_1471_113#_c_1013_n 3.8924e-19 $X=8.595 $Y=1.095
+ $X2=0 $Y2=0
cc_714 N_A_1669_87#_c_950_n N_A_1471_113#_c_1013_n 0.0125385f $X=9.37 $Y=1.19
+ $X2=0 $Y2=0
cc_715 N_A_1669_87#_c_951_n N_A_1471_113#_c_1013_n 0.00606452f $X=9.535 $Y=0.745
+ $X2=0 $Y2=0
cc_716 N_A_1669_87#_c_973_n N_A_1471_113#_c_1013_n 4.82138e-19 $X=9.165 $Y=1.225
+ $X2=0 $Y2=0
cc_717 N_A_1669_87#_c_953_n N_A_1471_113#_c_1013_n 0.0230596f $X=8.89 $Y=1.595
+ $X2=0 $Y2=0
cc_718 N_A_1669_87#_c_948_n N_A_1471_113#_c_1014_n 0.00129468f $X=8.595 $Y=1.095
+ $X2=0 $Y2=0
cc_719 N_A_1669_87#_c_953_n N_A_1471_113#_c_1015_n 0.00728824f $X=8.89 $Y=1.595
+ $X2=0 $Y2=0
cc_720 N_A_1669_87#_c_948_n N_A_1471_113#_c_1018_n 7.02965e-19 $X=8.595 $Y=1.095
+ $X2=0 $Y2=0
cc_721 N_A_1669_87#_c_949_n N_A_1471_113#_c_1020_n 0.00158116f $X=8.955 $Y=2.31
+ $X2=0 $Y2=0
cc_722 N_A_1669_87#_c_953_n N_A_1471_113#_c_1020_n 0.0178853f $X=8.89 $Y=1.595
+ $X2=0 $Y2=0
cc_723 N_A_1669_87#_c_954_n N_A_1471_113#_c_1021_n 0.0314637f $X=9.975 $Y=2.31
+ $X2=0 $Y2=0
cc_724 N_A_1669_87#_c_949_n N_A_1471_113#_c_1021_n 0.0589016f $X=8.955 $Y=2.31
+ $X2=0 $Y2=0
cc_725 N_A_1669_87#_c_965_n N_A_1471_113#_c_1021_n 0.0183589f $X=10.14 $Y=2.84
+ $X2=0 $Y2=0
cc_726 N_A_1669_87#_c_949_n N_A_1471_113#_c_1022_n 0.0130275f $X=8.955 $Y=2.31
+ $X2=0 $Y2=0
cc_727 N_A_1669_87#_c_950_n N_A_1471_113#_c_1022_n 0.021065f $X=9.37 $Y=1.19
+ $X2=0 $Y2=0
cc_728 N_A_1669_87#_c_973_n N_A_1471_113#_c_1022_n 0.0219469f $X=9.165 $Y=1.225
+ $X2=0 $Y2=0
cc_729 N_A_1669_87#_c_953_n N_A_1471_113#_c_1022_n 0.0151908f $X=8.89 $Y=1.595
+ $X2=0 $Y2=0
cc_730 N_A_1669_87#_c_950_n N_A_1471_113#_c_1110_n 0.013372f $X=9.37 $Y=1.19
+ $X2=0 $Y2=0
cc_731 N_A_1669_87#_c_953_n N_A_1471_113#_c_1110_n 4.69503e-19 $X=8.89 $Y=1.595
+ $X2=0 $Y2=0
cc_732 N_A_1669_87#_c_954_n N_SET_B_c_1156_n 0.0110317f $X=9.975 $Y=2.31 $X2=0
+ $Y2=0
cc_733 N_A_1669_87#_c_965_n N_SET_B_c_1156_n 0.0291022f $X=10.14 $Y=2.84 $X2=0
+ $Y2=0
cc_734 N_A_1669_87#_c_950_n N_SET_B_M1010_g 5.139e-19 $X=9.37 $Y=1.19 $X2=0
+ $Y2=0
cc_735 N_A_1669_87#_c_951_n N_SET_B_M1010_g 7.1237e-19 $X=9.535 $Y=0.745 $X2=0
+ $Y2=0
cc_736 N_A_1669_87#_c_949_n N_VPWR_c_1488_n 0.0378426f $X=8.955 $Y=2.31 $X2=0
+ $Y2=0
cc_737 N_A_1669_87#_c_948_n N_VGND_c_1766_n 0.0491045f $X=8.595 $Y=1.095 $X2=0
+ $Y2=0
cc_738 N_A_1669_87#_c_951_n N_VGND_c_1766_n 0.0283112f $X=9.535 $Y=0.745 $X2=0
+ $Y2=0
cc_739 N_A_1669_87#_c_973_n N_VGND_c_1766_n 0.0205415f $X=9.165 $Y=1.225 $X2=0
+ $Y2=0
cc_740 N_A_1669_87#_c_953_n N_VGND_c_1766_n 0.00810568f $X=8.89 $Y=1.595 $X2=0
+ $Y2=0
cc_741 N_A_1669_87#_c_951_n N_VGND_c_1768_n 0.00640403f $X=9.535 $Y=0.745 $X2=0
+ $Y2=0
cc_742 N_A_1669_87#_c_951_n N_VGND_c_1774_n 0.0272756f $X=9.535 $Y=0.745 $X2=0
+ $Y2=0
cc_743 N_A_1669_87#_c_973_n N_VGND_c_1774_n 0.00921454f $X=9.165 $Y=1.225 $X2=0
+ $Y2=0
cc_744 N_A_1669_87#_c_953_n N_VGND_c_1774_n 8.70972e-19 $X=8.89 $Y=1.595 $X2=0
+ $Y2=0
cc_745 N_A_1471_113#_M1016_g N_SET_B_c_1156_n 0.0585711f $X=11.425 $Y=3.215
+ $X2=0 $Y2=0
cc_746 N_A_1471_113#_c_1021_n N_SET_B_c_1156_n 0.040587f $X=9.685 $Y=1.575 $X2=0
+ $Y2=0
cc_747 N_A_1471_113#_M1011_g N_SET_B_c_1146_n 0.0220387f $X=11.51 $Y=0.91 $X2=0
+ $Y2=0
cc_748 N_A_1471_113#_c_1013_n N_SET_B_c_1146_n 9.16753e-19 $X=9.837 $Y=1.565
+ $X2=0 $Y2=0
cc_749 N_A_1471_113#_c_1016_n N_SET_B_c_1146_n 0.0670632f $X=11.36 $Y=1.61 $X2=0
+ $Y2=0
cc_750 N_A_1471_113#_c_1017_n N_SET_B_c_1146_n 0.00253167f $X=11.36 $Y=1.61
+ $X2=0 $Y2=0
cc_751 N_A_1471_113#_M1011_g N_SET_B_c_1165_n 0.0324908f $X=11.51 $Y=0.91 $X2=0
+ $Y2=0
cc_752 N_A_1471_113#_M1011_g N_SET_B_c_1147_n 0.00570881f $X=11.51 $Y=0.91 $X2=0
+ $Y2=0
cc_753 N_A_1471_113#_M1011_g N_SET_B_c_1149_n 0.00363307f $X=11.51 $Y=0.91 $X2=0
+ $Y2=0
cc_754 N_A_1471_113#_M1011_g N_SET_B_M1010_g 0.0281191f $X=11.51 $Y=0.91 $X2=0
+ $Y2=0
cc_755 N_A_1471_113#_c_1011_n N_SET_B_M1010_g 0.082526f $X=9.837 $Y=1.065 $X2=0
+ $Y2=0
cc_756 N_A_1471_113#_c_1016_n N_SET_B_M1010_g 0.0280953f $X=11.36 $Y=1.61 $X2=0
+ $Y2=0
cc_757 N_A_1471_113#_c_1017_n N_SET_B_M1010_g 0.0328325f $X=11.36 $Y=1.61 $X2=0
+ $Y2=0
cc_758 N_A_1471_113#_c_1021_n N_SET_B_M1010_g 0.0198672f $X=9.685 $Y=1.575 $X2=0
+ $Y2=0
cc_759 N_A_1471_113#_c_1110_n N_SET_B_M1010_g 2.68614e-19 $X=9.85 $Y=1.575 $X2=0
+ $Y2=0
cc_760 N_A_1471_113#_M1016_g N_A_2477_543#_c_1318_n 0.00108343f $X=11.425
+ $Y=3.215 $X2=0 $Y2=0
cc_761 N_A_1471_113#_c_1021_n N_VPWR_c_1488_n 0.00286454f $X=9.685 $Y=1.575
+ $X2=0 $Y2=0
cc_762 N_A_1471_113#_M1016_g N_VPWR_c_1491_n 0.0354328f $X=11.425 $Y=3.215 $X2=0
+ $Y2=0
cc_763 N_A_1471_113#_M1016_g N_VPWR_c_1503_n 0.00250239f $X=11.425 $Y=3.215
+ $X2=0 $Y2=0
cc_764 N_A_1471_113#_c_1027_n N_VPWR_c_1503_n 0.00214844f $X=7.79 $Y=2.925 $X2=0
+ $Y2=0
cc_765 N_A_1471_113#_c_1021_n N_VPWR_c_1503_n 0.00393471f $X=9.685 $Y=1.575
+ $X2=0 $Y2=0
cc_766 N_A_1471_113#_c_1011_n N_VGND_c_1766_n 0.00267849f $X=9.837 $Y=1.065
+ $X2=0 $Y2=0
cc_767 N_A_1471_113#_c_1015_n N_VGND_c_1766_n 0.00973359f $X=8.485 $Y=1.44 $X2=0
+ $Y2=0
cc_768 N_A_1471_113#_c_1018_n N_VGND_c_1766_n 0.0153246f $X=7.71 $Y=0.775 $X2=0
+ $Y2=0
cc_769 N_A_1471_113#_c_1020_n N_VGND_c_1766_n 0.00623408f $X=8.57 $Y=1.44 $X2=0
+ $Y2=0
cc_770 N_A_1471_113#_c_1022_n N_VGND_c_1766_n 0.00473013f $X=9.52 $Y=1.575 $X2=0
+ $Y2=0
cc_771 N_A_1471_113#_M1011_g N_VGND_c_1768_n 0.0121444f $X=11.51 $Y=0.91 $X2=0
+ $Y2=0
cc_772 N_A_1471_113#_c_1011_n N_VGND_c_1768_n 0.00444483f $X=9.837 $Y=1.065
+ $X2=0 $Y2=0
cc_773 N_A_1471_113#_c_1016_n N_VGND_c_1768_n 0.00632721f $X=11.36 $Y=1.61 $X2=0
+ $Y2=0
cc_774 N_A_1471_113#_M1034_d N_VGND_c_1774_n 0.00221032f $X=7.355 $Y=0.565 $X2=0
+ $Y2=0
cc_775 N_A_1471_113#_M1011_g N_VGND_c_1774_n 0.0114155f $X=11.51 $Y=0.91 $X2=0
+ $Y2=0
cc_776 N_A_1471_113#_c_1011_n N_VGND_c_1774_n 0.033371f $X=9.837 $Y=1.065 $X2=0
+ $Y2=0
cc_777 N_A_1471_113#_c_1014_n N_VGND_c_1774_n 4.27235e-19 $X=7.71 $Y=1.355 $X2=0
+ $Y2=0
cc_778 N_A_1471_113#_c_1018_n N_VGND_c_1774_n 0.0260656f $X=7.71 $Y=0.775 $X2=0
+ $Y2=0
cc_779 N_SET_B_c_1147_n N_A_2698_421#_M1014_g 0.0154529f $X=14.045 $Y=0.35 $X2=0
+ $Y2=0
cc_780 SET_B N_A_2698_421#_M1014_g 0.0135543f $X=14.075 $Y=0.84 $X2=0 $Y2=0
cc_781 SET_B N_A_2698_421#_M1014_g 0.0323398f $X=14.075 $Y=1.21 $X2=0 $Y2=0
cc_782 N_SET_B_M1015_g N_A_2698_421#_M1014_g 0.127564f $X=14.52 $Y=1.075 $X2=0
+ $Y2=0
cc_783 N_SET_B_c_1155_n N_A_2698_421#_M1014_g 0.00391751f $X=14.282 $Y=0.81
+ $X2=0 $Y2=0
cc_784 N_SET_B_M1015_g N_A_2698_421#_c_1237_n 0.0204714f $X=14.52 $Y=1.075 $X2=0
+ $Y2=0
cc_785 N_SET_B_M1015_g N_A_2698_421#_c_1239_n 0.036352f $X=14.52 $Y=1.075 $X2=0
+ $Y2=0
cc_786 N_SET_B_M1015_g N_A_2698_421#_c_1240_n 0.0090724f $X=14.52 $Y=1.075
+ $X2=9.36 $Y2=0
cc_787 N_SET_B_M1015_g N_A_2698_421#_c_1246_n 0.00378698f $X=14.52 $Y=1.075
+ $X2=0 $Y2=0
cc_788 N_SET_B_M1015_g N_A_2698_421#_c_1247_n 4.13202e-19 $X=14.52 $Y=1.075
+ $X2=0 $Y2=0
cc_789 N_SET_B_M1015_g N_A_2698_421#_c_1248_n 0.0125575f $X=14.52 $Y=1.075 $X2=0
+ $Y2=0
cc_790 SET_B N_A_2477_543#_M1023_g 2.51573e-19 $X=14.075 $Y=0.84 $X2=0 $Y2=0
cc_791 SET_B N_A_2477_543#_M1023_g 0.00195922f $X=14.075 $Y=1.21 $X2=0 $Y2=0
cc_792 N_SET_B_M1015_g N_A_2477_543#_M1023_g 0.0354509f $X=14.52 $Y=1.075 $X2=0
+ $Y2=0
cc_793 N_SET_B_M1015_g N_A_2477_543#_c_1323_n 0.0291748f $X=14.52 $Y=1.075 $X2=0
+ $Y2=0
cc_794 N_SET_B_M1015_g N_A_2477_543#_c_1324_n 0.00675269f $X=14.52 $Y=1.075
+ $X2=0 $Y2=0
cc_795 N_SET_B_M1015_g N_A_2477_543#_c_1370_n 0.00264961f $X=14.52 $Y=1.075
+ $X2=0 $Y2=0
cc_796 SET_B N_A_2477_543#_c_1326_n 0.0361634f $X=14.075 $Y=1.21 $X2=0 $Y2=0
cc_797 N_SET_B_M1015_g N_A_2477_543#_c_1326_n 0.0338381f $X=14.52 $Y=1.075 $X2=0
+ $Y2=0
cc_798 N_SET_B_M1015_g N_VPWR_c_1494_n 0.00179323f $X=14.52 $Y=1.075 $X2=0 $Y2=0
cc_799 N_SET_B_c_1156_n N_VPWR_c_1503_n 0.00398012f $X=10.582 $Y=2.605 $X2=0
+ $Y2=0
cc_800 N_SET_B_M1015_g N_VPWR_c_1503_n 0.00395199f $X=14.52 $Y=1.075 $X2=0 $Y2=0
cc_801 N_SET_B_c_1146_n N_VGND_M1010_d 0.00231484f $X=11.465 $Y=1.26 $X2=-0.33
+ $Y2=-0.265
cc_802 N_SET_B_c_1146_n N_VGND_c_1768_n 0.0504223f $X=11.465 $Y=1.26 $X2=0 $Y2=0
cc_803 N_SET_B_c_1165_n N_VGND_c_1768_n 0.0384016f $X=11.55 $Y=1.175 $X2=0 $Y2=0
cc_804 N_SET_B_c_1149_n N_VGND_c_1768_n 0.00465917f $X=11.635 $Y=0.35 $X2=0
+ $Y2=0
cc_805 N_SET_B_M1010_g N_VGND_c_1768_n 0.0548894f $X=10.635 $Y=0.745 $X2=0 $Y2=0
cc_806 N_SET_B_c_1147_n N_VGND_c_1770_n 0.00170665f $X=14.045 $Y=0.35 $X2=0
+ $Y2=0
cc_807 SET_B N_VGND_c_1770_n 0.0401019f $X=14.075 $Y=0.84 $X2=0 $Y2=0
cc_808 N_SET_B_M1015_g N_VGND_c_1770_n 0.0196486f $X=14.52 $Y=1.075 $X2=0 $Y2=0
cc_809 N_SET_B_c_1155_n N_VGND_c_1770_n 0.011667f $X=14.282 $Y=0.81 $X2=0 $Y2=0
cc_810 N_SET_B_c_1146_n N_VGND_c_1774_n 0.00754612f $X=11.465 $Y=1.26 $X2=0
+ $Y2=0
cc_811 N_SET_B_c_1165_n N_VGND_c_1774_n 0.0200609f $X=11.55 $Y=1.175 $X2=0 $Y2=0
cc_812 N_SET_B_c_1147_n N_VGND_c_1774_n 0.100677f $X=14.045 $Y=0.35 $X2=0 $Y2=0
cc_813 N_SET_B_c_1149_n N_VGND_c_1774_n 0.00774482f $X=11.635 $Y=0.35 $X2=0
+ $Y2=0
cc_814 SET_B N_VGND_c_1774_n 0.0161527f $X=14.075 $Y=0.84 $X2=0 $Y2=0
cc_815 N_SET_B_M1015_g N_VGND_c_1774_n 0.0140782f $X=14.52 $Y=1.075 $X2=0 $Y2=0
cc_816 N_SET_B_c_1155_n N_VGND_c_1774_n 0.0233663f $X=14.282 $Y=0.81 $X2=0 $Y2=0
cc_817 N_A_2698_421#_c_1235_n N_A_2477_543#_M1023_g 0.00719969f $X=15.855
+ $Y=1.075 $X2=0 $Y2=0
cc_818 N_A_2698_421#_c_1240_n N_A_2477_543#_M1020_g 0.00368185f $X=15.295
+ $Y=3.42 $X2=18.48 $Y2=0
cc_819 N_A_2698_421#_c_1246_n N_A_2477_543#_M1020_g 0.0178282f $X=15.46 $Y=3.275
+ $X2=18.48 $Y2=0
cc_820 N_A_2698_421#_c_1247_n N_A_2477_543#_M1020_g 0.0286759f $X=15.895
+ $Y=2.695 $X2=18.48 $Y2=0
cc_821 N_A_2698_421#_c_1235_n N_A_2477_543#_M1020_g 0.0410475f $X=15.855
+ $Y=1.075 $X2=18.48 $Y2=0
cc_822 N_A_2698_421#_M1014_g N_A_2477_543#_c_1310_n 0.00130453f $X=13.81
+ $Y=1.075 $X2=0 $Y2=0
cc_823 N_A_2698_421#_c_1238_n N_A_2477_543#_c_1322_n 0.00210957f $X=13.875
+ $Y=2.39 $X2=0 $Y2=0
cc_824 N_A_2698_421#_c_1237_n N_A_2477_543#_c_1323_n 0.0156266f $X=14.395
+ $Y=2.392 $X2=0 $Y2=0
cc_825 N_A_2698_421#_c_1238_n N_A_2477_543#_c_1323_n 4.41792e-19 $X=13.875
+ $Y=2.39 $X2=0 $Y2=0
cc_826 N_A_2698_421#_c_1239_n N_A_2477_543#_c_1323_n 0.0449883f $X=14.48
+ $Y=3.335 $X2=0 $Y2=0
cc_827 N_A_2698_421#_c_1240_n N_A_2477_543#_c_1323_n 0.0242156f $X=15.295
+ $Y=3.42 $X2=0 $Y2=0
cc_828 N_A_2698_421#_c_1246_n N_A_2477_543#_c_1323_n 0.0201625f $X=15.46
+ $Y=3.275 $X2=0 $Y2=0
cc_829 N_A_2698_421#_c_1247_n N_A_2477_543#_c_1323_n 0.012396f $X=15.895
+ $Y=2.695 $X2=0 $Y2=0
cc_830 N_A_2698_421#_c_1247_n N_A_2477_543#_c_1324_n 0.00917033f $X=15.895
+ $Y=2.695 $X2=0 $Y2=0
cc_831 N_A_2698_421#_c_1235_n N_A_2477_543#_c_1324_n 0.0170317f $X=15.855
+ $Y=1.075 $X2=0 $Y2=0
cc_832 N_A_2698_421#_c_1235_n N_A_2477_543#_c_1370_n 0.0298701f $X=15.855
+ $Y=1.075 $X2=0 $Y2=0
cc_833 N_A_2698_421#_M1014_g N_A_2477_543#_c_1326_n 0.0349115f $X=13.81 $Y=1.075
+ $X2=0 $Y2=0
cc_834 N_A_2698_421#_c_1237_n N_A_2477_543#_c_1326_n 0.0589434f $X=14.395
+ $Y=2.392 $X2=0 $Y2=0
cc_835 N_A_2698_421#_c_1238_n N_A_2477_543#_c_1326_n 0.0121971f $X=13.875
+ $Y=2.39 $X2=0 $Y2=0
cc_836 N_A_2698_421#_c_1247_n N_A_2477_543#_c_1311_n 0.00634828f $X=15.895
+ $Y=2.695 $X2=0 $Y2=0
cc_837 N_A_2698_421#_c_1235_n N_A_2477_543#_c_1311_n 0.0559653f $X=15.855
+ $Y=1.075 $X2=0 $Y2=0
cc_838 N_A_2698_421#_c_1235_n N_A_3321_173#_c_1432_n 0.0233603f $X=15.855
+ $Y=1.075 $X2=18.48 $Y2=0
cc_839 N_A_2698_421#_c_1235_n N_A_3321_173#_c_1442_n 0.00493656f $X=15.855
+ $Y=1.075 $X2=0 $Y2=0
cc_840 N_A_2698_421#_c_1247_n N_A_3321_173#_c_1438_n 0.00571777f $X=15.895
+ $Y=2.695 $X2=0 $Y2=0
cc_841 N_A_2698_421#_c_1235_n N_A_3321_173#_c_1439_n 0.031139f $X=15.855
+ $Y=1.075 $X2=0 $Y2=0
cc_842 N_A_2698_421#_c_1237_n N_VPWR_c_1494_n 0.0387617f $X=14.395 $Y=2.392
+ $X2=0 $Y2=0
cc_843 N_A_2698_421#_c_1238_n N_VPWR_c_1494_n 0.00216433f $X=13.875 $Y=2.39
+ $X2=0 $Y2=0
cc_844 N_A_2698_421#_c_1239_n N_VPWR_c_1494_n 0.0322093f $X=14.48 $Y=3.335 $X2=0
+ $Y2=0
cc_845 N_A_2698_421#_c_1243_n N_VPWR_c_1494_n 0.0140554f $X=14.565 $Y=3.42 $X2=0
+ $Y2=0
cc_846 N_A_2698_421#_c_1248_n N_VPWR_c_1494_n 0.0562761f $X=13.775 $Y=2.605
+ $X2=0 $Y2=0
cc_847 N_A_2698_421#_c_1240_n N_VPWR_c_1497_n 0.0118797f $X=15.295 $Y=3.42 $X2=0
+ $Y2=0
cc_848 N_A_2698_421#_c_1246_n N_VPWR_c_1497_n 0.020798f $X=15.46 $Y=3.275 $X2=0
+ $Y2=0
cc_849 N_A_2698_421#_c_1247_n N_VPWR_c_1497_n 0.0143675f $X=15.895 $Y=2.695
+ $X2=0 $Y2=0
cc_850 N_A_2698_421#_c_1240_n N_VPWR_c_1503_n 0.0535002f $X=15.295 $Y=3.42 $X2=0
+ $Y2=0
cc_851 N_A_2698_421#_c_1243_n N_VPWR_c_1503_n 0.00966809f $X=14.565 $Y=3.42
+ $X2=0 $Y2=0
cc_852 N_A_2698_421#_c_1247_n N_VPWR_c_1503_n 0.00641323f $X=15.895 $Y=2.695
+ $X2=0 $Y2=0
cc_853 N_A_2698_421#_M1014_g N_VGND_c_1770_n 2.31738e-19 $X=13.81 $Y=1.075 $X2=0
+ $Y2=0
cc_854 N_A_2698_421#_c_1235_n N_VGND_c_1770_n 0.0230119f $X=15.855 $Y=1.075
+ $X2=0 $Y2=0
cc_855 N_A_2698_421#_M1014_g N_VGND_c_1774_n 0.0158747f $X=13.81 $Y=1.075 $X2=0
+ $Y2=0
cc_856 N_A_2698_421#_c_1235_n N_VGND_c_1774_n 0.0137969f $X=15.855 $Y=1.075
+ $X2=0 $Y2=0
cc_857 N_A_2477_543#_M1032_g N_A_3321_173#_M1003_g 0.0145305f $X=17.14 $Y=1.075
+ $X2=0 $Y2=0
cc_858 N_A_2477_543#_M1033_g N_A_3321_173#_M1035_g 0.0192904f $X=17.18 $Y=2.75
+ $X2=0 $Y2=0
cc_859 N_A_2477_543#_c_1307_n N_A_3321_173#_c_1432_n 0.00993214f $X=16.89
+ $Y=1.665 $X2=18.48 $Y2=0
cc_860 N_A_2477_543#_M1032_g N_A_3321_173#_c_1432_n 0.01694f $X=17.14 $Y=1.075
+ $X2=18.48 $Y2=0
cc_861 N_A_2477_543#_c_1309_n N_A_3321_173#_c_1432_n 0.00421489f $X=17.16
+ $Y=1.665 $X2=18.48 $Y2=0
cc_862 N_A_2477_543#_c_1309_n N_A_3321_173#_c_1433_n 0.0453981f $X=17.16
+ $Y=1.665 $X2=9.36 $Y2=0.057
cc_863 N_A_2477_543#_c_1307_n N_A_3321_173#_c_1442_n 0.00965457f $X=16.89
+ $Y=1.665 $X2=0 $Y2=0
cc_864 N_A_2477_543#_c_1309_n N_A_3321_173#_c_1442_n 4.00199e-19 $X=17.16
+ $Y=1.665 $X2=0 $Y2=0
cc_865 N_A_2477_543#_M1020_g N_A_3321_173#_c_1438_n 0.0128134f $X=15.85 $Y=3.275
+ $X2=0 $Y2=0
cc_866 N_A_2477_543#_M1033_g N_A_3321_173#_c_1438_n 0.017148f $X=17.18 $Y=2.75
+ $X2=0 $Y2=0
cc_867 N_A_2477_543#_c_1307_n N_A_3321_173#_c_1439_n 0.0196679f $X=16.89
+ $Y=1.665 $X2=0 $Y2=0
cc_868 N_A_2477_543#_M1033_g N_A_3321_173#_c_1439_n 0.0220724f $X=17.18 $Y=2.75
+ $X2=0 $Y2=0
cc_869 N_A_2477_543#_c_1309_n N_A_3321_173#_c_1439_n 0.0113186f $X=17.16
+ $Y=1.665 $X2=0 $Y2=0
cc_870 N_A_2477_543#_c_1311_n N_A_3321_173#_c_1439_n 0.0125779f $X=16.1 $Y=1.805
+ $X2=0 $Y2=0
cc_871 N_A_2477_543#_c_1309_n N_A_3321_173#_c_1459_n 0.00344989f $X=17.16
+ $Y=1.665 $X2=0 $Y2=0
cc_872 N_A_2477_543#_c_1309_n N_A_3321_173#_c_1434_n 0.0420295f $X=17.16
+ $Y=1.665 $X2=0 $Y2=0
cc_873 N_A_2477_543#_c_1318_n N_VPWR_c_1491_n 0.00940837f $X=12.525 $Y=3.215
+ $X2=0 $Y2=0
cc_874 N_A_2477_543#_c_1318_n N_VPWR_c_1494_n 0.0251241f $X=12.525 $Y=3.215
+ $X2=0 $Y2=0
cc_875 N_A_2477_543#_c_1325_n N_VPWR_c_1494_n 0.00788907f $X=12.835 $Y=2.76
+ $X2=0 $Y2=0
cc_876 N_A_2477_543#_c_1326_n N_VPWR_c_1494_n 0.0143007f $X=14.745 $Y=2.057
+ $X2=0 $Y2=0
cc_877 N_A_2477_543#_M1020_g N_VPWR_c_1497_n 0.0394461f $X=15.85 $Y=3.275 $X2=0
+ $Y2=0
cc_878 N_A_2477_543#_M1033_g N_VPWR_c_1497_n 0.0036421f $X=17.18 $Y=2.75 $X2=0
+ $Y2=0
cc_879 N_A_2477_543#_M1033_g N_VPWR_c_1500_n 0.0769634f $X=17.18 $Y=2.75 $X2=0
+ $Y2=0
cc_880 N_A_2477_543#_M1020_g N_VPWR_c_1503_n 0.00733694f $X=15.85 $Y=3.275 $X2=0
+ $Y2=0
cc_881 N_A_2477_543#_M1033_g N_VPWR_c_1503_n 0.00641794f $X=17.18 $Y=2.75 $X2=0
+ $Y2=0
cc_882 N_A_2477_543#_c_1318_n N_VPWR_c_1503_n 0.0355816f $X=12.525 $Y=3.215
+ $X2=0 $Y2=0
cc_883 N_A_2477_543#_c_1323_n N_VPWR_c_1503_n 0.00209793f $X=14.91 $Y=2.925
+ $X2=0 $Y2=0
cc_884 N_A_2477_543#_c_1325_n N_VPWR_c_1503_n 0.00783169f $X=12.835 $Y=2.76
+ $X2=0 $Y2=0
cc_885 N_A_2477_543#_M1023_g N_VGND_c_1770_n 0.0530386f $X=15.465 $Y=1.075 $X2=0
+ $Y2=0
cc_886 N_A_2477_543#_c_1370_n N_VGND_c_1770_n 0.0256358f $X=15.42 $Y=1.67 $X2=0
+ $Y2=0
cc_887 N_A_2477_543#_c_1326_n N_VGND_c_1770_n 0.0185921f $X=14.745 $Y=2.057
+ $X2=0 $Y2=0
cc_888 N_A_2477_543#_M1032_g N_VGND_c_1772_n 0.0476742f $X=17.14 $Y=1.075 $X2=0
+ $Y2=0
cc_889 N_A_2477_543#_c_1309_n N_VGND_c_1772_n 0.00120691f $X=17.16 $Y=1.665
+ $X2=0 $Y2=0
cc_890 N_A_2477_543#_M1023_g N_VGND_c_1774_n 0.00411567f $X=15.465 $Y=1.075
+ $X2=0 $Y2=0
cc_891 N_A_2477_543#_M1032_g N_VGND_c_1774_n 0.00672879f $X=17.14 $Y=1.075 $X2=0
+ $Y2=0
cc_892 N_A_2477_543#_c_1332_n N_VGND_c_1774_n 0.00250938f $X=12.75 $Y=1.06 $X2=0
+ $Y2=0
cc_893 N_A_3321_173#_c_1438_n N_VPWR_c_1497_n 0.00843468f $X=16.79 $Y=2.52 $X2=0
+ $Y2=0
cc_894 N_A_3321_173#_M1035_g N_VPWR_c_1500_n 0.061155f $X=18.055 $Y=2.875 $X2=0
+ $Y2=0
cc_895 N_A_3321_173#_c_1438_n N_VPWR_c_1500_n 0.0604153f $X=16.79 $Y=2.52 $X2=0
+ $Y2=0
cc_896 N_A_3321_173#_c_1459_n N_VPWR_c_1500_n 0.0267222f $X=17.915 $Y=1.67 $X2=0
+ $Y2=0
cc_897 N_A_3321_173#_c_1434_n N_VPWR_c_1500_n 0.00267375f $X=17.915 $Y=1.67
+ $X2=0 $Y2=0
cc_898 N_A_3321_173#_M1035_g N_VPWR_c_1503_n 0.0125532f $X=18.055 $Y=2.875 $X2=0
+ $Y2=0
cc_899 N_A_3321_173#_c_1438_n N_VPWR_c_1503_n 0.0184574f $X=16.79 $Y=2.52 $X2=0
+ $Y2=0
cc_900 N_A_3321_173#_M1003_g N_Q_c_1748_n 0.0243202f $X=18.035 $Y=0.91 $X2=0
+ $Y2=0
cc_901 N_A_3321_173#_M1035_g N_Q_c_1748_n 0.0283531f $X=18.055 $Y=2.875 $X2=0
+ $Y2=0
cc_902 N_A_3321_173#_c_1459_n N_Q_c_1748_n 0.0489817f $X=17.915 $Y=1.67 $X2=0
+ $Y2=0
cc_903 N_A_3321_173#_c_1434_n N_Q_c_1748_n 0.03769f $X=17.915 $Y=1.67 $X2=0
+ $Y2=0
cc_904 N_A_3321_173#_M1003_g N_VGND_c_1772_n 0.0500684f $X=18.035 $Y=0.91 $X2=0
+ $Y2=0
cc_905 N_A_3321_173#_c_1432_n N_VGND_c_1772_n 0.0379441f $X=16.75 $Y=1.075 $X2=0
+ $Y2=0
cc_906 N_A_3321_173#_c_1433_n N_VGND_c_1772_n 0.0503224f $X=17.75 $Y=1.59 $X2=0
+ $Y2=0
cc_907 N_A_3321_173#_c_1459_n N_VGND_c_1772_n 0.0238914f $X=17.915 $Y=1.67 $X2=0
+ $Y2=0
cc_908 N_A_3321_173#_c_1434_n N_VGND_c_1772_n 0.00165882f $X=17.915 $Y=1.67
+ $X2=0 $Y2=0
cc_909 N_A_3321_173#_M1003_g N_VGND_c_1774_n 0.0136923f $X=18.035 $Y=0.91 $X2=0
+ $Y2=0
cc_910 N_A_3321_173#_c_1432_n N_VGND_c_1774_n 0.0181496f $X=16.75 $Y=1.075 $X2=0
+ $Y2=0
cc_911 N_VPWR_c_1503_n N_A_481_107#_c_1649_n 0.0206009f $X=17.965 $Y=3.59
+ $X2=18.48 $Y2=4.07
cc_912 N_VPWR_c_1482_n N_A_481_107#_c_1617_n 0.00461337f $X=4.15 $Y=2.97
+ $X2=9.36 $Y2=4.013
cc_913 N_VPWR_c_1482_n N_A_481_107#_c_1618_n 0.0678227f $X=4.15 $Y=2.97 $X2=0
+ $Y2=0
cc_914 N_VPWR_c_1482_n N_A_481_107#_c_1673_n 0.0579547f $X=4.15 $Y=2.97 $X2=0
+ $Y2=0
cc_915 N_VPWR_c_1503_n N_A_481_107#_c_1673_n 0.0190146f $X=17.965 $Y=3.59 $X2=0
+ $Y2=0
cc_916 N_VPWR_c_1485_n N_A_481_107#_c_1619_n 0.0047991f $X=5.64 $Y=2.79 $X2=0
+ $Y2=0
cc_917 N_VPWR_c_1503_n N_A_481_107#_c_1619_n 0.0279566f $X=17.965 $Y=3.59 $X2=0
+ $Y2=0
cc_918 N_VPWR_c_1482_n N_A_481_107#_c_1622_n 0.00433879f $X=4.15 $Y=2.97 $X2=0
+ $Y2=0
cc_919 N_VPWR_c_1503_n N_A_481_107#_c_1622_n 0.00754921f $X=17.965 $Y=3.59 $X2=0
+ $Y2=0
cc_920 N_VPWR_c_1485_n N_A_481_107#_c_1625_n 0.0711742f $X=5.64 $Y=2.79 $X2=0
+ $Y2=0
cc_921 N_VPWR_c_1503_n N_A_481_107#_c_1625_n 0.0194693f $X=17.965 $Y=3.59 $X2=0
+ $Y2=0
cc_922 N_VPWR_c_1485_n N_A_481_107#_c_1626_n 0.0137562f $X=5.64 $Y=2.79 $X2=0
+ $Y2=0
cc_923 N_VPWR_c_1485_n N_A_481_107#_c_1628_n 0.0413753f $X=5.64 $Y=2.79 $X2=0
+ $Y2=0
cc_924 N_VPWR_c_1503_n N_A_481_107#_c_1628_n 0.0195984f $X=17.965 $Y=3.59 $X2=0
+ $Y2=0
cc_925 N_VPWR_c_1503_n N_A_481_107#_c_1629_n 0.0399246f $X=17.965 $Y=3.59 $X2=0
+ $Y2=0
cc_926 N_VPWR_c_1485_n N_A_481_107#_c_1632_n 0.0047991f $X=5.64 $Y=2.79 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1503_n N_A_481_107#_c_1632_n 0.00659047f $X=17.965 $Y=3.59 $X2=0
+ $Y2=0
cc_928 N_VPWR_c_1503_n N_A_481_107#_c_1636_n 0.0395567f $X=17.965 $Y=3.59 $X2=0
+ $Y2=0
cc_929 N_VPWR_c_1503_n N_A_481_107#_c_1637_n 0.0182755f $X=17.965 $Y=3.59 $X2=0
+ $Y2=0
cc_930 N_VPWR_c_1488_n A_1686_543# 0.00285177f $X=9.28 $Y=3.01 $X2=0 $Y2=3.985
cc_931 N_VPWR_c_1491_n A_2335_543# 0.00617484f $X=11.67 $Y=3.59 $X2=0 $Y2=3.985
cc_932 N_VPWR_c_1503_n A_2335_543# 0.00106357f $X=17.965 $Y=3.59 $X2=0 $Y2=3.985
cc_933 N_VPWR_c_1500_n N_Q_c_1748_n 0.0792609f $X=17.665 $Y=2.52 $X2=9.36
+ $Y2=4.07
cc_934 N_VPWR_c_1503_n N_Q_c_1748_n 0.0152638f $X=17.965 $Y=3.59 $X2=9.36
+ $Y2=4.07
cc_935 N_A_481_107#_c_1611_n N_VGND_c_1762_n 0.00461337f $X=3.155 $Y=2.455 $X2=0
+ $Y2=0
cc_936 N_A_481_107#_c_1610_n N_VGND_c_1774_n 0.01835f $X=3.07 $Y=0.83 $X2=0
+ $Y2=0
cc_937 N_A_481_107#_c_1612_n N_VGND_c_1774_n 0.0273048f $X=2.545 $Y=0.745 $X2=0
+ $Y2=0
cc_938 N_A_481_107#_c_1614_n N_VGND_c_1774_n 0.0220791f $X=6.715 $Y=0.78 $X2=0
+ $Y2=0
cc_939 N_Q_c_1748_n N_VGND_c_1772_n 0.0528446f $X=18.425 $Y=0.66 $X2=0 $Y2=0
cc_940 N_Q_c_1748_n N_VGND_c_1774_n 0.0351041f $X=18.425 $Y=0.66 $X2=0 $Y2=0
cc_941 N_VGND_c_1774_n A_339_107# 0.00261802f $X=17.93 $Y=0.48 $X2=0 $Y2=0
cc_942 N_VGND_c_1774_n A_637_107# 0.00691792f $X=17.93 $Y=0.48 $X2=0 $Y2=0
cc_943 N_VGND_c_1766_n A_1627_113# 0.00576077f $X=9.035 $Y=0.48 $X2=0 $Y2=0
cc_944 N_VGND_c_1774_n A_1627_113# 0.00271077f $X=17.93 $Y=0.48 $X2=0 $Y2=0
cc_945 N_VGND_c_1774_n A_2035_107# 0.00663096f $X=17.93 $Y=0.48 $X2=0 $Y2=0
cc_946 N_VGND_c_1774_n A_2352_107# 0.00875788f $X=17.93 $Y=0.48 $X2=0 $Y2=0
