* File: sky130_fd_sc_hvl__a21oi_1.pex.spice
* Created: Fri Aug 28 09:32:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__A21OI_1%VNB 5 7 11 25
c20 11 0 1.16365e-19 $X=0.24 $Y=0
r21 7 25 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0.058
r22 7 11 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0
r23 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r24 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__A21OI_1%VPB 4 6 14 21
r28 10 21 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=4.07
+ $X2=1.68 $Y2=4.013
r29 10 14 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=4.07
+ $X2=3.12 $Y2=4.07
r30 9 14 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=3.12 $Y2=4.07
r31 9 10 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r32 6 21 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=4.012
+ $X2=1.68 $Y2=4.013
r33 4 14 52 $w=1.7e-07 $l=3.16221e-06 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=3.12 $Y2=4.07
r34 4 9 52 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__A21OI_1%A2 3 7 9 10 11 20
r23 19 20 23.158 $w=6.7e-07 $l=2.9e-07 $layer=POLY_cond $X=0.815 $Y=1.75
+ $X2=1.105 $Y2=1.75
r24 16 19 5.19058 $w=6.7e-07 $l=6.5e-08 $layer=POLY_cond $X=0.75 $Y=1.75
+ $X2=0.815 $Y2=1.75
r25 10 11 22.5785 $w=2.43e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.627
+ $X2=1.2 $Y2=1.627
r26 10 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.625 $X2=0.75 $Y2=1.625
r27 9 10 22.5785 $w=2.43e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.627
+ $X2=0.72 $Y2=1.627
r28 5 20 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.105 $Y=1.415
+ $X2=1.105 $Y2=1.75
r29 5 7 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.105 $Y=1.415 $X2=1.105
+ $Y2=0.91
r30 1 19 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.815 $Y=2.085
+ $X2=0.815 $Y2=1.75
r31 1 3 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.815 $Y=2.085 $X2=0.815
+ $Y2=2.965
.ends

.subckt PM_SKY130_FD_SC_HVL__A21OI_1%A1 1 4 10
c26 4 0 1.16365e-19 $X=1.815 $Y=0.91
r27 7 10 142.853 $w=5e-07 $l=1.335e-06 $layer=POLY_cond $X=1.815 $Y=1.63
+ $X2=1.815 $Y2=2.965
r28 4 7 77.0442 $w=5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.815 $Y=0.91 $X2=1.815
+ $Y2=1.63
r29 1 7 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75 $Y=1.63
+ $X2=1.75 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HVL__A21OI_1%B1 3 6 7 8 9 10 16 17 18 19
r28 16 19 20.8158 $w=6e-07 $l=2.15e-07 $layer=POLY_cond $X=2.645 $Y=1.89
+ $X2=2.645 $Y2=2.105
r29 16 18 45.7838 $w=6e-07 $l=4.95e-07 $layer=POLY_cond $X=2.645 $Y=1.89
+ $X2=2.645 $Y2=1.395
r30 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.635
+ $Y=1.89 $X2=2.635 $Y2=1.89
r31 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.635 $Y=2.775
+ $X2=2.635 $Y2=3.145
r32 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.635 $Y=2.405
+ $X2=2.635 $Y2=2.775
r33 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.635 $Y=2.035
+ $X2=2.635 $Y2=2.405
r34 7 17 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.635 $Y=2.035
+ $X2=2.635 $Y2=1.89
r35 6 18 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.695 $Y=0.91 $X2=2.695
+ $Y2=1.395
r36 3 19 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.595 $Y=2.965 $X2=2.595
+ $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_HVL__A21OI_1%A_56_443# 1 2 9 13 14 17
r29 17 19 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.205 $Y=2.34
+ $X2=2.205 $Y2=3.59
r30 15 17 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.205 $Y=2.1
+ $X2=2.205 $Y2=2.34
r31 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.12 $Y=2.015
+ $X2=2.205 $Y2=2.1
r32 13 14 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=2.12 $Y=2.015
+ $X2=0.51 $Y2=2.015
r33 9 11 57.6222 $w=2.48e-07 $l=1.25e-06 $layer=LI1_cond $X=0.385 $Y=2.34
+ $X2=0.385 $Y2=3.59
r34 7 14 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.385 $Y=2.1
+ $X2=0.51 $Y2=2.015
r35 7 9 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=0.385 $Y=2.1 $X2=0.385
+ $Y2=2.34
r36 2 19 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.065
+ $Y=2.215 $X2=2.205 $Y2=3.59
r37 2 17 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.065
+ $Y=2.215 $X2=2.205 $Y2=2.34
r38 1 11 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.28
+ $Y=2.215 $X2=0.425 $Y2=3.59
r39 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.28
+ $Y=2.215 $X2=0.425 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__A21OI_1%VPWR 1 4 7 14
r22 10 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.855 $Y=3.59
+ $X2=1.855 $Y2=3.59
r23 10 11 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.775 $Y=3.59
+ $X2=0.775 $Y2=3.59
r24 7 10 11.956 $w=1.248e-06 $l=1.225e-06 $layer=LI1_cond $X=1.315 $Y=2.365
+ $X2=1.315 $Y2=3.59
r25 4 14 0.0671834 $w=3.7e-07 $l=1.75e-07 $layer=MET1_cond $X=1.68 $Y=3.63
+ $X2=1.855 $Y2=3.63
r26 4 11 0.347434 $w=3.7e-07 $l=9.05e-07 $layer=MET1_cond $X=1.68 $Y=3.63
+ $X2=0.775 $Y2=3.63
r27 1 10 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.065
+ $Y=2.215 $X2=1.205 $Y2=3.59
r28 1 7 300 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=2 $X=1.065
+ $Y=2.215 $X2=1.205 $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_HVL__A21OI_1%Y 1 2 9 11 12 13 14 15 16 17 24 26
r29 24 26 1.80775 $w=2.53e-07 $l=4e-08 $layer=LI1_cond $X=3.107 $Y=1.625
+ $X2=3.107 $Y2=1.665
r30 17 38 20.1113 $w=2.53e-07 $l=4.45e-07 $layer=LI1_cond $X=3.107 $Y=3.145
+ $X2=3.107 $Y2=3.59
r31 16 17 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.107 $Y=2.775
+ $X2=3.107 $Y2=3.145
r32 15 16 19.6593 $w=2.53e-07 $l=4.35e-07 $layer=LI1_cond $X=3.107 $Y=2.34
+ $X2=3.107 $Y2=2.775
r33 14 15 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=3.107 $Y=2.035
+ $X2=3.107 $Y2=2.34
r34 13 24 2.87766 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.107 $Y=1.54
+ $X2=3.107 $Y2=1.625
r35 13 14 15.7275 $w=2.53e-07 $l=3.48e-07 $layer=LI1_cond $X=3.107 $Y=1.687
+ $X2=3.107 $Y2=2.035
r36 13 26 0.994265 $w=2.53e-07 $l=2.2e-08 $layer=LI1_cond $X=3.107 $Y=1.687
+ $X2=3.107 $Y2=1.665
r37 11 13 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.98 $Y=1.54
+ $X2=3.107 $Y2=1.54
r38 11 12 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.98 $Y=1.54
+ $X2=2.47 $Y2=1.54
r39 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.345 $Y=1.455
+ $X2=2.47 $Y2=1.54
r40 7 9 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=2.345 $Y=1.455
+ $X2=2.345 $Y2=0.66
r41 2 38 300 $w=1.7e-07 $l=1.48092e-06 $layer=licon1_PDIFF $count=2 $X=2.845
+ $Y=2.215 $X2=3.065 $Y2=3.59
r42 2 15 300 $w=1.7e-07 $l=2.755e-07 $layer=licon1_PDIFF $count=2 $X=2.845
+ $Y=2.215 $X2=3.065 $Y2=2.34
r43 1 9 91 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=2 $X=2.065
+ $Y=0.535 $X2=2.305 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__A21OI_1%VGND 1 2 7 16 20 21
r23 20 24 4.0545 $w=5.88e-07 $l=2e-07 $layer=LI1_cond $X=2.97 $Y=0.48 $X2=2.97
+ $Y2=0.68
r24 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.15 $Y=0.48
+ $X2=3.15 $Y2=0.48
r25 17 21 0.477962 $w=3.7e-07 $l=1.245e-06 $layer=MET1_cond $X=1.905 $Y=0.44
+ $X2=3.15 $Y2=0.44
r26 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.905 $Y=0.48
+ $X2=1.905 $Y2=0.48
r27 14 16 15.1229 $w=9.58e-07 $l=1.19e-06 $layer=LI1_cond $X=0.715 $Y=0.845
+ $X2=1.905 $Y2=0.845
r28 10 14 3.17708 $w=9.58e-07 $l=2.5e-07 $layer=LI1_cond $X=0.465 $Y=0.845
+ $X2=0.715 $Y2=0.845
r29 10 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.465 $Y=0.48
+ $X2=0.465 $Y2=0.48
r30 7 17 0.0863787 $w=3.7e-07 $l=2.25e-07 $layer=MET1_cond $X=1.68 $Y=0.44
+ $X2=1.905 $Y2=0.44
r31 7 11 0.466445 $w=3.7e-07 $l=1.215e-06 $layer=MET1_cond $X=1.68 $Y=0.44
+ $X2=0.465 $Y2=0.44
r32 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.535 $X2=3.085 $Y2=0.68
r33 1 14 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.535 $X2=0.715 $Y2=0.66
.ends

