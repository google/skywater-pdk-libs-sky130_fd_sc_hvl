* File: sky130_fd_sc_hvl__probec_p_8.pex.spice
* Created: Fri Aug 28 09:39:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__PROBEC_P_8%VNB 5 7 11 25
r49 7 25 1.30208e-05 $w=9.6e-06 $l=1e-09 $layer=MET1_cond $X=4.8 $Y=0.057
+ $X2=4.8 $Y2=0.058
r50 7 11 0.000742187 $w=9.6e-06 $l=5.7e-08 $layer=MET1_cond $X=4.8 $Y=0.057
+ $X2=4.8 $Y2=0
r51 5 11 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r52 5 11 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBEC_P_8%VPB 4 6 14 21
c91 4 0 1.06581e-19 $X=-0.33 $Y=1.885
r92 10 21 0.000742187 $w=9.6e-06 $l=5.7e-08 $layer=MET1_cond $X=4.8 $Y=4.07
+ $X2=4.8 $Y2=4.013
r93 10 14 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=9.36 $Y=4.07
+ $X2=9.36 $Y2=4.07
r94 9 14 594.995 $w=1.68e-07 $l=9.12e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=9.36 $Y2=4.07
r95 9 10 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r96 6 21 1.30208e-05 $w=9.6e-06 $l=1e-09 $layer=MET1_cond $X=4.8 $Y=4.012
+ $X2=4.8 $Y2=4.013
r97 4 14 18.2 $w=1.7e-07 $l=9.4024e-06 $layer=licon1_NTAP_notbjt $count=10 $X=0
+ $Y=3.985 $X2=9.36 $Y2=4.07
r98 4 9 18.2 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=10 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBEC_P_8%A 3 5 7 8 10 12 15 17 19 22 24 25 26 27
+ 28 37
c85 15 0 1.43567e-19 $X=1.82 $Y=2.965
r86 36 37 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.82 $Y=1.815 $X2=2.6
+ $Y2=1.815
r87 34 36 9.0955 $w=5e-07 $l=8.5e-08 $layer=POLY_cond $X=1.735 $Y=1.815 $X2=1.82
+ $Y2=1.815
r88 27 28 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.697
+ $X2=2.16 $Y2=1.697
r89 27 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.735
+ $Y=1.73 $X2=1.735 $Y2=1.73
r90 26 27 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.697
+ $X2=1.68 $Y2=1.697
r91 25 26 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.697
+ $X2=1.2 $Y2=1.697
r92 20 37 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.6 $Y=2.065 $X2=2.6
+ $Y2=1.815
r93 20 22 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=2.6 $Y=2.065 $X2=2.6
+ $Y2=2.965
r94 17 37 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.6 $Y=1.565 $X2=2.6
+ $Y2=1.815
r95 17 19 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.6 $Y=1.565 $X2=2.6
+ $Y2=1.08
r96 13 36 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.82 $Y=2.065 $X2=1.82
+ $Y2=1.815
r97 13 15 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=1.82 $Y=2.065 $X2=1.82
+ $Y2=2.965
r98 10 36 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.82 $Y=1.565 $X2=1.82
+ $Y2=1.815
r99 10 12 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.82 $Y=1.565 $X2=1.82
+ $Y2=1.08
r100 9 24 5.30422 $w=5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.03 $Y=1.815 $X2=0.77
+ $Y2=1.815
r101 8 34 17.656 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.815
+ $X2=1.735 $Y2=1.815
r102 8 9 57.7832 $w=5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.57 $Y=1.815 $X2=1.03
+ $Y2=1.815
r103 5 24 20.4101 $w=5e-07 $l=2.54951e-07 $layer=POLY_cond $X=0.78 $Y=1.565
+ $X2=0.77 $Y2=1.815
r104 5 7 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.78 $Y=1.565 $X2=0.78
+ $Y2=1.08
r105 1 24 20.4101 $w=5e-07 $l=2.54951e-07 $layer=POLY_cond $X=0.76 $Y=2.065
+ $X2=0.77 $Y2=1.815
r106 1 3 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=0.76 $Y=2.065 $X2=0.76
+ $Y2=2.965
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBEC_P_8%A_45_443# 1 2 3 4 15 17 19 22 24 26 29
+ 31 33 36 38 40 43 45 47 50 52 54 57 59 61 64 66 68 71 74 77 81 85 91 94 96 99
+ 102 103 104 107 109 119
c260 94 0 1.82353e-19 $X=2.51 $Y=1.625
c261 91 0 6.98013e-20 $X=2.21 $Y=0.895
c262 71 0 1.17159e-19 $X=0.37 $Y=0.97
c263 59 0 1.125e-19 $X=8.06 $Y=2.105
c264 57 0 1.2129e-19 $X=8.06 $Y=1.08
c265 52 0 1.29061e-19 $X=7.28 $Y=2.105
r266 118 119 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=8.06 $Y=1.855
+ $X2=8.84 $Y2=1.855
r267 117 118 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.28 $Y=1.855
+ $X2=8.06 $Y2=1.855
r268 116 117 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=6.5 $Y=1.855
+ $X2=7.28 $Y2=1.855
r269 115 116 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=5.72 $Y=1.855
+ $X2=6.5 $Y2=1.855
r270 114 115 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=4.94 $Y=1.855
+ $X2=5.72 $Y2=1.855
r271 113 114 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=4.16 $Y=1.855
+ $X2=4.94 $Y2=1.855
r272 112 113 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.38 $Y=1.855
+ $X2=4.16 $Y2=1.855
r273 100 112 9.0955 $w=5e-07 $l=8.5e-08 $layer=POLY_cond $X=3.295 $Y=1.855
+ $X2=3.38 $Y2=1.855
r274 99 100 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.295
+ $Y=1.79 $X2=3.295 $Y2=1.79
r275 97 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.79
+ $X2=2.51 $Y2=1.79
r276 97 99 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.595 $Y=1.79
+ $X2=3.295 $Y2=1.79
r277 96 104 2.66603 $w=3.6e-07 $l=2.28583e-07 $layer=LI1_cond $X=2.51 $Y=2.095
+ $X2=2.32 $Y2=2.18
r278 95 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=1.955
+ $X2=2.51 $Y2=1.79
r279 95 96 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.51 $Y=1.955
+ $X2=2.51 $Y2=2.095
r280 94 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=1.625
+ $X2=2.51 $Y2=1.79
r281 93 107 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=1.4
+ $X2=2.51 $Y2=1.315
r282 93 94 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.51 $Y=1.4
+ $X2=2.51 $Y2=1.625
r283 89 107 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.21 $Y=1.315
+ $X2=2.51 $Y2=1.315
r284 89 91 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=2.21 $Y=1.23
+ $X2=2.21 $Y2=0.895
r285 85 87 22.1818 $w=5.48e-07 $l=1.02e-06 $layer=LI1_cond $X=2.32 $Y=2.34
+ $X2=2.32 $Y2=3.36
r286 83 104 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.32 $Y=2.265
+ $X2=2.32 $Y2=2.18
r287 83 85 1.63102 $w=5.48e-07 $l=7.5e-08 $layer=LI1_cond $X=2.32 $Y=2.265
+ $X2=2.32 $Y2=2.34
r288 82 103 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.435 $Y=2.18
+ $X2=0.34 $Y2=2.18
r289 81 104 4.14084 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.045 $Y=2.18
+ $X2=2.32 $Y2=2.18
r290 81 82 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=2.045 $Y=2.18
+ $X2=0.435 $Y2=2.18
r291 77 79 59.5407 $w=1.88e-07 $l=1.02e-06 $layer=LI1_cond $X=0.34 $Y=2.36
+ $X2=0.34 $Y2=3.38
r292 75 103 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.34 $Y=2.265
+ $X2=0.34 $Y2=2.18
r293 75 77 5.54545 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=0.34 $Y=2.265
+ $X2=0.34 $Y2=2.36
r294 74 103 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.34 $Y=2.095
+ $X2=0.34 $Y2=2.18
r295 74 102 36.1914 $w=1.88e-07 $l=6.2e-07 $layer=LI1_cond $X=0.34 $Y=2.095
+ $X2=0.34 $Y2=1.475
r296 69 102 5.66915 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=0.35 $Y=1.37
+ $X2=0.35 $Y2=1.475
r297 69 71 21.1255 $w=2.08e-07 $l=4e-07 $layer=LI1_cond $X=0.35 $Y=1.37 $X2=0.35
+ $Y2=0.97
r298 66 119 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.84 $Y=2.105
+ $X2=8.84 $Y2=1.855
r299 66 68 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.84 $Y=2.105 $X2=8.84
+ $Y2=2.965
r300 62 119 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.84 $Y=1.605
+ $X2=8.84 $Y2=1.855
r301 62 64 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=8.84 $Y=1.605
+ $X2=8.84 $Y2=1.08
r302 59 118 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.06 $Y=2.105
+ $X2=8.06 $Y2=1.855
r303 59 61 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.06 $Y=2.105 $X2=8.06
+ $Y2=2.965
r304 55 118 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.06 $Y=1.605
+ $X2=8.06 $Y2=1.855
r305 55 57 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=8.06 $Y=1.605
+ $X2=8.06 $Y2=1.08
r306 52 117 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.28 $Y=2.105
+ $X2=7.28 $Y2=1.855
r307 52 54 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.28 $Y=2.105 $X2=7.28
+ $Y2=2.965
r308 48 117 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.28 $Y=1.605
+ $X2=7.28 $Y2=1.855
r309 48 50 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=7.28 $Y=1.605
+ $X2=7.28 $Y2=1.08
r310 45 116 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.5 $Y=2.105 $X2=6.5
+ $Y2=1.855
r311 45 47 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.5 $Y=2.105 $X2=6.5
+ $Y2=2.965
r312 41 116 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.5 $Y=1.605 $X2=6.5
+ $Y2=1.855
r313 41 43 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=6.5 $Y=1.605 $X2=6.5
+ $Y2=1.08
r314 38 115 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.72 $Y=2.105
+ $X2=5.72 $Y2=1.855
r315 38 40 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.72 $Y=2.105 $X2=5.72
+ $Y2=2.965
r316 34 115 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.72 $Y=1.605
+ $X2=5.72 $Y2=1.855
r317 34 36 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=5.72 $Y=1.605
+ $X2=5.72 $Y2=1.08
r318 31 114 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.94 $Y=2.105
+ $X2=4.94 $Y2=1.855
r319 31 33 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.94 $Y=2.105 $X2=4.94
+ $Y2=2.965
r320 27 114 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.94 $Y=1.605
+ $X2=4.94 $Y2=1.855
r321 27 29 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.94 $Y=1.605
+ $X2=4.94 $Y2=1.08
r322 24 113 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.16 $Y=2.105
+ $X2=4.16 $Y2=1.855
r323 24 26 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.16 $Y=2.105 $X2=4.16
+ $Y2=2.965
r324 20 113 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.16 $Y=1.605
+ $X2=4.16 $Y2=1.855
r325 20 22 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.16 $Y=1.605
+ $X2=4.16 $Y2=1.08
r326 17 112 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.38 $Y=2.105
+ $X2=3.38 $Y2=1.855
r327 17 19 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.38 $Y=2.105 $X2=3.38
+ $Y2=2.965
r328 13 112 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.38 $Y=1.605
+ $X2=3.38 $Y2=1.855
r329 13 15 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.38 $Y=1.605
+ $X2=3.38 $Y2=1.08
r330 4 87 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=2.07
+ $Y=2.215 $X2=2.21 $Y2=3.36
r331 4 85 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.07
+ $Y=2.215 $X2=2.21 $Y2=2.34
r332 3 79 300 $w=1.7e-07 $l=1.22591e-06 $layer=licon1_PDIFF $count=2 $X=0.225
+ $Y=2.215 $X2=0.35 $Y2=3.38
r333 3 77 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.225
+ $Y=2.215 $X2=0.35 $Y2=2.36
r334 2 91 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=2.07
+ $Y=0.705 $X2=2.21 $Y2=0.895
r335 1 71 91 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=2 $X=0.245
+ $Y=0.705 $X2=0.37 $Y2=0.97
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBEC_P_8%VPWR 1 2 3 4 5 6 19 21 23 25 29 31 36 38
+ 40 42 43 58 68 80 92 102 117 124 125 127 142
c159 125 0 1.86017e-19 $X=9.76 $Y=3.635
r160 125 130 0.16865 $w=2.8e-07 $l=3.2e-07 $layer=MET2_cond $X=9.76 $Y=3.645
+ $X2=9.44 $Y2=3.645
r161 124 125 4.5 $w=1.5e-07 $l=1.5e-07 $layer=via $count=1 $X=9.76 $Y=3.635
+ $X2=9.76 $Y2=3.635
r162 120 127 0.0249539 $w=3.7e-07 $l=6.5e-08 $layer=MET1_cond $X=9.35 $Y=3.63
+ $X2=9.415 $Y2=3.63
r163 116 117 14.2225 $w=3.18e-07 $l=3.25e-07 $layer=LI1_cond $X=9.23 $Y=3.635
+ $X2=8.905 $Y2=3.635
r164 112 113 1.3664 $w=1.248e-06 $l=1.4e-07 $layer=LI1_cond $X=1.24 $Y=3.57
+ $X2=1.24 $Y2=3.71
r165 108 110 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=1.42 $Y=3.63
+ $X2=1.78 $Y2=3.63
r166 106 108 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.7 $Y=3.63
+ $X2=1.42 $Y2=3.63
r167 105 112 0.0976 $w=1.248e-06 $l=1e-08 $layer=LI1_cond $X=1.24 $Y=3.56
+ $X2=1.24 $Y2=3.57
r168 105 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.78 $Y=3.56
+ $X2=1.78 $Y2=3.56
r169 105 108 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.42 $Y=3.56
+ $X2=1.42 $Y2=3.56
r170 105 106 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.7 $Y=3.56
+ $X2=0.7 $Y2=3.56
r171 102 105 9.8576 $w=1.248e-06 $l=1.01e-06 $layer=LI1_cond $X=1.24 $Y=2.55
+ $X2=1.24 $Y2=3.56
r172 98 120 0.506755 $w=3.7e-07 $l=1.32e-06 $layer=MET1_cond $X=8.03 $Y=3.63
+ $X2=9.35 $Y2=3.63
r173 96 98 0.274492 $w=3.7e-07 $l=7.15e-07 $layer=MET1_cond $X=7.315 $Y=3.63
+ $X2=8.03 $Y2=3.63
r174 95 100 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=7.67 $Y=3.56
+ $X2=7.67 $Y2=3.57
r175 95 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.03 $Y=3.56
+ $X2=8.03 $Y2=3.56
r176 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.315 $Y=3.56
+ $X2=7.315 $Y2=3.56
r177 92 95 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=7.67 $Y=2.55
+ $X2=7.67 $Y2=3.56
r178 88 96 0.3244 $w=3.7e-07 $l=8.45e-07 $layer=MET1_cond $X=6.47 $Y=3.63
+ $X2=7.315 $Y2=3.63
r179 86 88 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=6.11 $Y=3.63
+ $X2=6.47 $Y2=3.63
r180 84 86 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=5.75 $Y=3.63
+ $X2=6.11 $Y2=3.63
r181 83 90 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=6.11 $Y=3.56
+ $X2=6.11 $Y2=3.57
r182 83 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.47 $Y=3.56
+ $X2=6.47 $Y2=3.56
r183 83 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.11 $Y=3.56
+ $X2=6.11 $Y2=3.56
r184 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=3.56
+ $X2=5.75 $Y2=3.56
r185 80 83 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=6.11 $Y=2.55
+ $X2=6.11 $Y2=3.56
r186 76 84 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=4.91 $Y=3.63
+ $X2=5.75 $Y2=3.63
r187 76 142 0.0422296 $w=3.7e-07 $l=1.1e-07 $layer=MET1_cond $X=4.91 $Y=3.63
+ $X2=4.8 $Y2=3.63
r188 72 74 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=4.19 $Y=3.63
+ $X2=4.55 $Y2=3.63
r189 71 78 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=4.55 $Y=3.56
+ $X2=4.55 $Y2=3.57
r190 71 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.91 $Y=3.56
+ $X2=4.91 $Y2=3.56
r191 71 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.55 $Y=3.56
+ $X2=4.55 $Y2=3.56
r192 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.19 $Y=3.56
+ $X2=4.19 $Y2=3.56
r193 68 71 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=4.55 $Y=2.55
+ $X2=4.55 $Y2=3.56
r194 64 72 0.374308 $w=3.7e-07 $l=9.75e-07 $layer=MET1_cond $X=3.215 $Y=3.63
+ $X2=4.19 $Y2=3.63
r195 62 64 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=2.855 $Y=3.63
+ $X2=3.215 $Y2=3.63
r196 62 110 0.412698 $w=3.7e-07 $l=1.075e-06 $layer=MET1_cond $X=2.855 $Y=3.63
+ $X2=1.78 $Y2=3.63
r197 61 66 0.178519 $w=6.68e-07 $l=1e-08 $layer=LI1_cond $X=3.1 $Y=3.56 $X2=3.1
+ $Y2=3.57
r198 61 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.215 $Y=3.56
+ $X2=3.215 $Y2=3.56
r199 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.855 $Y=3.56
+ $X2=2.855 $Y2=3.56
r200 58 61 18.0304 $w=6.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.1 $Y=2.55
+ $X2=3.1 $Y2=3.56
r201 43 142 0.0357032 $w=3.7e-07 $l=9.3e-08 $layer=MET1_cond $X=4.707 $Y=3.63
+ $X2=4.8 $Y2=3.63
r202 43 74 0.0602731 $w=3.7e-07 $l=1.57e-07 $layer=MET1_cond $X=4.707 $Y=3.63
+ $X2=4.55 $Y2=3.63
r203 43 127 0.00959763 $w=3.7e-07 $l=2.5e-08 $layer=MET1_cond $X=9.44 $Y=3.63
+ $X2=9.415 $Y2=3.63
r204 43 130 4.5 $w=1.5e-07 $l=1.5e-07 $layer=via $count=1 $X=9.44 $Y=3.635
+ $X2=9.44 $Y2=3.635
r205 43 124 0.0761468 $w=5.2e-07 $l=1.6e-07 $layer=MET1_cond $X=9.6 $Y=3.635
+ $X2=9.76 $Y2=3.635
r206 41 100 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=7.67 $Y=3.625
+ $X2=7.67 $Y2=3.57
r207 41 42 3.33002 $w=8.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.67 $Y=3.625
+ $X2=7.67 $Y2=3.71
r208 39 90 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6.11 $Y=3.625
+ $X2=6.11 $Y2=3.57
r209 39 40 3.33002 $w=8.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.11 $Y=3.625
+ $X2=6.11 $Y2=3.71
r210 37 78 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=4.55 $Y=3.625
+ $X2=4.55 $Y2=3.57
r211 37 38 3.33002 $w=8.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=3.625
+ $X2=4.55 $Y2=3.71
r212 35 66 0.981855 $w=6.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.1 $Y=3.625
+ $X2=3.1 $Y2=3.57
r213 35 36 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=3.625 $X2=3.1
+ $Y2=3.71
r214 31 34 21.18 $w=3.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.32 $Y=2.55 $X2=9.32
+ $Y2=3.23
r215 29 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.35 $Y=3.56
+ $X2=9.35 $Y2=3.56
r216 29 116 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=9.32 $Y=3.635
+ $X2=9.23 $Y2=3.635
r217 29 34 7.63104 $w=3.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.32 $Y=3.475
+ $X2=9.32 $Y2=3.23
r218 28 42 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=8.115 $Y=3.71
+ $X2=7.67 $Y2=3.71
r219 28 117 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.115 $Y=3.71
+ $X2=8.905 $Y2=3.71
r220 26 40 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=6.555 $Y=3.71
+ $X2=6.11 $Y2=3.71
r221 25 42 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=7.225 $Y=3.71
+ $X2=7.67 $Y2=3.71
r222 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.225 $Y=3.71
+ $X2=6.555 $Y2=3.71
r223 24 38 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=4.995 $Y=3.71
+ $X2=4.55 $Y2=3.71
r224 23 40 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=5.665 $Y=3.71
+ $X2=6.11 $Y2=3.71
r225 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.665 $Y=3.71
+ $X2=4.995 $Y2=3.71
r226 22 36 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.435 $Y=3.71
+ $X2=3.1 $Y2=3.71
r227 21 38 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=4.105 $Y=3.71
+ $X2=4.55 $Y2=3.71
r228 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.105 $Y=3.71
+ $X2=3.435 $Y2=3.71
r229 20 113 13.277 $w=1.7e-07 $l=6.25e-07 $layer=LI1_cond $X=1.865 $Y=3.71
+ $X2=1.24 $Y2=3.71
r230 19 36 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.765 $Y=3.71
+ $X2=3.1 $Y2=3.71
r231 19 20 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.765 $Y=3.71
+ $X2=1.865 $Y2=3.71
r232 6 116 600 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=1 $X=9.09
+ $Y=2.215 $X2=9.23 $Y2=3.57
r233 6 34 400 $w=1.7e-07 $l=1.08274e-06 $layer=licon1_PDIFF $count=1 $X=9.09
+ $Y=2.215 $X2=9.23 $Y2=3.23
r234 6 31 400 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=9.09
+ $Y=2.215 $X2=9.23 $Y2=2.55
r235 5 100 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=7.53
+ $Y=2.215 $X2=7.67 $Y2=3.57
r236 5 92 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=7.53
+ $Y=2.215 $X2=7.67 $Y2=2.55
r237 4 90 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=5.97
+ $Y=2.215 $X2=6.11 $Y2=3.57
r238 4 80 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=5.97
+ $Y=2.215 $X2=6.11 $Y2=2.55
r239 3 78 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=4.41
+ $Y=2.215 $X2=4.55 $Y2=3.57
r240 3 68 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=4.41
+ $Y=2.215 $X2=4.55 $Y2=2.55
r241 2 66 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=2.85
+ $Y=2.215 $X2=2.99 $Y2=3.57
r242 2 58 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=2.85
+ $Y=2.215 $X2=2.99 $Y2=2.55
r243 1 112 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=2.215 $X2=1.15 $Y2=3.57
r244 1 102 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=2.215 $X2=1.15 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBEC_P_8%noxref_6 1 2 3 4 5 6 7 8 27 33 35 39 45
+ 49 55 57 60 62 65 67 69 70 71 72 76 80 82 88 93
c159 82 0 5.55441e-20 $X=4.26 $Y=2.035
c160 76 0 1.06581e-19 $X=5.6 $Y=2.035
r161 88 93 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=6.05 $Y=2.035
+ $X2=6.05 $Y2=2.035
r162 85 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.065 $Y=2.035
+ $X2=6.065 $Y2=2.035
r163 80 93 1.705 $w=2e-07 $l=4e-07 $layer=via2 $count=2 $X=6.025 $Y=2.035
+ $X2=6.025 $Y2=2.035
r164 77 82 0.0203094 $w=4.097e-06 $l=1.34e-06 $layer=MET5_cond $X=5.6 $Y=2.035
+ $X2=4.26 $Y2=2.035
r165 76 80 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=6.025
+ $Y=2.035 $X2=6.025 $Y2=2.035
r166 76 77 0.38 $w=8e-07 $l=8e-07 $layer=via4_notcap2m $count=1 $X=5.6 $Y=2.035
+ $X2=5.6 $Y2=2.035
r167 70 85 13.6105 $w=5.78e-07 $l=6.6e-07 $layer=LI1_cond $X=6.725 $Y=1.915
+ $X2=6.065 $Y2=1.915
r168 70 71 1.08702 $w=5.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=1.915
+ $X2=6.89 $Y2=1.915
r169 68 85 11.7546 $w=5.78e-07 $l=5.7e-07 $layer=LI1_cond $X=5.495 $Y=1.915
+ $X2=6.065 $Y2=1.915
r170 68 69 1.08702 $w=5.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.495 $Y=1.915
+ $X2=5.33 $Y2=1.915
r171 63 72 4.69387 $w=6.5e-07 $l=3.04631e-07 $layer=LI1_cond $X=8.655 $Y=1.625
+ $X2=8.625 $Y2=1.915
r172 63 65 12.636 $w=6.18e-07 $l=6.55e-07 $layer=LI1_cond $X=8.655 $Y=1.625
+ $X2=8.655 $Y2=0.97
r173 60 74 8.67899 $w=6.8e-07 $l=4.7e-07 $layer=LI1_cond $X=8.625 $Y=2.89
+ $X2=8.625 $Y2=3.36
r174 60 62 9.67416 $w=6.78e-07 $l=5.5e-07 $layer=LI1_cond $X=8.625 $Y=2.89
+ $X2=8.625 $Y2=2.34
r175 59 72 4.69387 $w=6.5e-07 $l=2.9e-07 $layer=LI1_cond $X=8.625 $Y=2.205
+ $X2=8.625 $Y2=1.915
r176 59 62 2.37457 $w=6.78e-07 $l=1.35e-07 $layer=LI1_cond $X=8.625 $Y=2.205
+ $X2=8.625 $Y2=2.34
r177 58 71 1.08702 $w=5.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.055 $Y=1.915
+ $X2=6.89 $Y2=1.915
r178 57 72 1.75591 $w=5.8e-07 $l=3.4e-07 $layer=LI1_cond $X=8.285 $Y=1.915
+ $X2=8.625 $Y2=1.915
r179 57 58 25.3651 $w=5.78e-07 $l=1.23e-06 $layer=LI1_cond $X=8.285 $Y=1.915
+ $X2=7.055 $Y2=1.915
r180 53 71 5.63874 $w=2.1e-07 $l=2.9e-07 $layer=LI1_cond $X=6.89 $Y=1.625
+ $X2=6.89 $Y2=1.915
r181 53 55 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=6.89 $Y=1.625
+ $X2=6.89 $Y2=0.97
r182 49 51 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=6.89 $Y=2.34
+ $X2=6.89 $Y2=3.36
r183 47 71 5.63874 $w=3.3e-07 $l=2.9e-07 $layer=LI1_cond $X=6.89 $Y=2.205
+ $X2=6.89 $Y2=1.915
r184 47 49 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.89 $Y=2.205
+ $X2=6.89 $Y2=2.34
r185 43 69 5.63874 $w=2.1e-07 $l=2.9e-07 $layer=LI1_cond $X=5.33 $Y=1.625
+ $X2=5.33 $Y2=1.915
r186 43 45 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=5.33 $Y=1.625
+ $X2=5.33 $Y2=0.97
r187 39 41 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=5.33 $Y=2.34
+ $X2=5.33 $Y2=3.36
r188 37 69 5.63874 $w=3.3e-07 $l=2.9e-07 $layer=LI1_cond $X=5.33 $Y=2.205
+ $X2=5.33 $Y2=1.915
r189 37 39 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.33 $Y=2.205
+ $X2=5.33 $Y2=2.34
r190 36 67 1.2027 $w=5.8e-07 $l=3.49428e-07 $layer=LI1_cond $X=3.935 $Y=1.915
+ $X2=3.605 $Y2=1.955
r191 35 69 1.08702 $w=5.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=1.915
+ $X2=5.33 $Y2=1.915
r192 35 36 25.3651 $w=5.78e-07 $l=1.23e-06 $layer=LI1_cond $X=5.165 $Y=1.915
+ $X2=3.935 $Y2=1.915
r193 31 67 9.23321 $w=2.7e-07 $l=4.04166e-07 $layer=LI1_cond $X=3.77 $Y=1.625
+ $X2=3.605 $Y2=1.955
r194 31 33 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=3.77 $Y=1.625
+ $X2=3.77 $Y2=0.97
r195 27 29 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3.77 $Y=2.34
+ $X2=3.77 $Y2=3.36
r196 25 67 9.23321 $w=2.7e-07 $l=3.22102e-07 $layer=LI1_cond $X=3.77 $Y=2.205
+ $X2=3.605 $Y2=1.955
r197 25 27 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.77 $Y=2.205
+ $X2=3.77 $Y2=2.34
r198 8 74 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=8.31
+ $Y=2.215 $X2=8.45 $Y2=3.36
r199 8 62 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=8.31
+ $Y=2.215 $X2=8.45 $Y2=2.34
r200 7 51 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=6.75
+ $Y=2.215 $X2=6.89 $Y2=3.36
r201 7 49 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=6.75
+ $Y=2.215 $X2=6.89 $Y2=2.34
r202 6 41 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=5.19
+ $Y=2.215 $X2=5.33 $Y2=3.36
r203 6 39 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=5.19
+ $Y=2.215 $X2=5.33 $Y2=2.34
r204 5 29 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=3.63
+ $Y=2.215 $X2=3.77 $Y2=3.36
r205 5 27 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=3.63
+ $Y=2.215 $X2=3.77 $Y2=2.34
r206 4 65 91 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=2 $X=8.31
+ $Y=0.705 $X2=8.45 $Y2=0.97
r207 3 55 91 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=2 $X=6.75
+ $Y=0.705 $X2=6.89 $Y2=0.97
r208 2 45 91 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=2 $X=5.19
+ $Y=0.705 $X2=5.33 $Y2=0.97
r209 1 33 91 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=2 $X=3.63
+ $Y=0.705 $X2=3.77 $Y2=0.97
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBEC_P_8%VGND 1 2 3 4 5 6 19 31 33 56 58 67 73 77
+ 83 87 93 95 97 102 103 105 118
c123 97 0 1.2129e-19 $X=9.42 $Y=0.465
r124 103 108 0.16865 $w=2.8e-07 $l=3.2e-07 $layer=MET2_cond $X=9.76 $Y=0.425
+ $X2=9.44 $Y2=0.425
r125 102 103 4.5 $w=1.5e-07 $l=1.5e-07 $layer=via $count=1 $X=9.76 $Y=0.435
+ $X2=9.76 $Y2=0.435
r126 93 95 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=8.175 $Y=0.465
+ $X2=8.975 $Y2=0.465
r127 92 105 0.52787 $w=3.7e-07 $l=1.375e-06 $layer=MET1_cond $X=8.04 $Y=0.44
+ $X2=9.415 $Y2=0.44
r128 91 93 12.8638 $w=1.063e-06 $l=1.35e-07 $layer=LI1_cond $X=8.04 $Y=0.912
+ $X2=8.175 $Y2=0.912
r129 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.04 $Y=0.465
+ $X2=8.04 $Y2=0.465
r130 89 91 4.2385 $w=1.063e-06 $l=3.7e-07 $layer=LI1_cond $X=7.67 $Y=0.912
+ $X2=8.04 $Y2=0.912
r131 86 92 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.32 $Y=0.44
+ $X2=8.04 $Y2=0.44
r132 85 89 4.00939 $w=1.063e-06 $l=3.5e-07 $layer=LI1_cond $X=7.32 $Y=0.912
+ $X2=7.67 $Y2=0.912
r133 85 87 13.0929 $w=1.063e-06 $l=1.55e-07 $layer=LI1_cond $X=7.32 $Y=0.912
+ $X2=7.165 $Y2=0.912
r134 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.32 $Y=0.465
+ $X2=7.32 $Y2=0.465
r135 83 87 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.615 $Y=0.465
+ $X2=7.165 $Y2=0.465
r136 82 86 0.3244 $w=3.7e-07 $l=8.45e-07 $layer=MET1_cond $X=6.475 $Y=0.44
+ $X2=7.32 $Y2=0.44
r137 81 83 12.9211 $w=1.063e-06 $l=1.4e-07 $layer=LI1_cond $X=6.475 $Y=0.912
+ $X2=6.615 $Y2=0.912
r138 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.475 $Y=0.465
+ $X2=6.475 $Y2=0.465
r139 79 81 4.18122 $w=1.063e-06 $l=3.65e-07 $layer=LI1_cond $X=6.11 $Y=0.912
+ $X2=6.475 $Y2=0.912
r140 76 82 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.755 $Y=0.44
+ $X2=6.475 $Y2=0.44
r141 76 118 0.36663 $w=3.7e-07 $l=9.55e-07 $layer=MET1_cond $X=5.755 $Y=0.44
+ $X2=4.8 $Y2=0.44
r142 75 79 4.06667 $w=1.063e-06 $l=3.55e-07 $layer=LI1_cond $X=5.755 $Y=0.912
+ $X2=6.11 $Y2=0.912
r143 75 77 13.0357 $w=1.063e-06 $l=1.5e-07 $layer=LI1_cond $X=5.755 $Y=0.912
+ $X2=5.605 $Y2=0.912
r144 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.755 $Y=0.465
+ $X2=5.755 $Y2=0.465
r145 73 77 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.055 $Y=0.465
+ $X2=5.605 $Y2=0.465
r146 71 73 13.3793 $w=1.063e-06 $l=1.8e-07 $layer=LI1_cond $X=4.875 $Y=0.912
+ $X2=5.055 $Y2=0.912
r147 71 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.875 $Y=0.465
+ $X2=4.875 $Y2=0.465
r148 69 71 3.723 $w=1.063e-06 $l=3.25e-07 $layer=LI1_cond $X=4.55 $Y=0.912
+ $X2=4.875 $Y2=0.912
r149 65 69 4.52488 $w=1.063e-06 $l=3.95e-07 $layer=LI1_cond $X=4.155 $Y=0.912
+ $X2=4.55 $Y2=0.912
r150 65 67 12.5774 $w=1.063e-06 $l=1.1e-07 $layer=LI1_cond $X=4.155 $Y=0.912
+ $X2=4.045 $Y2=0.912
r151 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.155 $Y=0.465
+ $X2=4.155 $Y2=0.465
r152 61 66 0.28601 $w=3.7e-07 $l=7.45e-07 $layer=MET1_cond $X=3.41 $Y=0.44
+ $X2=4.155 $Y2=0.44
r153 59 61 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.69 $Y=0.44
+ $X2=3.41 $Y2=0.44
r154 58 63 7.36341 $w=7.87e-07 $l=4.75e-07 $layer=LI1_cond $X=3.05 $Y=0.465
+ $X2=3.05 $Y2=0.94
r155 58 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.41 $Y=0.465
+ $X2=3.41 $Y2=0.465
r156 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.69 $Y=0.465
+ $X2=2.69 $Y2=0.465
r157 55 59 0.32632 $w=3.7e-07 $l=8.5e-07 $layer=MET1_cond $X=1.84 $Y=0.44
+ $X2=2.69 $Y2=0.44
r158 54 56 11.907 $w=1.003e-06 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=0.882
+ $X2=1.925 $Y2=0.882
r159 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.84 $Y=0.465
+ $X2=1.84 $Y2=0.465
r160 52 54 7.64776 $w=1.003e-06 $l=6.3e-07 $layer=LI1_cond $X=1.21 $Y=0.882
+ $X2=1.84 $Y2=0.882
r161 49 55 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=0.76 $Y=0.44
+ $X2=1.84 $Y2=0.44
r162 48 52 5.46269 $w=1.003e-06 $l=4.5e-07 $layer=LI1_cond $X=0.76 $Y=0.882
+ $X2=1.21 $Y2=0.882
r163 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.76 $Y=0.465
+ $X2=0.76 $Y2=0.465
r164 33 118 0.0357032 $w=3.7e-07 $l=9.3e-08 $layer=MET1_cond $X=4.707 $Y=0.44
+ $X2=4.8 $Y2=0.44
r165 33 66 0.211916 $w=3.7e-07 $l=5.52e-07 $layer=MET1_cond $X=4.707 $Y=0.44
+ $X2=4.155 $Y2=0.44
r166 33 108 4.5 $w=1.5e-07 $l=1.5e-07 $layer=via $count=1 $X=9.44 $Y=0.435
+ $X2=9.44 $Y2=0.435
r167 33 105 0.00191953 $w=3.7e-07 $l=5e-09 $layer=MET1_cond $X=9.42 $Y=0.44
+ $X2=9.415 $Y2=0.44
r168 33 102 0.0761468 $w=5.2e-07 $l=1.6e-07 $layer=MET1_cond $X=9.6 $Y=0.435
+ $X2=9.76 $Y2=0.435
r169 33 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.42 $Y=0.465
+ $X2=9.42 $Y2=0.465
r170 29 97 5.23838 $w=2.18e-07 $l=1e-07 $layer=LI1_cond $X=9.32 $Y=0.49 $X2=9.42
+ $Y2=0.49
r171 29 95 18.6977 $w=2.18e-07 $l=3.45e-07 $layer=LI1_cond $X=9.32 $Y=0.49
+ $X2=8.975 $Y2=0.49
r172 29 31 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.32 $Y=0.6 $X2=9.32
+ $Y2=0.94
r173 22 58 10.0992 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=3.495 $Y=0.465
+ $X2=3.05 $Y2=0.465
r174 22 67 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.495 $Y=0.465
+ $X2=4.045 $Y2=0.465
r175 19 58 10.0992 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=2.605 $Y=0.465
+ $X2=3.05 $Y2=0.465
r176 19 56 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.605 $Y=0.465
+ $X2=1.925 $Y2=0.465
r177 6 31 91 $w=1.7e-07 $l=3.04672e-07 $layer=licon1_NDIFF $count=2 $X=9.09
+ $Y=0.705 $X2=9.25 $Y2=0.94
r178 5 89 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=7.53
+ $Y=0.705 $X2=7.67 $Y2=0.94
r179 4 79 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=5.97
+ $Y=0.705 $X2=6.11 $Y2=0.94
r180 3 69 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=4.41
+ $Y=0.705 $X2=4.55 $Y2=0.94
r181 2 63 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.705 $X2=2.99 $Y2=0.94
r182 1 52 91 $w=1.7e-07 $l=3.1229e-07 $layer=licon1_NDIFF $count=2 $X=1.03
+ $Y=0.705 $X2=1.21 $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBEC_P_8%X 1 4 8 10
c64 10 0 3.69313e-19 $X=4.16 $Y=2.035
c65 4 0 1.43567e-19 $X=3 $Y=2.035
r66 5 10 0.0218943 $w=1.6e-06 $l=1.16e-06 $layer=MET5_cond $X=3 $Y=2.035
+ $X2=4.16 $Y2=2.035
r67 4 8 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=3.425 $Y=2.035
+ $X2=3.425 $Y2=2.035
r68 4 5 0.38 $w=8e-07 $l=8e-07 $layer=via4_notcap2m $count=1 $X=3 $Y=2.035 $X2=3
+ $Y2=2.035
r69 1 8 0.0552787 $w=3.2e-07 $l=3.45e-07 $layer=MET3_cond $X=3.08 $Y=2.035
+ $X2=3.425 $Y2=2.035
.ends

