* File: sky130_fd_sc_hvl__dfrtp_1.pxi.spice
* Created: Wed Sep  2 09:05:05 2020
* 
x_PM_SKY130_FD_SC_HVL__DFRTP_1%VNB N_VNB_M1016_b VNB N_VNB_c_3_p
+ PM_SKY130_FD_SC_HVL__DFRTP_1%VNB
x_PM_SKY130_FD_SC_HVL__DFRTP_1%VPB N_VPB_M1018_b VPB N_VPB_c_101_p
+ PM_SKY130_FD_SC_HVL__DFRTP_1%VPB
x_PM_SKY130_FD_SC_HVL__DFRTP_1%CLK N_CLK_M1018_g N_CLK_M1016_g CLK CLK CLK
+ N_CLK_c_264_n PM_SKY130_FD_SC_HVL__DFRTP_1%CLK
x_PM_SKY130_FD_SC_HVL__DFRTP_1%A_30_107# N_A_30_107#_M1016_s N_A_30_107#_M1018_s
+ N_A_30_107#_M1000_g N_A_30_107#_M1028_g N_A_30_107#_c_307_n
+ N_A_30_107#_M1008_g N_A_30_107#_c_309_n N_A_30_107#_M1007_g
+ N_A_30_107#_c_294_n N_A_30_107#_M1030_g N_A_30_107#_c_295_n
+ N_A_30_107#_c_296_n N_A_30_107#_c_313_n N_A_30_107#_c_316_n
+ N_A_30_107#_c_356_n N_A_30_107#_c_298_n N_A_30_107#_c_318_n
+ N_A_30_107#_c_319_n N_A_30_107#_c_322_n N_A_30_107#_c_364_p
+ N_A_30_107#_c_325_n N_A_30_107#_c_366_p N_A_30_107#_c_367_p
+ N_A_30_107#_c_326_n N_A_30_107#_c_329_n N_A_30_107#_c_450_p
+ N_A_30_107#_c_412_p N_A_30_107#_c_332_n N_A_30_107#_c_369_p
+ N_A_30_107#_c_333_n N_A_30_107#_c_336_n N_A_30_107#_c_339_n
+ N_A_30_107#_c_340_n N_A_30_107#_c_341_n N_A_30_107#_c_299_n
+ N_A_30_107#_c_300_n N_A_30_107#_c_301_n N_A_30_107#_c_302_n
+ N_A_30_107#_c_386_p N_A_30_107#_c_303_n N_A_30_107#_c_343_n
+ N_A_30_107#_c_404_p N_A_30_107#_c_344_n N_A_30_107#_M1013_g
+ PM_SKY130_FD_SC_HVL__DFRTP_1%A_30_107#
x_PM_SKY130_FD_SC_HVL__DFRTP_1%RESET_B N_RESET_B_M1024_g N_RESET_B_M1012_g
+ N_RESET_B_M1029_g N_RESET_B_c_598_n N_RESET_B_M1006_g N_RESET_B_M1005_g
+ N_RESET_B_M1011_g N_RESET_B_c_603_n N_RESET_B_c_576_n N_RESET_B_c_578_n
+ N_RESET_B_c_580_n N_RESET_B_c_581_n N_RESET_B_c_658_p N_RESET_B_c_582_n
+ N_RESET_B_c_583_n N_RESET_B_c_631_p N_RESET_B_c_669_p N_RESET_B_c_584_n
+ N_RESET_B_c_586_n N_RESET_B_c_622_n N_RESET_B_c_588_n N_RESET_B_c_696_p
+ N_RESET_B_c_589_n N_RESET_B_c_590_n N_RESET_B_c_591_n N_RESET_B_c_667_p
+ N_RESET_B_c_697_p N_RESET_B_c_592_n RESET_B N_RESET_B_c_593_n
+ N_RESET_B_c_594_n PM_SKY130_FD_SC_HVL__DFRTP_1%RESET_B
x_PM_SKY130_FD_SC_HVL__DFRTP_1%D N_D_M1009_g N_D_c_767_n D D D N_D_M1014_g
+ PM_SKY130_FD_SC_HVL__DFRTP_1%D
x_PM_SKY130_FD_SC_HVL__DFRTP_1%A_339_537# N_A_339_537#_M1028_d
+ N_A_339_537#_M1000_d N_A_339_537#_c_804_n N_A_339_537#_M1017_g
+ N_A_339_537#_M1027_g N_A_339_537#_c_805_n N_A_339_537#_c_806_n
+ N_A_339_537#_c_808_n N_A_339_537#_c_814_n N_A_339_537#_c_850_n
+ N_A_339_537#_c_809_n N_A_339_537#_c_815_n N_A_339_537#_c_816_n
+ N_A_339_537#_c_818_n N_A_339_537#_c_860_n N_A_339_537#_c_819_n
+ N_A_339_537#_c_820_n N_A_339_537#_c_821_n N_A_339_537#_c_822_n
+ N_A_339_537#_c_823_n N_A_339_537#_c_824_n N_A_339_537#_c_825_n
+ N_A_339_537#_c_826_n N_A_339_537#_M1001_g N_A_339_537#_M1020_g
+ N_A_339_537#_c_828_n N_A_339_537#_c_811_n
+ PM_SKY130_FD_SC_HVL__DFRTP_1%A_339_537#
x_PM_SKY130_FD_SC_HVL__DFRTP_1%A_1119_506# N_A_1119_506#_M1004_d
+ N_A_1119_506#_M1022_d N_A_1119_506#_M1026_g N_A_1119_506#_M1003_g
+ N_A_1119_506#_c_1010_n N_A_1119_506#_c_1002_n N_A_1119_506#_c_1003_n
+ N_A_1119_506#_c_1042_n N_A_1119_506#_c_1004_n N_A_1119_506#_c_1012_n
+ N_A_1119_506#_c_1074_p N_A_1119_506#_c_1023_n N_A_1119_506#_c_1048_n
+ N_A_1119_506#_c_1005_n N_A_1119_506#_c_1030_n N_A_1119_506#_c_1006_n
+ PM_SKY130_FD_SC_HVL__DFRTP_1%A_1119_506#
x_PM_SKY130_FD_SC_HVL__DFRTP_1%A_921_632# N_A_921_632#_M1008_d
+ N_A_921_632#_M1001_d N_A_921_632#_M1006_d N_A_921_632#_M1022_g
+ N_A_921_632#_c_1097_n N_A_921_632#_M1004_g N_A_921_632#_c_1108_n
+ N_A_921_632#_c_1109_n N_A_921_632#_c_1154_n N_A_921_632#_c_1099_n
+ N_A_921_632#_c_1100_n N_A_921_632#_c_1101_n N_A_921_632#_c_1111_n
+ N_A_921_632#_c_1112_n N_A_921_632#_c_1132_n N_A_921_632#_c_1113_n
+ N_A_921_632#_c_1102_n N_A_921_632#_c_1103_n N_A_921_632#_c_1114_n
+ N_A_921_632#_c_1104_n PM_SKY130_FD_SC_HVL__DFRTP_1%A_921_632#
x_PM_SKY130_FD_SC_HVL__DFRTP_1%A_2096_417# N_A_2096_417#_M1023_d
+ N_A_2096_417#_M1005_d N_A_2096_417#_M1021_g N_A_2096_417#_c_1242_n
+ N_A_2096_417#_c_1249_n N_A_2096_417#_c_1234_n N_A_2096_417#_c_1293_p
+ N_A_2096_417#_c_1244_n N_A_2096_417#_c_1245_n N_A_2096_417#_c_1246_n
+ N_A_2096_417#_c_1235_n N_A_2096_417#_c_1237_n N_A_2096_417#_c_1247_n
+ N_A_2096_417#_c_1238_n N_A_2096_417#_c_1282_p N_A_2096_417#_M1031_g
+ PM_SKY130_FD_SC_HVL__DFRTP_1%A_2096_417#
x_PM_SKY130_FD_SC_HVL__DFRTP_1%A_1875_543# N_A_1875_543#_M1017_d
+ N_A_1875_543#_M1007_d N_A_1875_543#_M1023_g N_A_1875_543#_c_1324_n
+ N_A_1875_543#_M1015_g N_A_1875_543#_M1019_g N_A_1875_543#_c_1326_n
+ N_A_1875_543#_c_1327_n N_A_1875_543#_c_1364_n N_A_1875_543#_c_1328_n
+ N_A_1875_543#_c_1334_n N_A_1875_543#_c_1335_n N_A_1875_543#_c_1338_n
+ N_A_1875_543#_c_1351_n N_A_1875_543#_c_1339_n N_A_1875_543#_c_1329_n
+ N_A_1875_543#_c_1341_n N_A_1875_543#_c_1342_n N_A_1875_543#_c_1343_n
+ N_A_1875_543#_M1025_g PM_SKY130_FD_SC_HVL__DFRTP_1%A_1875_543#
x_PM_SKY130_FD_SC_HVL__DFRTP_1%A_2649_207# N_A_2649_207#_M1015_s
+ N_A_2649_207#_M1019_s N_A_2649_207#_M1002_g N_A_2649_207#_M1010_g
+ N_A_2649_207#_c_1457_n N_A_2649_207#_c_1458_n N_A_2649_207#_c_1465_n
+ N_A_2649_207#_c_1459_n N_A_2649_207#_c_1460_n N_A_2649_207#_c_1461_n
+ N_A_2649_207#_c_1472_n PM_SKY130_FD_SC_HVL__DFRTP_1%A_2649_207#
x_PM_SKY130_FD_SC_HVL__DFRTP_1%VPWR N_VPWR_M1018_d N_VPWR_M1024_d N_VPWR_M1026_d
+ N_VPWR_M1022_s N_VPWR_M1021_d N_VPWR_M1025_d N_VPWR_M1019_d VPWR
+ N_VPWR_c_1507_n N_VPWR_c_1510_n N_VPWR_c_1513_n N_VPWR_c_1516_n
+ N_VPWR_c_1519_n N_VPWR_c_1522_n N_VPWR_c_1525_n N_VPWR_c_1528_n
+ PM_SKY130_FD_SC_HVL__DFRTP_1%VPWR
x_PM_SKY130_FD_SC_HVL__DFRTP_1%A_452_632# N_A_452_632#_M1014_d
+ N_A_452_632#_M1024_s N_A_452_632#_M1009_d N_A_452_632#_c_1634_n
+ N_A_452_632#_c_1635_n N_A_452_632#_c_1636_n N_A_452_632#_c_1637_n
+ N_A_452_632#_c_1638_n N_A_452_632#_c_1631_n N_A_452_632#_c_1632_n
+ N_A_452_632#_c_1640_n N_A_452_632#_c_1641_n N_A_452_632#_c_1633_n
+ PM_SKY130_FD_SC_HVL__DFRTP_1%A_452_632#
x_PM_SKY130_FD_SC_HVL__DFRTP_1%Q N_Q_M1002_d N_Q_M1010_d Q Q Q Q Q Q Q
+ N_Q_c_1696_n PM_SKY130_FD_SC_HVL__DFRTP_1%Q
x_PM_SKY130_FD_SC_HVL__DFRTP_1%VGND N_VGND_M1016_d N_VGND_M1012_s N_VGND_M1029_d
+ N_VGND_M1031_d N_VGND_M1015_d VGND N_VGND_c_1708_n N_VGND_c_1710_n
+ N_VGND_c_1712_n N_VGND_c_1714_n N_VGND_c_1716_n N_VGND_c_1718_n
+ PM_SKY130_FD_SC_HVL__DFRTP_1%VGND
cc_1 N_VNB_M1016_b N_CLK_M1018_g 0.00183817f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=3.06
cc_2 N_VNB_M1016_b N_CLK_M1016_g 0.04492f $X=-0.33 $Y=-0.265 $X2=0.685 $Y2=0.745
cc_3 N_VNB_c_3_p N_CLK_M1016_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.685 $Y2=0.745
cc_4 N_VNB_M1016_b N_CLK_c_264_n 0.0787707f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=1.34
cc_5 N_VNB_M1016_b N_A_30_107#_M1028_g 0.11909f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_c_3_p N_A_30_107#_M1028_g 9.58849e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_7 N_VNB_M1016_b N_A_30_107#_M1008_g 0.0792881f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=1.34
cc_8 N_VNB_M1016_b N_A_30_107#_c_294_n 0.0274493f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_M1016_b N_A_30_107#_c_295_n 0.0212608f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_10 N_VNB_M1016_b N_A_30_107#_c_296_n 0.0734121f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_c_3_p N_A_30_107#_c_296_n 6.28066e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_12 N_VNB_M1016_b N_A_30_107#_c_298_n 0.00603047f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1016_b N_A_30_107#_c_299_n 0.00191258f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_M1016_b N_A_30_107#_c_300_n 0.009108f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_15 N_VNB_M1016_b N_A_30_107#_c_301_n 0.0103681f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_16 N_VNB_M1016_b N_A_30_107#_c_302_n 7.13236e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_17 N_VNB_M1016_b N_A_30_107#_c_303_n 0.0588414f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1016_b N_RESET_B_M1029_g 0.0898229f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.58
cc_19 N_VNB_M1016_b N_RESET_B_M1005_g 0.010911f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=1.295
cc_20 N_VNB_M1016_b N_RESET_B_c_576_n 0.149549f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_21 N_VNB_c_3_p N_RESET_B_c_576_n 0.00699185f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_22 N_VNB_M1016_b N_RESET_B_c_578_n 0.00794781f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_23 N_VNB_c_3_p N_RESET_B_c_578_n 4.18973e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_24 N_VNB_M1016_b N_RESET_B_c_580_n 0.00714554f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_25 N_VNB_M1016_b N_RESET_B_c_581_n 0.012826f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_26 N_VNB_M1016_b N_RESET_B_c_582_n 0.00851024f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_27 N_VNB_M1016_b N_RESET_B_c_583_n 0.0206369f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_28 N_VNB_M1016_b N_RESET_B_c_584_n 0.179338f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_29 N_VNB_c_3_p N_RESET_B_c_584_n 0.00840003f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_30 N_VNB_M1016_b N_RESET_B_c_586_n 0.0135577f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_31 N_VNB_c_3_p N_RESET_B_c_586_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_32 N_VNB_M1016_b N_RESET_B_c_588_n 0.00506015f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_33 N_VNB_M1016_b N_RESET_B_c_589_n 0.00164515f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_34 N_VNB_M1016_b N_RESET_B_c_590_n 0.0581971f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_35 N_VNB_M1016_b N_RESET_B_c_591_n 0.00778724f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_36 N_VNB_M1016_b N_RESET_B_c_592_n 0.0675542f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_37 N_VNB_M1016_b N_RESET_B_c_593_n 0.0453905f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_38 N_VNB_M1016_b N_RESET_B_c_594_n 0.0364404f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_39 N_VNB_M1016_b N_D_M1014_g 0.0778363f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_40 N_VNB_M1016_b N_A_339_537#_c_804_n 0.0382086f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=0.745
cc_41 N_VNB_M1016_b N_A_339_537#_c_805_n 0.049762f $X=-0.33 $Y=-0.265 $X2=0.675
+ $Y2=1.085
cc_42 N_VNB_M1016_b N_A_339_537#_c_806_n 0.0138837f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_c_3_p N_A_339_537#_c_806_n 8.16848e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_44 N_VNB_M1016_b N_A_339_537#_c_808_n 0.0269863f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=2.035
cc_45 N_VNB_M1016_b N_A_339_537#_c_809_n 0.00295213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_M1016_b N_A_339_537#_M1020_g 0.077847f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_47 N_VNB_M1016_b N_A_339_537#_c_811_n 0.0160658f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_M1016_b N_A_1119_506#_c_1002_n 0.0217779f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=1.34
cc_49 N_VNB_M1016_b N_A_1119_506#_c_1003_n 0.0396957f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=1.085
cc_50 N_VNB_M1016_b N_A_1119_506#_c_1004_n 0.0202923f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_51 N_VNB_M1016_b N_A_1119_506#_c_1005_n 0.00487839f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_52 N_VNB_M1016_b N_A_1119_506#_c_1006_n 7.12344e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_53 N_VNB_M1016_b N_A_921_632#_c_1097_n 0.045275f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_54 N_VNB_c_3_p N_A_921_632#_c_1097_n 5.98017e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_55 N_VNB_M1016_b N_A_921_632#_c_1099_n 0.00321392f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_56 N_VNB_M1016_b N_A_921_632#_c_1100_n 0.00375955f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_57 N_VNB_M1016_b N_A_921_632#_c_1101_n 0.0225307f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_58 N_VNB_M1016_b N_A_921_632#_c_1102_n 0.00223884f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_59 N_VNB_M1016_b N_A_921_632#_c_1103_n 0.00102919f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_60 N_VNB_M1016_b N_A_921_632#_c_1104_n 0.0876728f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_61 N_VNB_M1016_b N_A_2096_417#_c_1234_n 0.0111045f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=1.865
cc_62 N_VNB_M1016_b N_A_2096_417#_c_1235_n 0.0208938f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_63 N_VNB_c_3_p N_A_2096_417#_c_1235_n 8.21372e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_64 N_VNB_M1016_b N_A_2096_417#_c_1237_n 0.00657723f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_65 N_VNB_M1016_b N_A_2096_417#_c_1238_n 0.00605718f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_66 N_VNB_M1016_b N_A_2096_417#_M1031_g 0.111026f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_67 N_VNB_c_3_p N_A_2096_417#_M1031_g 8.54021e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_68 N_VNB_M1016_b N_A_1875_543#_M1023_g 0.102697f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.21
cc_69 N_VNB_c_3_p N_A_1875_543#_M1023_g 0.0023273f $X=0.24 $Y=0 $X2=0.635
+ $Y2=1.21
cc_70 N_VNB_M1016_b N_A_1875_543#_c_1324_n 0.0550779f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=1.95
cc_71 N_VNB_M1016_b N_A_1875_543#_M1015_g 0.0430857f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=1.34
cc_72 N_VNB_M1016_b N_A_1875_543#_c_1326_n 0.021099f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_73 N_VNB_M1016_b N_A_1875_543#_c_1327_n 0.0230454f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=1.665
cc_74 N_VNB_M1016_b N_A_1875_543#_c_1328_n 0.00526301f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_75 N_VNB_M1016_b N_A_1875_543#_c_1329_n 0.00778568f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_76 N_VNB_M1016_b N_A_2649_207#_M1002_g 0.0492564f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=1.21
cc_77 N_VNB_c_3_p N_A_2649_207#_M1002_g 9.28887e-19 $X=0.24 $Y=0 $X2=0.635
+ $Y2=1.21
cc_78 N_VNB_M1016_b N_A_2649_207#_c_1457_n 0.00863758f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=1.34
cc_79 N_VNB_M1016_b N_A_2649_207#_c_1458_n 0.00129586f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=1.295
cc_80 N_VNB_M1016_b N_A_2649_207#_c_1459_n 0.0028368f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_81 N_VNB_M1016_b N_A_2649_207#_c_1460_n 0.0336135f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_82 N_VNB_M1016_b N_A_2649_207#_c_1461_n 0.00296628f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_83 N_VNB_M1016_b N_A_452_632#_c_1631_n 0.00229087f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_84 N_VNB_M1016_b N_A_452_632#_c_1632_n 0.0112012f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_85 N_VNB_M1016_b N_A_452_632#_c_1633_n 0.003269f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_86 N_VNB_M1016_b N_Q_c_1696_n 0.0565391f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_87 N_VNB_M1016_b N_VGND_c_1708_n 0.058257f $X=-0.33 $Y=-0.265 $X2=0.675
+ $Y2=1.865
cc_88 N_VNB_c_3_p N_VGND_c_1708_n 0.00269373f $X=0.24 $Y=0 $X2=0.675 $Y2=1.865
cc_89 N_VNB_M1016_b N_VGND_c_1710_n 0.0553697f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_90 N_VNB_c_3_p N_VGND_c_1710_n 0.00166879f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_91 N_VNB_M1016_b N_VGND_c_1712_n 0.0695943f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_92 N_VNB_c_3_p N_VGND_c_1712_n 0.002699f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_93 N_VNB_M1016_b N_VGND_c_1714_n 0.0479288f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_94 N_VNB_c_3_p N_VGND_c_1714_n 0.00270129f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_95 N_VNB_M1016_b N_VGND_c_1716_n 0.0741524f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_96 N_VNB_c_3_p N_VGND_c_1716_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_97 N_VNB_M1016_b N_VGND_c_1718_n 0.243951f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_98 N_VNB_c_3_p N_VGND_c_1718_n 1.64226f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_99 N_VPB_M1018_b N_CLK_M1018_g 0.106066f $X=-0.33 $Y=1.885 $X2=0.665 $Y2=3.06
cc_100 VPB N_CLK_M1018_g 8.9764e-19 $X=0 $Y=3.955 $X2=0.665 $Y2=3.06
cc_101 N_VPB_c_101_p N_CLK_M1018_g 0.00515583f $X=15.12 $Y=4.07 $X2=0.665
+ $Y2=3.06
cc_102 N_VPB_M1018_b N_A_30_107#_M1000_g 0.0413251f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.21
cc_103 VPB N_A_30_107#_M1000_g 7.58639e-19 $X=0 $Y=3.955 $X2=0.635 $Y2=1.21
cc_104 N_VPB_c_101_p N_A_30_107#_M1000_g 0.00432362f $X=15.12 $Y=4.07 $X2=0.635
+ $Y2=1.21
cc_105 N_VPB_M1018_b N_A_30_107#_c_307_n 0.105413f $X=-0.33 $Y=1.885 $X2=0.675
+ $Y2=1.34
cc_106 N_VPB_M1018_b N_A_30_107#_M1008_g 0.0158199f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=1.34
cc_107 N_VPB_M1018_b N_A_30_107#_c_309_n 0.040306f $X=-0.33 $Y=1.885 $X2=0.675
+ $Y2=1.865
cc_108 VPB N_A_30_107#_c_309_n 0.00970178f $X=0 $Y=3.955 $X2=0.675 $Y2=1.865
cc_109 N_VPB_c_101_p N_A_30_107#_c_309_n 0.0196751f $X=15.12 $Y=4.07 $X2=0.675
+ $Y2=1.865
cc_110 N_VPB_M1018_b N_A_30_107#_c_296_n 0.0242711f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_111 N_VPB_M1018_b N_A_30_107#_c_313_n 0.0387844f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_112 VPB N_A_30_107#_c_313_n 7.0347e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_113 N_VPB_c_101_p N_A_30_107#_c_313_n 0.00639736f $X=15.12 $Y=4.07 $X2=0
+ $Y2=0
cc_114 N_VPB_M1018_b N_A_30_107#_c_316_n 0.0119027f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_115 N_VPB_M1018_b N_A_30_107#_c_298_n 0.0663276f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_116 N_VPB_M1018_b N_A_30_107#_c_318_n 0.00113164f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_117 N_VPB_M1018_b N_A_30_107#_c_319_n 0.0178951f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_118 VPB N_A_30_107#_c_319_n 0.00428557f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_119 N_VPB_c_101_p N_A_30_107#_c_319_n 0.0837795f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_120 N_VPB_M1018_b N_A_30_107#_c_322_n 0.00252874f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_121 VPB N_A_30_107#_c_322_n 5.70856e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_122 N_VPB_c_101_p N_A_30_107#_c_322_n 0.0114989f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_123 N_VPB_M1018_b N_A_30_107#_c_325_n 0.00262232f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_124 N_VPB_M1018_b N_A_30_107#_c_326_n 0.00989982f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_125 VPB N_A_30_107#_c_326_n 0.00529907f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_126 N_VPB_c_101_p N_A_30_107#_c_326_n 0.103511f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_127 N_VPB_M1018_b N_A_30_107#_c_329_n 0.00183475f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_128 VPB N_A_30_107#_c_329_n 5.70856e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_129 N_VPB_c_101_p N_A_30_107#_c_329_n 0.0114989f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_130 N_VPB_M1018_b N_A_30_107#_c_332_n 0.00975788f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_131 N_VPB_M1018_b N_A_30_107#_c_333_n 0.0105162f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_132 VPB N_A_30_107#_c_333_n 0.00290029f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_133 N_VPB_c_101_p N_A_30_107#_c_333_n 0.0568193f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_134 N_VPB_M1018_b N_A_30_107#_c_336_n 0.00183475f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_135 VPB N_A_30_107#_c_336_n 5.70856e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_136 N_VPB_c_101_p N_A_30_107#_c_336_n 0.0114989f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_137 N_VPB_M1018_b N_A_30_107#_c_339_n 0.00869251f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_138 N_VPB_M1018_b N_A_30_107#_c_340_n 0.0101952f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_139 N_VPB_M1018_b N_A_30_107#_c_341_n 0.00927491f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_140 N_VPB_M1018_b N_A_30_107#_c_300_n 0.0552152f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_141 N_VPB_M1018_b N_A_30_107#_c_343_n 0.0091351f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_142 N_VPB_M1018_b N_A_30_107#_c_344_n 0.0675017f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_143 VPB N_A_30_107#_c_344_n 5.81702e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_144 N_VPB_c_101_p N_A_30_107#_c_344_n 0.00477198f $X=15.12 $Y=4.07 $X2=0
+ $Y2=0
cc_145 N_VPB_M1018_b N_RESET_B_M1024_g 0.111633f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=3.06
cc_146 VPB N_RESET_B_M1024_g 0.00102394f $X=0 $Y=3.955 $X2=0.665 $Y2=3.06
cc_147 N_VPB_c_101_p N_RESET_B_M1024_g 0.0063482f $X=15.12 $Y=4.07 $X2=0.665
+ $Y2=3.06
cc_148 N_VPB_M1018_b N_RESET_B_c_598_n 0.0821685f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_149 N_VPB_M1018_b N_RESET_B_M1006_g 0.0413116f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=1.34
cc_150 VPB N_RESET_B_M1006_g 6.30839e-19 $X=0 $Y=3.955 $X2=0.725 $Y2=1.34
cc_151 N_VPB_c_101_p N_RESET_B_M1006_g 0.00497186f $X=15.12 $Y=4.07 $X2=0.725
+ $Y2=1.34
cc_152 N_VPB_M1018_b N_RESET_B_M1005_g 0.10037f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=1.295
cc_153 N_VPB_M1018_b N_RESET_B_c_603_n 0.0294483f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=2.035
cc_154 N_VPB_M1018_b N_RESET_B_c_582_n 0.005894f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_155 N_VPB_M1018_b N_RESET_B_c_583_n 0.0120245f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_156 N_VPB_M1018_b N_RESET_B_c_590_n 0.0509273f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_157 N_VPB_M1018_b RESET_B 0.00683375f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_158 N_VPB_M1018_b N_D_c_767_n 0.0864139f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=0.745
cc_159 VPB N_D_c_767_n 0.00102394f $X=0 $Y=3.955 $X2=0.685 $Y2=0.745
cc_160 N_VPB_c_101_p N_D_c_767_n 0.0063482f $X=15.12 $Y=4.07 $X2=0.685 $Y2=0.745
cc_161 N_VPB_M1018_b N_D_M1014_g 0.0588822f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_162 N_VPB_M1018_b N_A_339_537#_M1027_g 0.0559056f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_163 N_VPB_M1018_b N_A_339_537#_c_808_n 0.00174272f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=2.035
cc_164 N_VPB_M1018_b N_A_339_537#_c_814_n 0.0247339f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_165 N_VPB_M1018_b N_A_339_537#_c_815_n 2.56298e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_166 N_VPB_M1018_b N_A_339_537#_c_816_n 0.0774673f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_167 N_VPB_c_101_p N_A_339_537#_c_816_n 0.00245646f $X=15.12 $Y=4.07 $X2=0
+ $Y2=0
cc_168 N_VPB_M1018_b N_A_339_537#_c_818_n 0.00294868f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_169 N_VPB_M1018_b N_A_339_537#_c_819_n 0.00836553f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_170 N_VPB_M1018_b N_A_339_537#_c_820_n 0.0241389f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_171 N_VPB_M1018_b N_A_339_537#_c_821_n 0.0206022f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_172 N_VPB_M1018_b N_A_339_537#_c_822_n 0.0201127f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_173 N_VPB_M1018_b N_A_339_537#_c_823_n 0.00111649f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_174 N_VPB_M1018_b N_A_339_537#_c_824_n 0.0155856f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_175 N_VPB_M1018_b N_A_339_537#_c_825_n 0.0034041f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_176 N_VPB_M1018_b N_A_339_537#_c_826_n 0.00337819f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_177 N_VPB_M1018_b N_A_339_537#_M1020_g 0.0221427f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_178 N_VPB_M1018_b N_A_339_537#_c_828_n 0.0559818f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_179 N_VPB_M1018_b N_A_339_537#_c_811_n 0.0130633f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_180 N_VPB_M1018_b N_A_1119_506#_M1026_g 0.0390185f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=1.21
cc_181 VPB N_A_1119_506#_M1026_g 0.00245686f $X=0 $Y=3.955 $X2=0.635 $Y2=1.21
cc_182 N_VPB_c_101_p N_A_1119_506#_M1026_g 0.00781374f $X=15.12 $Y=4.07
+ $X2=0.635 $Y2=1.21
cc_183 N_VPB_M1018_b N_A_1119_506#_c_1010_n 0.0488658f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=1.34
cc_184 N_VPB_M1018_b N_A_1119_506#_c_1004_n 0.0573179f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_185 N_VPB_M1018_b N_A_1119_506#_c_1012_n 0.0481697f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_186 N_VPB_M1018_b N_A_1119_506#_c_1005_n 0.00259335f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_187 N_VPB_M1018_b N_A_921_632#_M1022_g 0.116587f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_188 VPB N_A_921_632#_M1022_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_189 N_VPB_c_101_p N_A_921_632#_M1022_g 0.013715f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_190 N_VPB_M1018_b N_A_921_632#_c_1108_n 0.00278383f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=1.865
cc_191 N_VPB_M1018_b N_A_921_632#_c_1109_n 3.83023e-19 $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=1.295
cc_192 N_VPB_M1018_b N_A_921_632#_c_1100_n 0.0110108f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_193 N_VPB_M1018_b N_A_921_632#_c_1111_n 0.0141742f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_194 N_VPB_M1018_b N_A_921_632#_c_1112_n 0.0209008f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_195 N_VPB_M1018_b N_A_921_632#_c_1113_n 0.011703f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_196 N_VPB_M1018_b N_A_921_632#_c_1114_n 0.00485221f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_197 N_VPB_M1018_b N_A_921_632#_c_1104_n 0.0128668f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_198 N_VPB_M1018_b N_A_2096_417#_M1021_g 0.0373198f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=1.21
cc_199 N_VPB_M1018_b N_A_2096_417#_c_1242_n 0.0607077f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_200 N_VPB_M1018_b N_A_2096_417#_c_1234_n 0.00458905f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=1.865
cc_201 N_VPB_M1018_b N_A_2096_417#_c_1244_n 0.0036003f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=1.665
cc_202 N_VPB_M1018_b N_A_2096_417#_c_1245_n 0.00729768f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=2.035
cc_203 N_VPB_M1018_b N_A_2096_417#_c_1246_n 0.00214269f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_204 N_VPB_M1018_b N_A_2096_417#_c_1247_n 0.0107216f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_205 N_VPB_M1018_b N_A_2096_417#_M1031_g 0.0179113f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_206 N_VPB_M1018_b N_A_1875_543#_c_1324_n 0.0524137f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=1.95
cc_207 N_VPB_M1018_b N_A_1875_543#_M1019_g 0.0428329f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=1.865
cc_208 N_VPB_M1018_b N_A_1875_543#_c_1326_n 0.01382f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_209 N_VPB_M1018_b N_A_1875_543#_c_1327_n 0.0148285f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=1.665
cc_210 N_VPB_M1018_b N_A_1875_543#_c_1334_n 0.00353331f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_211 N_VPB_M1018_b N_A_1875_543#_c_1335_n 0.0141006f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_212 VPB N_A_1875_543#_c_1335_n 7.60114e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_213 N_VPB_c_101_p N_A_1875_543#_c_1335_n 0.0131049f $X=15.12 $Y=4.07 $X2=0
+ $Y2=0
cc_214 N_VPB_M1018_b N_A_1875_543#_c_1338_n 8.18961e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_215 N_VPB_M1018_b N_A_1875_543#_c_1339_n 0.00315273f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_216 N_VPB_M1018_b N_A_1875_543#_c_1329_n 0.00451223f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_217 N_VPB_M1018_b N_A_1875_543#_c_1341_n 0.00817511f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_218 N_VPB_M1018_b N_A_1875_543#_c_1342_n 0.00950759f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_219 N_VPB_M1018_b N_A_1875_543#_c_1343_n 0.0884972f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_220 N_VPB_M1018_b N_A_2649_207#_M1010_g 0.0427937f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_221 VPB N_A_2649_207#_M1010_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_222 N_VPB_c_101_p N_A_2649_207#_M1010_g 0.0159423f $X=15.12 $Y=4.07 $X2=0
+ $Y2=0
cc_223 N_VPB_M1018_b N_A_2649_207#_c_1465_n 0.00627736f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=1.665
cc_224 N_VPB_M1018_b N_A_2649_207#_c_1459_n 0.002891f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_225 N_VPB_M1018_b N_A_2649_207#_c_1460_n 0.023126f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_226 N_VPB_M1018_b N_VPWR_c_1507_n 0.00540376f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=2.035
cc_227 VPB N_VPWR_c_1507_n 0.00166879f $X=0 $Y=3.955 $X2=0.725 $Y2=2.035
cc_228 N_VPB_c_101_p N_VPWR_c_1507_n 0.0254284f $X=15.12 $Y=4.07 $X2=0.725
+ $Y2=2.035
cc_229 N_VPB_M1018_b N_VPWR_c_1510_n 0.00146585f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1510_n 0.00101701f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_231 N_VPB_c_101_p N_VPWR_c_1510_n 0.0138495f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_232 N_VPB_M1018_b N_VPWR_c_1513_n 0.0038263f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1513_n 0.00357564f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_234 N_VPB_c_101_p N_VPWR_c_1513_n 0.0388009f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_235 N_VPB_M1018_b N_VPWR_c_1516_n 0.00402905f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1516_n 0.00363414f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_237 N_VPB_c_101_p N_VPWR_c_1516_n 0.0476105f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_238 N_VPB_M1018_b N_VPWR_c_1519_n 0.0396388f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1519_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_240 N_VPB_c_101_p N_VPWR_c_1519_n 0.0409968f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_241 N_VPB_M1018_b N_VPWR_c_1522_n 0.0486034f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1522_n 0.0025344f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_243 N_VPB_c_101_p N_VPWR_c_1522_n 0.0386183f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_244 N_VPB_M1018_b N_VPWR_c_1525_n 0.0212428f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1525_n 0.00329801f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_246 N_VPB_c_101_p N_VPWR_c_1525_n 0.0447253f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_247 N_VPB_M1018_b N_VPWR_c_1528_n 0.16685f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1528_n 1.63915f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_249 N_VPB_c_101_p N_VPWR_c_1528_n 0.0739966f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_250 N_VPB_M1018_b N_A_452_632#_c_1634_n 0.00995153f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_251 N_VPB_M1018_b N_A_452_632#_c_1635_n 0.00719275f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_252 N_VPB_M1018_b N_A_452_632#_c_1636_n 0.00694031f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=1.34
cc_253 N_VPB_M1018_b N_A_452_632#_c_1637_n 0.00182304f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=1.34
cc_254 N_VPB_M1018_b N_A_452_632#_c_1638_n 0.00300765f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=1.295
cc_255 N_VPB_M1018_b N_A_452_632#_c_1632_n 0.00694928f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_256 N_VPB_M1018_b N_A_452_632#_c_1640_n 0.00373805f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_257 N_VPB_M1018_b N_A_452_632#_c_1641_n 0.00102342f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_258 N_VPB_M1018_b N_Q_c_1696_n 0.0661062f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_259 VPB N_Q_c_1696_n 0.00106913f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_260 N_VPB_c_101_p N_Q_c_1696_n 0.0160028f $X=15.12 $Y=4.07 $X2=0 $Y2=0
cc_261 N_CLK_M1016_g N_A_30_107#_M1028_g 0.0556732f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_262 CLK N_A_30_107#_M1028_g 0.00427849f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_263 N_CLK_M1016_g N_A_30_107#_c_296_n 0.0069987f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_264 CLK N_A_30_107#_c_296_n 0.0727029f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_265 N_CLK_c_264_n N_A_30_107#_c_296_n 0.0427696f $X=0.725 $Y=1.34 $X2=0 $Y2=0
cc_266 N_CLK_M1018_g N_A_30_107#_c_313_n 0.0270173f $X=0.665 $Y=3.06 $X2=0 $Y2=0
cc_267 N_CLK_M1018_g N_A_30_107#_c_316_n 0.0335161f $X=0.665 $Y=3.06 $X2=0 $Y2=0
cc_268 CLK N_A_30_107#_c_316_n 0.0214916f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_269 N_CLK_c_264_n N_A_30_107#_c_316_n 5.93306e-19 $X=0.725 $Y=1.34 $X2=0
+ $Y2=0
cc_270 N_CLK_M1018_g N_A_30_107#_c_356_n 0.00245392f $X=0.665 $Y=3.06 $X2=0
+ $Y2=0
cc_271 CLK N_A_30_107#_c_356_n 0.0123828f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_272 N_CLK_M1018_g N_A_30_107#_c_298_n 0.051902f $X=0.665 $Y=3.06 $X2=0 $Y2=0
cc_273 CLK N_A_30_107#_c_298_n 0.00135612f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_274 N_CLK_c_264_n N_A_30_107#_c_298_n 0.00168194f $X=0.725 $Y=1.34 $X2=0
+ $Y2=0
cc_275 N_CLK_M1018_g N_A_30_107#_c_318_n 0.0011946f $X=0.665 $Y=3.06 $X2=0 $Y2=0
cc_276 N_CLK_M1018_g N_A_30_107#_c_343_n 0.00513266f $X=0.665 $Y=3.06 $X2=0
+ $Y2=0
cc_277 N_CLK_M1018_g N_VPWR_c_1507_n 0.0479648f $X=0.665 $Y=3.06 $X2=0 $Y2=0
cc_278 N_CLK_M1018_g N_VPWR_c_1528_n 0.0127317f $X=0.665 $Y=3.06 $X2=0 $Y2=0
cc_279 N_CLK_M1016_g N_VGND_c_1708_n 0.0414858f $X=0.685 $Y=0.745 $X2=0 $Y2=0
cc_280 CLK N_VGND_c_1708_n 0.0254652f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_281 N_CLK_M1016_g N_VGND_c_1718_n 0.00891597f $X=0.685 $Y=0.745 $X2=0 $Y2=0
cc_282 CLK N_VGND_c_1718_n 0.00119919f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_283 N_CLK_c_264_n N_VGND_c_1718_n 5.19894e-19 $X=0.725 $Y=1.34 $X2=0 $Y2=0
cc_284 N_A_30_107#_c_319_n N_RESET_B_M1024_g 0.0122842f $X=2.67 $Y=3.72 $X2=0
+ $Y2=0
cc_285 N_A_30_107#_c_364_p N_RESET_B_M1024_g 0.0181814f $X=2.755 $Y=3.635 $X2=0
+ $Y2=0
cc_286 N_A_30_107#_c_325_n N_RESET_B_M1024_g 0.0113379f $X=3.53 $Y=3.105 $X2=0
+ $Y2=0
cc_287 N_A_30_107#_c_366_p N_RESET_B_M1024_g 0.00673779f $X=2.84 $Y=3.105 $X2=0
+ $Y2=0
cc_288 N_A_30_107#_c_367_p N_RESET_B_M1024_g 7.37579e-19 $X=3.615 $Y=3.635 $X2=0
+ $Y2=0
cc_289 N_A_30_107#_c_332_n N_RESET_B_M1006_g 0.00317598f $X=6.58 $Y=2.96
+ $X2=15.12 $Y2=0
cc_290 N_A_30_107#_c_369_p N_RESET_B_M1006_g 0.0242843f $X=6.665 $Y=3.635
+ $X2=15.12 $Y2=0
cc_291 N_A_30_107#_c_333_n N_RESET_B_M1006_g 0.0109716f $X=7.44 $Y=3.72
+ $X2=15.12 $Y2=0
cc_292 N_A_30_107#_c_336_n N_RESET_B_M1006_g 0.00438942f $X=6.75 $Y=3.72
+ $X2=15.12 $Y2=0
cc_293 N_A_30_107#_c_339_n N_RESET_B_M1006_g 0.00243209f $X=7.525 $Y=3.635
+ $X2=15.12 $Y2=0
cc_294 N_A_30_107#_c_341_n N_RESET_B_M1006_g 4.32489e-19 $X=7.61 $Y=3.19
+ $X2=15.12 $Y2=0
cc_295 N_A_30_107#_c_332_n N_RESET_B_c_603_n 0.0146364f $X=6.58 $Y=2.96 $X2=0
+ $Y2=0
cc_296 N_A_30_107#_M1008_g N_RESET_B_c_576_n 0.0215138f $X=4.425 $Y=1.075 $X2=0
+ $Y2=0
cc_297 N_A_30_107#_c_294_n N_RESET_B_c_584_n 0.0147224f $X=10.195 $Y=0.935 $X2=0
+ $Y2=0
cc_298 N_A_30_107#_c_294_n N_RESET_B_c_622_n 0.00185701f $X=10.195 $Y=0.935
+ $X2=0 $Y2=0
cc_299 N_A_30_107#_c_364_p N_D_c_767_n 7.37579e-19 $X=2.755 $Y=3.635 $X2=0 $Y2=0
cc_300 N_A_30_107#_c_325_n N_D_c_767_n 0.0180984f $X=3.53 $Y=3.105 $X2=0 $Y2=0
cc_301 N_A_30_107#_c_367_p N_D_c_767_n 0.0180349f $X=3.615 $Y=3.635 $X2=0 $Y2=0
cc_302 N_A_30_107#_c_326_n N_D_c_767_n 0.00800543f $X=5.1 $Y=3.72 $X2=0 $Y2=0
cc_303 N_A_30_107#_c_329_n N_D_c_767_n 0.00459958f $X=3.7 $Y=3.72 $X2=0 $Y2=0
cc_304 N_A_30_107#_M1008_g D 2.6823e-19 $X=4.425 $Y=1.075 $X2=0 $Y2=0
cc_305 N_A_30_107#_M1008_g N_D_M1014_g 0.0597828f $X=4.425 $Y=1.075 $X2=0 $Y2=0
cc_306 N_A_30_107#_c_294_n N_A_339_537#_c_804_n 0.0102134f $X=10.195 $Y=0.935
+ $X2=0 $Y2=0
cc_307 N_A_30_107#_c_386_p N_A_339_537#_c_804_n 5.17359e-19 $X=10.13 $Y=1.25
+ $X2=0 $Y2=0
cc_308 N_A_30_107#_c_303_n N_A_339_537#_c_804_n 0.00350483f $X=10.13 $Y=1.25
+ $X2=0 $Y2=0
cc_309 N_A_30_107#_c_309_n N_A_339_537#_M1027_g 0.011707f $X=9.125 $Y=2.835
+ $X2=0 $Y2=0
cc_310 N_A_30_107#_c_299_n N_A_339_537#_M1027_g 0.00152271f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_311 N_A_30_107#_c_300_n N_A_339_537#_M1027_g 0.00503362f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_312 N_A_30_107#_c_300_n N_A_339_537#_c_805_n 0.0274207f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_313 N_A_30_107#_c_301_n N_A_339_537#_c_805_n 0.0196817f $X=9.965 $Y=1.67
+ $X2=0 $Y2=0
cc_314 N_A_30_107#_c_302_n N_A_339_537#_c_805_n 0.0120928f $X=9.25 $Y=1.67 $X2=0
+ $Y2=0
cc_315 N_A_30_107#_c_386_p N_A_339_537#_c_805_n 0.00145983f $X=10.13 $Y=1.25
+ $X2=0 $Y2=0
cc_316 N_A_30_107#_c_303_n N_A_339_537#_c_805_n 0.0264591f $X=10.13 $Y=1.25
+ $X2=0 $Y2=0
cc_317 N_A_30_107#_M1028_g N_A_339_537#_c_806_n 0.00602693f $X=1.465 $Y=0.745
+ $X2=0 $Y2=0
cc_318 N_A_30_107#_M1028_g N_A_339_537#_c_808_n 0.0432552f $X=1.465 $Y=0.745
+ $X2=0 $Y2=0
cc_319 N_A_30_107#_c_356_n N_A_339_537#_c_808_n 0.00484925f $X=1.405 $Y=2.02
+ $X2=0 $Y2=0
cc_320 N_A_30_107#_M1000_g N_A_339_537#_c_814_n 0.00592745f $X=1.445 $Y=3.06
+ $X2=0 $Y2=0
cc_321 N_A_30_107#_c_356_n N_A_339_537#_c_814_n 0.0151658f $X=1.405 $Y=2.02
+ $X2=0 $Y2=0
cc_322 N_A_30_107#_c_298_n N_A_339_537#_c_814_n 0.0118804f $X=1.405 $Y=2.02
+ $X2=0 $Y2=0
cc_323 N_A_30_107#_c_318_n N_A_339_537#_c_814_n 0.0367959f $X=1.485 $Y=3.635
+ $X2=0 $Y2=0
cc_324 N_A_30_107#_c_319_n N_A_339_537#_c_814_n 0.0169875f $X=2.67 $Y=3.72 $X2=0
+ $Y2=0
cc_325 N_A_30_107#_c_404_p N_A_339_537#_c_814_n 0.0133773f $X=1.405 $Y=2.44
+ $X2=0 $Y2=0
cc_326 N_A_30_107#_M1008_g N_A_339_537#_c_850_n 0.00337673f $X=4.425 $Y=1.075
+ $X2=0 $Y2=0
cc_327 N_A_30_107#_M1028_g N_A_339_537#_c_809_n 0.00506999f $X=1.465 $Y=0.745
+ $X2=0 $Y2=0
cc_328 N_A_30_107#_c_307_n N_A_339_537#_c_815_n 3.77728e-19 $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_329 N_A_30_107#_c_326_n N_A_339_537#_c_815_n 0.00247889f $X=5.1 $Y=3.72 $X2=0
+ $Y2=0
cc_330 N_A_30_107#_c_307_n N_A_339_537#_c_816_n 0.031436f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_331 N_A_30_107#_c_367_p N_A_339_537#_c_816_n 0.00139996f $X=3.615 $Y=3.635
+ $X2=0 $Y2=0
cc_332 N_A_30_107#_c_326_n N_A_339_537#_c_816_n 0.0239927f $X=5.1 $Y=3.72 $X2=0
+ $Y2=0
cc_333 N_A_30_107#_c_412_p N_A_339_537#_c_816_n 0.00105383f $X=5.185 $Y=3.635
+ $X2=0 $Y2=0
cc_334 N_A_30_107#_c_344_n N_A_339_537#_c_816_n 0.0299805f $X=5.145 $Y=2.835
+ $X2=0 $Y2=0
cc_335 N_A_30_107#_c_307_n N_A_339_537#_c_818_n 0.0184349f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_336 N_A_30_107#_c_307_n N_A_339_537#_c_860_n 0.00166743f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_337 N_A_30_107#_M1008_g N_A_339_537#_c_860_n 0.0111039f $X=4.425 $Y=1.075
+ $X2=0 $Y2=0
cc_338 N_A_30_107#_c_307_n N_A_339_537#_c_819_n 0.0176977f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_339 N_A_30_107#_M1008_g N_A_339_537#_c_819_n 0.0103311f $X=4.425 $Y=1.075
+ $X2=0 $Y2=0
cc_340 N_A_30_107#_c_307_n N_A_339_537#_c_820_n 0.00181964f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_341 N_A_30_107#_M1008_g N_A_339_537#_c_820_n 0.00501159f $X=4.425 $Y=1.075
+ $X2=0 $Y2=0
cc_342 N_A_30_107#_c_356_n N_A_339_537#_c_821_n 9.17742e-19 $X=1.405 $Y=2.02
+ $X2=0 $Y2=0
cc_343 N_A_30_107#_c_307_n N_A_339_537#_c_822_n 0.00104214f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_344 N_A_30_107#_c_309_n N_A_339_537#_c_822_n 0.00104513f $X=9.125 $Y=2.835
+ $X2=0 $Y2=0
cc_345 N_A_30_107#_c_299_n N_A_339_537#_c_822_n 0.0194463f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_346 N_A_30_107#_c_300_n N_A_339_537#_c_822_n 0.0159729f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_347 N_A_30_107#_c_301_n N_A_339_537#_c_822_n 0.0159105f $X=9.965 $Y=1.67
+ $X2=0 $Y2=0
cc_348 N_A_30_107#_c_307_n N_A_339_537#_c_823_n 0.00440683f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_349 N_A_30_107#_M1008_g N_A_339_537#_c_823_n 0.0111861f $X=4.425 $Y=1.075
+ $X2=0 $Y2=0
cc_350 N_A_30_107#_c_356_n N_A_339_537#_c_824_n 0.017227f $X=1.405 $Y=2.02 $X2=0
+ $Y2=0
cc_351 N_A_30_107#_c_298_n N_A_339_537#_c_824_n 0.00683577f $X=1.405 $Y=2.02
+ $X2=0 $Y2=0
cc_352 N_A_30_107#_c_299_n N_A_339_537#_c_825_n 8.52356e-19 $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_353 N_A_30_107#_c_301_n N_A_339_537#_c_825_n 0.00843551f $X=9.965 $Y=1.67
+ $X2=0 $Y2=0
cc_354 N_A_30_107#_c_303_n N_A_339_537#_c_825_n 3.26023e-19 $X=10.13 $Y=1.25
+ $X2=0 $Y2=0
cc_355 N_A_30_107#_c_299_n N_A_339_537#_c_826_n 0.0166663f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_356 N_A_30_107#_c_300_n N_A_339_537#_c_826_n 0.00171229f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_357 N_A_30_107#_c_301_n N_A_339_537#_c_826_n 0.0204906f $X=9.965 $Y=1.67
+ $X2=0 $Y2=0
cc_358 N_A_30_107#_c_307_n N_A_339_537#_M1020_g 0.0292792f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_359 N_A_30_107#_M1008_g N_A_339_537#_M1020_g 0.0509791f $X=4.425 $Y=1.075
+ $X2=0 $Y2=0
cc_360 N_A_30_107#_c_301_n N_A_339_537#_c_828_n 0.00293162f $X=9.965 $Y=1.67
+ $X2=0 $Y2=0
cc_361 N_A_30_107#_c_303_n N_A_339_537#_c_828_n 0.0147062f $X=10.13 $Y=1.25
+ $X2=0 $Y2=0
cc_362 N_A_30_107#_c_299_n N_A_339_537#_c_811_n 0.00562685f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_363 N_A_30_107#_c_300_n N_A_339_537#_c_811_n 0.0390777f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_364 N_A_30_107#_c_301_n N_A_339_537#_c_811_n 0.00818113f $X=9.965 $Y=1.67
+ $X2=0 $Y2=0
cc_365 N_A_30_107#_c_340_n N_A_1119_506#_M1022_d 0.00368877f $X=9.08 $Y=3.19
+ $X2=0 $Y2=0
cc_366 N_A_30_107#_c_412_p N_A_1119_506#_M1026_g 0.00144913f $X=5.185 $Y=3.635
+ $X2=0 $Y2=0
cc_367 N_A_30_107#_c_332_n N_A_1119_506#_M1026_g 0.00788541f $X=6.58 $Y=2.96
+ $X2=0 $Y2=0
cc_368 N_A_30_107#_c_369_p N_A_1119_506#_M1026_g 0.00104405f $X=6.665 $Y=3.635
+ $X2=0 $Y2=0
cc_369 N_A_30_107#_c_344_n N_A_1119_506#_M1026_g 0.0402139f $X=5.145 $Y=2.835
+ $X2=0 $Y2=0
cc_370 N_A_30_107#_c_307_n N_A_1119_506#_c_1010_n 0.0402139f $X=4.425 $Y=2.075
+ $X2=15.12 $Y2=0
cc_371 N_A_30_107#_c_450_p N_A_1119_506#_c_1010_n 0.00115694f $X=5.185 $Y=3.045
+ $X2=15.12 $Y2=0
cc_372 N_A_30_107#_c_332_n N_A_1119_506#_c_1010_n 0.021157f $X=6.58 $Y=2.96
+ $X2=15.12 $Y2=0
cc_373 N_A_30_107#_c_307_n N_A_1119_506#_c_1004_n 0.0106778f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_374 N_A_30_107#_c_309_n N_A_1119_506#_c_1023_n 0.00754106f $X=9.125 $Y=2.835
+ $X2=0 $Y2=0
cc_375 N_A_30_107#_c_340_n N_A_1119_506#_c_1023_n 0.0156718f $X=9.08 $Y=3.19
+ $X2=0 $Y2=0
cc_376 N_A_30_107#_c_299_n N_A_1119_506#_c_1023_n 0.0393914f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_377 N_A_30_107#_c_300_n N_A_1119_506#_c_1023_n 0.00677989f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_378 N_A_30_107#_c_299_n N_A_1119_506#_c_1005_n 0.0280683f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_379 N_A_30_107#_c_300_n N_A_1119_506#_c_1005_n 0.00763373f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_380 N_A_30_107#_c_302_n N_A_1119_506#_c_1005_n 0.0138765f $X=9.25 $Y=1.67
+ $X2=0 $Y2=0
cc_381 N_A_30_107#_c_299_n N_A_1119_506#_c_1030_n 0.0123662f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_382 N_A_30_107#_c_300_n N_A_1119_506#_c_1030_n 0.0048839f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_383 N_A_30_107#_c_300_n N_A_1119_506#_c_1006_n 0.00157228f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_384 N_A_30_107#_c_333_n N_A_921_632#_M1022_g 0.00114127f $X=7.44 $Y=3.72
+ $X2=0 $Y2=0
cc_385 N_A_30_107#_c_339_n N_A_921_632#_M1022_g 0.00370885f $X=7.525 $Y=3.635
+ $X2=0 $Y2=0
cc_386 N_A_30_107#_c_340_n N_A_921_632#_M1022_g 0.0420274f $X=9.08 $Y=3.19 $X2=0
+ $Y2=0
cc_387 N_A_30_107#_c_299_n N_A_921_632#_M1022_g 9.79519e-19 $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_388 N_A_30_107#_c_300_n N_A_921_632#_M1022_g 0.0797305f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_389 N_A_30_107#_c_307_n N_A_921_632#_c_1108_n 0.0275976f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_390 N_A_30_107#_c_450_p N_A_921_632#_c_1108_n 0.0225517f $X=5.185 $Y=3.045
+ $X2=0 $Y2=0
cc_391 N_A_30_107#_c_332_n N_A_921_632#_c_1108_n 0.00725053f $X=6.58 $Y=2.96
+ $X2=0 $Y2=0
cc_392 N_A_30_107#_c_307_n N_A_921_632#_c_1109_n 0.0102121f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_393 N_A_30_107#_c_307_n N_A_921_632#_c_1100_n 0.00108736f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_394 N_A_30_107#_c_332_n N_A_921_632#_c_1111_n 0.0734907f $X=6.58 $Y=2.96
+ $X2=0 $Y2=0
cc_395 N_A_30_107#_c_332_n N_A_921_632#_c_1112_n 0.0128825f $X=6.58 $Y=2.96
+ $X2=0 $Y2=0
cc_396 N_A_30_107#_c_369_p N_A_921_632#_c_1112_n 0.0278635f $X=6.665 $Y=3.635
+ $X2=0 $Y2=0
cc_397 N_A_30_107#_c_333_n N_A_921_632#_c_1112_n 0.0209781f $X=7.44 $Y=3.72
+ $X2=0 $Y2=0
cc_398 N_A_30_107#_c_339_n N_A_921_632#_c_1112_n 0.0135834f $X=7.525 $Y=3.635
+ $X2=0 $Y2=0
cc_399 N_A_30_107#_c_341_n N_A_921_632#_c_1112_n 0.0144409f $X=7.61 $Y=3.19
+ $X2=0 $Y2=0
cc_400 N_A_30_107#_c_307_n N_A_921_632#_c_1132_n 0.00117793f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_401 N_A_30_107#_c_326_n N_A_921_632#_c_1132_n 0.0198579f $X=5.1 $Y=3.72 $X2=0
+ $Y2=0
cc_402 N_A_30_107#_c_412_p N_A_921_632#_c_1132_n 0.0165797f $X=5.185 $Y=3.635
+ $X2=0 $Y2=0
cc_403 N_A_30_107#_c_344_n N_A_921_632#_c_1132_n 0.00545322f $X=5.145 $Y=2.835
+ $X2=0 $Y2=0
cc_404 N_A_30_107#_c_307_n N_A_921_632#_c_1113_n 0.00808691f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_405 N_A_30_107#_c_450_p N_A_921_632#_c_1113_n 0.0260081f $X=5.185 $Y=3.045
+ $X2=0 $Y2=0
cc_406 N_A_30_107#_c_412_p N_A_921_632#_c_1113_n 0.00715901f $X=5.185 $Y=3.635
+ $X2=0 $Y2=0
cc_407 N_A_30_107#_c_344_n N_A_921_632#_c_1113_n 0.00447517f $X=5.145 $Y=2.835
+ $X2=0 $Y2=0
cc_408 N_A_30_107#_M1008_g N_A_921_632#_c_1102_n 0.0125685f $X=4.425 $Y=1.075
+ $X2=0 $Y2=0
cc_409 N_A_30_107#_c_307_n N_A_921_632#_c_1114_n 0.00443849f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_410 N_A_30_107#_c_450_p N_A_921_632#_c_1114_n 0.00108474f $X=5.185 $Y=3.045
+ $X2=0 $Y2=0
cc_411 N_A_30_107#_c_332_n N_A_921_632#_c_1114_n 0.0130905f $X=6.58 $Y=2.96
+ $X2=0 $Y2=0
cc_412 N_A_30_107#_c_299_n N_A_921_632#_c_1104_n 4.65016e-19 $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_413 N_A_30_107#_c_300_n N_A_921_632#_c_1104_n 0.00195765f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_414 N_A_30_107#_c_302_n N_A_921_632#_c_1104_n 5.14133e-19 $X=9.25 $Y=1.67
+ $X2=0 $Y2=0
cc_415 N_A_30_107#_c_303_n N_A_2096_417#_c_1249_n 2.52298e-19 $X=10.13 $Y=1.25
+ $X2=15.12 $Y2=0
cc_416 N_A_30_107#_c_294_n N_A_2096_417#_M1031_g 0.0888416f $X=10.195 $Y=0.935
+ $X2=0 $Y2=0
cc_417 N_A_30_107#_c_294_n N_A_1875_543#_c_1328_n 0.00551221f $X=10.195 $Y=0.935
+ $X2=0 $Y2=0
cc_418 N_A_30_107#_c_301_n N_A_1875_543#_c_1328_n 0.0190032f $X=9.965 $Y=1.67
+ $X2=0 $Y2=0
cc_419 N_A_30_107#_c_386_p N_A_1875_543#_c_1328_n 0.0163067f $X=10.13 $Y=1.25
+ $X2=0 $Y2=0
cc_420 N_A_30_107#_c_303_n N_A_1875_543#_c_1328_n 0.00135986f $X=10.13 $Y=1.25
+ $X2=0 $Y2=0
cc_421 N_A_30_107#_c_309_n N_A_1875_543#_c_1334_n 4.57034e-19 $X=9.125 $Y=2.835
+ $X2=0 $Y2=0
cc_422 N_A_30_107#_c_299_n N_A_1875_543#_c_1334_n 0.00724111f $X=9.165 $Y=2.05
+ $X2=0 $Y2=0
cc_423 N_A_30_107#_c_309_n N_A_1875_543#_c_1335_n 0.00382302f $X=9.125 $Y=2.835
+ $X2=0 $Y2=0
cc_424 N_A_30_107#_c_294_n N_A_1875_543#_c_1351_n 0.0299299f $X=10.195 $Y=0.935
+ $X2=0 $Y2=0
cc_425 N_A_30_107#_c_386_p N_A_1875_543#_c_1351_n 0.0118387f $X=10.13 $Y=1.25
+ $X2=0 $Y2=0
cc_426 N_A_30_107#_c_294_n N_A_1875_543#_c_1329_n 0.00486075f $X=10.195 $Y=0.935
+ $X2=0 $Y2=0
cc_427 N_A_30_107#_c_295_n N_A_1875_543#_c_1329_n 0.00704333f $X=10.195 $Y=1.185
+ $X2=0 $Y2=0
cc_428 N_A_30_107#_c_301_n N_A_1875_543#_c_1329_n 0.0123662f $X=9.965 $Y=1.67
+ $X2=0 $Y2=0
cc_429 N_A_30_107#_c_386_p N_A_1875_543#_c_1329_n 0.0336062f $X=10.13 $Y=1.25
+ $X2=0 $Y2=0
cc_430 N_A_30_107#_c_303_n N_A_1875_543#_c_1329_n 0.0127338f $X=10.13 $Y=1.25
+ $X2=0 $Y2=0
cc_431 N_A_30_107#_c_301_n N_A_1875_543#_c_1341_n 0.00410048f $X=9.965 $Y=1.67
+ $X2=0 $Y2=0
cc_432 N_A_30_107#_c_303_n N_A_1875_543#_c_1341_n 0.00580522f $X=10.13 $Y=1.25
+ $X2=0 $Y2=0
cc_433 N_A_30_107#_c_325_n N_VPWR_M1024_d 0.00167928f $X=3.53 $Y=3.105 $X2=0
+ $Y2=0
cc_434 N_A_30_107#_c_340_n N_VPWR_M1022_s 0.0119303f $X=9.08 $Y=3.19 $X2=0 $Y2=0
cc_435 N_A_30_107#_M1000_g N_VPWR_c_1507_n 0.0171307f $X=1.445 $Y=3.06 $X2=0
+ $Y2=0
cc_436 N_A_30_107#_c_313_n N_VPWR_c_1507_n 0.0522997f $X=0.275 $Y=2.83 $X2=0
+ $Y2=0
cc_437 N_A_30_107#_c_316_n N_VPWR_c_1507_n 0.03655f $X=1.24 $Y=2.44 $X2=0 $Y2=0
cc_438 N_A_30_107#_c_318_n N_VPWR_c_1507_n 0.0635801f $X=1.485 $Y=3.635 $X2=0
+ $Y2=0
cc_439 N_A_30_107#_c_322_n N_VPWR_c_1507_n 0.00488837f $X=1.57 $Y=3.72 $X2=0
+ $Y2=0
cc_440 N_A_30_107#_c_319_n N_VPWR_c_1510_n 0.00432581f $X=2.67 $Y=3.72 $X2=0
+ $Y2=0
cc_441 N_A_30_107#_c_364_p N_VPWR_c_1510_n 0.0166877f $X=2.755 $Y=3.635 $X2=0
+ $Y2=0
cc_442 N_A_30_107#_c_325_n N_VPWR_c_1510_n 0.0141955f $X=3.53 $Y=3.105 $X2=0
+ $Y2=0
cc_443 N_A_30_107#_c_367_p N_VPWR_c_1510_n 0.0166877f $X=3.615 $Y=3.635 $X2=0
+ $Y2=0
cc_444 N_A_30_107#_c_329_n N_VPWR_c_1510_n 0.00432581f $X=3.7 $Y=3.72 $X2=0
+ $Y2=0
cc_445 N_A_30_107#_c_326_n N_VPWR_c_1513_n 0.00457995f $X=5.1 $Y=3.72 $X2=0
+ $Y2=0
cc_446 N_A_30_107#_c_412_p N_VPWR_c_1513_n 0.0287713f $X=5.185 $Y=3.635 $X2=0
+ $Y2=0
cc_447 N_A_30_107#_c_332_n N_VPWR_c_1513_n 0.0612799f $X=6.58 $Y=2.96 $X2=0
+ $Y2=0
cc_448 N_A_30_107#_c_369_p N_VPWR_c_1513_n 0.017181f $X=6.665 $Y=3.635 $X2=0
+ $Y2=0
cc_449 N_A_30_107#_c_336_n N_VPWR_c_1513_n 0.00457995f $X=6.75 $Y=3.72 $X2=0
+ $Y2=0
cc_450 N_A_30_107#_c_344_n N_VPWR_c_1513_n 0.00335868f $X=5.145 $Y=2.835 $X2=0
+ $Y2=0
cc_451 N_A_30_107#_c_309_n N_VPWR_c_1516_n 0.00619189f $X=9.125 $Y=2.835 $X2=0
+ $Y2=0
cc_452 N_A_30_107#_c_333_n N_VPWR_c_1516_n 0.00837555f $X=7.44 $Y=3.72 $X2=0
+ $Y2=0
cc_453 N_A_30_107#_c_339_n N_VPWR_c_1516_n 0.0122276f $X=7.525 $Y=3.635 $X2=0
+ $Y2=0
cc_454 N_A_30_107#_c_340_n N_VPWR_c_1516_n 0.0504084f $X=9.08 $Y=3.19 $X2=0
+ $Y2=0
cc_455 N_A_30_107#_M1000_g N_VPWR_c_1528_n 0.019492f $X=1.445 $Y=3.06 $X2=0
+ $Y2=0
cc_456 N_A_30_107#_c_309_n N_VPWR_c_1528_n 0.0220138f $X=9.125 $Y=2.835 $X2=0
+ $Y2=0
cc_457 N_A_30_107#_c_313_n N_VPWR_c_1528_n 0.0261499f $X=0.275 $Y=2.83 $X2=0
+ $Y2=0
cc_458 N_A_30_107#_c_318_n N_VPWR_c_1528_n 0.0205319f $X=1.485 $Y=3.635 $X2=0
+ $Y2=0
cc_459 N_A_30_107#_c_319_n N_VPWR_c_1528_n 0.0510104f $X=2.67 $Y=3.72 $X2=0
+ $Y2=0
cc_460 N_A_30_107#_c_322_n N_VPWR_c_1528_n 0.00776931f $X=1.57 $Y=3.72 $X2=0
+ $Y2=0
cc_461 N_A_30_107#_c_364_p N_VPWR_c_1528_n 0.0138576f $X=2.755 $Y=3.635 $X2=0
+ $Y2=0
cc_462 N_A_30_107#_c_325_n N_VPWR_c_1528_n 0.0158496f $X=3.53 $Y=3.105 $X2=0
+ $Y2=0
cc_463 N_A_30_107#_c_367_p N_VPWR_c_1528_n 0.0138576f $X=3.615 $Y=3.635 $X2=0
+ $Y2=0
cc_464 N_A_30_107#_c_326_n N_VPWR_c_1528_n 0.0583295f $X=5.1 $Y=3.72 $X2=0 $Y2=0
cc_465 N_A_30_107#_c_329_n N_VPWR_c_1528_n 0.00766613f $X=3.7 $Y=3.72 $X2=0
+ $Y2=0
cc_466 N_A_30_107#_c_450_p N_VPWR_c_1528_n 0.00408181f $X=5.185 $Y=3.045 $X2=0
+ $Y2=0
cc_467 N_A_30_107#_c_412_p N_VPWR_c_1528_n 0.0199583f $X=5.185 $Y=3.635 $X2=0
+ $Y2=0
cc_468 N_A_30_107#_c_332_n N_VPWR_c_1528_n 0.015416f $X=6.58 $Y=2.96 $X2=0 $Y2=0
cc_469 N_A_30_107#_c_369_p N_VPWR_c_1528_n 0.0199533f $X=6.665 $Y=3.635 $X2=0
+ $Y2=0
cc_470 N_A_30_107#_c_333_n N_VPWR_c_1528_n 0.0323485f $X=7.44 $Y=3.72 $X2=0
+ $Y2=0
cc_471 N_A_30_107#_c_336_n N_VPWR_c_1528_n 0.00767994f $X=6.75 $Y=3.72 $X2=0
+ $Y2=0
cc_472 N_A_30_107#_c_339_n N_VPWR_c_1528_n 0.0205954f $X=7.525 $Y=3.635 $X2=0
+ $Y2=0
cc_473 N_A_30_107#_c_340_n N_VPWR_c_1528_n 0.0589936f $X=9.08 $Y=3.19 $X2=0
+ $Y2=0
cc_474 N_A_30_107#_c_344_n N_VPWR_c_1528_n 0.00950786f $X=5.145 $Y=2.835 $X2=0
+ $Y2=0
cc_475 N_A_30_107#_c_319_n N_A_452_632#_c_1634_n 0.016639f $X=2.67 $Y=3.72 $X2=0
+ $Y2=0
cc_476 N_A_30_107#_c_364_p N_A_452_632#_c_1634_n 0.00869555f $X=2.755 $Y=3.635
+ $X2=0 $Y2=0
cc_477 N_A_30_107#_c_366_p N_A_452_632#_c_1634_n 0.012185f $X=2.84 $Y=3.105
+ $X2=0 $Y2=0
cc_478 N_A_30_107#_c_325_n N_A_452_632#_c_1635_n 0.0574665f $X=3.53 $Y=3.105
+ $X2=0 $Y2=0
cc_479 N_A_30_107#_c_366_p N_A_452_632#_c_1635_n 0.0120584f $X=2.84 $Y=3.105
+ $X2=0 $Y2=0
cc_480 N_A_30_107#_c_325_n N_A_452_632#_c_1638_n 0.0117279f $X=3.53 $Y=3.105
+ $X2=0 $Y2=0
cc_481 N_A_30_107#_c_367_p N_A_452_632#_c_1638_n 0.00869352f $X=3.615 $Y=3.635
+ $X2=0 $Y2=0
cc_482 N_A_30_107#_c_326_n N_A_452_632#_c_1638_n 0.0112539f $X=5.1 $Y=3.72 $X2=0
+ $Y2=0
cc_483 N_A_30_107#_M1008_g N_A_452_632#_c_1631_n 0.0101889f $X=4.425 $Y=1.075
+ $X2=0 $Y2=0
cc_484 N_A_30_107#_M1008_g N_A_452_632#_c_1632_n 0.00942298f $X=4.425 $Y=1.075
+ $X2=0 $Y2=0
cc_485 N_A_30_107#_c_307_n N_A_452_632#_c_1640_n 0.00942298f $X=4.425 $Y=2.075
+ $X2=0 $Y2=0
cc_486 N_A_30_107#_M1008_g N_A_452_632#_c_1633_n 0.0068356f $X=4.425 $Y=1.075
+ $X2=0 $Y2=0
cc_487 N_A_30_107#_M1028_g N_VGND_c_1708_n 0.0465728f $X=1.465 $Y=0.745 $X2=0
+ $Y2=0
cc_488 N_A_30_107#_c_296_n N_VGND_c_1708_n 0.0231898f $X=0.295 $Y=0.745 $X2=0
+ $Y2=0
cc_489 N_A_30_107#_M1028_g N_VGND_c_1710_n 0.00264212f $X=1.465 $Y=0.745 $X2=0
+ $Y2=0
cc_490 N_A_30_107#_M1016_s N_VGND_c_1718_n 0.00177616f $X=0.15 $Y=0.535 $X2=0
+ $Y2=0
cc_491 N_A_30_107#_M1028_g N_VGND_c_1718_n 0.0118525f $X=1.465 $Y=0.745 $X2=0
+ $Y2=0
cc_492 N_A_30_107#_c_294_n N_VGND_c_1718_n 0.00266367f $X=10.195 $Y=0.935 $X2=0
+ $Y2=0
cc_493 N_A_30_107#_c_296_n N_VGND_c_1718_n 0.0280027f $X=0.295 $Y=0.745 $X2=0
+ $Y2=0
cc_494 N_A_30_107#_c_386_p N_VGND_c_1718_n 0.001544f $X=10.13 $Y=1.25 $X2=0
+ $Y2=0
cc_495 N_RESET_B_M1024_g N_D_c_767_n 0.0434886f $X=2.795 $Y=3.37 $X2=0 $Y2=0
cc_496 N_RESET_B_c_576_n D 0.0224538f $X=5.84 $Y=0.545 $X2=0 $Y2=0
cc_497 N_RESET_B_c_591_n D 0.0793197f $X=2.965 $Y=1.62 $X2=0 $Y2=0
cc_498 N_RESET_B_c_593_n D 0.00149734f $X=2.865 $Y=1.395 $X2=0 $Y2=0
cc_499 N_RESET_B_M1024_g N_D_M1014_g 0.0088148f $X=2.795 $Y=3.37 $X2=0 $Y2=0
cc_500 N_RESET_B_c_576_n N_D_M1014_g 0.0170287f $X=5.84 $Y=0.545 $X2=0 $Y2=0
cc_501 N_RESET_B_c_591_n N_D_M1014_g 0.0163429f $X=2.965 $Y=1.62 $X2=0 $Y2=0
cc_502 N_RESET_B_c_593_n N_D_M1014_g 0.102199f $X=2.865 $Y=1.395 $X2=0 $Y2=0
cc_503 N_RESET_B_c_631_p N_A_339_537#_c_804_n 0.00120637f $X=8.375 $Y=1.125
+ $X2=0 $Y2=0
cc_504 N_RESET_B_c_584_n N_A_339_537#_c_804_n 0.0221897f $X=10.78 $Y=0.35 $X2=0
+ $Y2=0
cc_505 N_RESET_B_c_593_n N_A_339_537#_c_806_n 8.03799e-19 $X=2.865 $Y=1.395
+ $X2=0 $Y2=0
cc_506 N_RESET_B_c_589_n N_A_339_537#_c_808_n 0.0084279f $X=2.86 $Y=1.785 $X2=0
+ $Y2=0
cc_507 N_RESET_B_c_590_n N_A_339_537#_c_808_n 0.0128174f $X=2.86 $Y=1.785 $X2=0
+ $Y2=0
cc_508 N_RESET_B_c_593_n N_A_339_537#_c_808_n 0.00339212f $X=2.865 $Y=1.395
+ $X2=0 $Y2=0
cc_509 N_RESET_B_M1024_g N_A_339_537#_c_814_n 0.0016637f $X=2.795 $Y=3.37 $X2=0
+ $Y2=0
cc_510 N_RESET_B_c_590_n N_A_339_537#_c_814_n 0.0146212f $X=2.86 $Y=1.785 $X2=0
+ $Y2=0
cc_511 N_RESET_B_c_590_n N_A_339_537#_c_820_n 0.0106462f $X=2.86 $Y=1.785 $X2=0
+ $Y2=0
cc_512 RESET_B N_A_339_537#_c_820_n 0.0493112f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_513 N_RESET_B_c_590_n N_A_339_537#_c_821_n 0.00258034f $X=2.86 $Y=1.785 $X2=0
+ $Y2=0
cc_514 RESET_B N_A_339_537#_c_821_n 0.00231338f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_515 N_RESET_B_c_598_n N_A_339_537#_c_822_n 0.007479f $X=6.677 $Y=2.753 $X2=0
+ $Y2=0
cc_516 N_RESET_B_c_582_n N_A_339_537#_c_822_n 0.0543498f $X=8.29 $Y=1.91 $X2=0
+ $Y2=0
cc_517 N_RESET_B_c_583_n N_A_339_537#_c_822_n 0.00268397f $X=6.77 $Y=1.91 $X2=0
+ $Y2=0
cc_518 N_RESET_B_c_590_n N_A_339_537#_c_824_n 0.00453639f $X=2.86 $Y=1.785 $X2=0
+ $Y2=0
cc_519 RESET_B N_A_339_537#_c_824_n 0.00582333f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_520 N_RESET_B_c_576_n N_A_339_537#_M1020_g 0.0158202f $X=5.84 $Y=0.545 $X2=0
+ $Y2=0
cc_521 N_RESET_B_c_580_n N_A_339_537#_M1020_g 0.00178023f $X=5.925 $Y=1.125
+ $X2=0 $Y2=0
cc_522 N_RESET_B_M1006_g N_A_1119_506#_M1026_g 0.0179982f $X=6.705 $Y=3.37 $X2=0
+ $Y2=0
cc_523 N_RESET_B_c_598_n N_A_1119_506#_c_1010_n 0.0392419f $X=6.677 $Y=2.753
+ $X2=15.12 $Y2=0
cc_524 N_RESET_B_M1029_g N_A_1119_506#_c_1002_n 0.0392419f $X=6.65 $Y=1.075
+ $X2=15.12 $Y2=0
cc_525 N_RESET_B_c_581_n N_A_1119_506#_c_1002_n 7.18539e-19 $X=8.29 $Y=1.21
+ $X2=15.12 $Y2=0
cc_526 N_RESET_B_M1029_g N_A_1119_506#_c_1003_n 0.0424628f $X=6.65 $Y=1.075
+ $X2=0 $Y2=0
cc_527 N_RESET_B_c_576_n N_A_1119_506#_c_1003_n 0.0077764f $X=5.84 $Y=0.545
+ $X2=0 $Y2=0
cc_528 N_RESET_B_c_580_n N_A_1119_506#_c_1003_n 0.0207401f $X=5.925 $Y=1.125
+ $X2=0 $Y2=0
cc_529 N_RESET_B_c_581_n N_A_1119_506#_c_1003_n 0.00946316f $X=8.29 $Y=1.21
+ $X2=0 $Y2=0
cc_530 N_RESET_B_c_658_p N_A_1119_506#_c_1003_n 0.00678279f $X=6.01 $Y=1.21
+ $X2=0 $Y2=0
cc_531 N_RESET_B_c_582_n N_A_1119_506#_c_1042_n 0.00575289f $X=8.29 $Y=1.91
+ $X2=7.68 $Y2=0
cc_532 N_RESET_B_c_583_n N_A_1119_506#_c_1042_n 0.00240669f $X=6.77 $Y=1.91
+ $X2=7.68 $Y2=0
cc_533 N_RESET_B_c_582_n N_A_1119_506#_c_1004_n 4.72845e-19 $X=8.29 $Y=1.91
+ $X2=0 $Y2=0
cc_534 N_RESET_B_c_583_n N_A_1119_506#_c_1004_n 0.0392419f $X=6.77 $Y=1.91 $X2=0
+ $Y2=0
cc_535 N_RESET_B_c_598_n N_A_1119_506#_c_1012_n 0.0316179f $X=6.677 $Y=2.753
+ $X2=0 $Y2=0
cc_536 N_RESET_B_c_582_n N_A_1119_506#_c_1012_n 0.108896f $X=8.29 $Y=1.91 $X2=0
+ $Y2=0
cc_537 N_RESET_B_c_631_p N_A_1119_506#_c_1048_n 0.0346849f $X=8.375 $Y=1.125
+ $X2=0 $Y2=0
cc_538 N_RESET_B_c_584_n N_A_1119_506#_c_1048_n 0.0199335f $X=10.78 $Y=0.35
+ $X2=0 $Y2=0
cc_539 N_RESET_B_c_667_p N_A_1119_506#_c_1048_n 0.0129227f $X=8.375 $Y=1.21
+ $X2=0 $Y2=0
cc_540 N_RESET_B_c_582_n N_A_1119_506#_c_1005_n 0.012678f $X=8.29 $Y=1.91 $X2=0
+ $Y2=0
cc_541 N_RESET_B_c_669_p N_A_1119_506#_c_1006_n 0.0353439f $X=8.375 $Y=1.825
+ $X2=0 $Y2=0
cc_542 N_RESET_B_c_582_n N_A_921_632#_M1022_g 0.00945079f $X=8.29 $Y=1.91 $X2=0
+ $Y2=0
cc_543 N_RESET_B_c_581_n N_A_921_632#_c_1097_n 0.0119619f $X=8.29 $Y=1.21 $X2=0
+ $Y2=0
cc_544 N_RESET_B_c_631_p N_A_921_632#_c_1097_n 0.0318677f $X=8.375 $Y=1.125
+ $X2=0 $Y2=0
cc_545 N_RESET_B_c_669_p N_A_921_632#_c_1097_n 0.00659601f $X=8.375 $Y=1.825
+ $X2=0 $Y2=0
cc_546 N_RESET_B_c_584_n N_A_921_632#_c_1097_n 0.00891555f $X=10.78 $Y=0.35
+ $X2=0 $Y2=0
cc_547 N_RESET_B_c_586_n N_A_921_632#_c_1097_n 0.00353941f $X=8.46 $Y=0.35 $X2=0
+ $Y2=0
cc_548 N_RESET_B_c_667_p N_A_921_632#_c_1097_n 0.00513124f $X=8.375 $Y=1.21
+ $X2=0 $Y2=0
cc_549 N_RESET_B_c_576_n N_A_921_632#_c_1154_n 0.0189379f $X=5.84 $Y=0.545
+ $X2=7.68 $Y2=0
cc_550 N_RESET_B_c_658_p N_A_921_632#_c_1099_n 0.00233777f $X=6.01 $Y=1.21 $X2=0
+ $Y2=0
cc_551 N_RESET_B_M1029_g N_A_921_632#_c_1101_n 0.0296912f $X=6.65 $Y=1.075 $X2=0
+ $Y2=0
cc_552 N_RESET_B_c_581_n N_A_921_632#_c_1101_n 0.145457f $X=8.29 $Y=1.21 $X2=0
+ $Y2=0
cc_553 N_RESET_B_c_658_p N_A_921_632#_c_1101_n 0.0122858f $X=6.01 $Y=1.21 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_582_n N_A_921_632#_c_1101_n 0.0962274f $X=8.29 $Y=1.91 $X2=0
+ $Y2=0
cc_555 N_RESET_B_c_583_n N_A_921_632#_c_1101_n 0.00161874f $X=6.77 $Y=1.91 $X2=0
+ $Y2=0
cc_556 N_RESET_B_c_669_p N_A_921_632#_c_1101_n 0.0122207f $X=8.375 $Y=1.825
+ $X2=0 $Y2=0
cc_557 N_RESET_B_c_598_n N_A_921_632#_c_1111_n 0.0343338f $X=6.677 $Y=2.753
+ $X2=0 $Y2=0
cc_558 N_RESET_B_c_598_n N_A_921_632#_c_1112_n 0.0037888f $X=6.677 $Y=2.753
+ $X2=0 $Y2=0
cc_559 N_RESET_B_M1006_g N_A_921_632#_c_1112_n 0.00976932f $X=6.705 $Y=3.37
+ $X2=0 $Y2=0
cc_560 N_RESET_B_c_603_n N_A_921_632#_c_1112_n 0.0139618f $X=6.677 $Y=3.03 $X2=0
+ $Y2=0
cc_561 N_RESET_B_c_576_n N_A_921_632#_c_1102_n 0.0211665f $X=5.84 $Y=0.545 $X2=0
+ $Y2=0
cc_562 N_RESET_B_c_581_n N_A_921_632#_c_1104_n 0.0111689f $X=8.29 $Y=1.21 $X2=0
+ $Y2=0
cc_563 N_RESET_B_c_582_n N_A_921_632#_c_1104_n 0.0219928f $X=8.29 $Y=1.91 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_669_p N_A_921_632#_c_1104_n 0.0259698f $X=8.375 $Y=1.825
+ $X2=0 $Y2=0
cc_565 N_RESET_B_M1005_g N_A_2096_417#_M1021_g 0.0157965f $X=11.615 $Y=2.925
+ $X2=0 $Y2=0
cc_566 N_RESET_B_M1005_g N_A_2096_417#_c_1242_n 0.0544346f $X=11.615 $Y=2.925
+ $X2=0 $Y2=0
cc_567 N_RESET_B_c_588_n N_A_2096_417#_c_1249_n 0.0131366f $X=11.455 $Y=1.18
+ $X2=15.12 $Y2=0
cc_568 N_RESET_B_c_696_p N_A_2096_417#_c_1249_n 0.0114678f $X=10.95 $Y=1.18
+ $X2=15.12 $Y2=0
cc_569 N_RESET_B_c_697_p N_A_2096_417#_c_1249_n 0.00949758f $X=11.62 $Y=1.23
+ $X2=15.12 $Y2=0
cc_570 N_RESET_B_c_592_n N_A_2096_417#_c_1249_n 0.00210584f $X=11.62 $Y=1.23
+ $X2=15.12 $Y2=0
cc_571 N_RESET_B_M1005_g N_A_2096_417#_c_1234_n 0.0290733f $X=11.615 $Y=2.925
+ $X2=0 $Y2=0
cc_572 N_RESET_B_c_588_n N_A_2096_417#_c_1234_n 0.00955743f $X=11.455 $Y=1.18
+ $X2=0 $Y2=0
cc_573 N_RESET_B_c_697_p N_A_2096_417#_c_1234_n 0.0234754f $X=11.62 $Y=1.23
+ $X2=0 $Y2=0
cc_574 N_RESET_B_c_592_n N_A_2096_417#_c_1234_n 0.00320447f $X=11.62 $Y=1.23
+ $X2=0 $Y2=0
cc_575 N_RESET_B_M1005_g N_A_2096_417#_c_1244_n 0.0126705f $X=11.615 $Y=2.925
+ $X2=7.68 $Y2=0.057
cc_576 N_RESET_B_M1005_g N_A_2096_417#_c_1246_n 0.00905379f $X=11.615 $Y=2.925
+ $X2=0 $Y2=0
cc_577 N_RESET_B_c_594_n N_A_2096_417#_c_1235_n 3.15636e-19 $X=11.65 $Y=1.065
+ $X2=0 $Y2=0
cc_578 N_RESET_B_c_592_n N_A_2096_417#_c_1237_n 0.00130113f $X=11.62 $Y=1.23
+ $X2=0 $Y2=0
cc_579 N_RESET_B_c_594_n N_A_2096_417#_c_1238_n 0.00130113f $X=11.65 $Y=1.065
+ $X2=0 $Y2=0
cc_580 N_RESET_B_c_584_n N_A_2096_417#_M1031_g 0.00934051f $X=10.78 $Y=0.35
+ $X2=0 $Y2=0
cc_581 N_RESET_B_c_622_n N_A_2096_417#_M1031_g 0.0259581f $X=10.865 $Y=1.095
+ $X2=0 $Y2=0
cc_582 N_RESET_B_c_588_n N_A_2096_417#_M1031_g 0.0120023f $X=11.455 $Y=1.18
+ $X2=0 $Y2=0
cc_583 N_RESET_B_c_696_p N_A_2096_417#_M1031_g 0.00757277f $X=10.95 $Y=1.18
+ $X2=0 $Y2=0
cc_584 N_RESET_B_c_697_p N_A_2096_417#_M1031_g 0.00177972f $X=11.62 $Y=1.23
+ $X2=0 $Y2=0
cc_585 N_RESET_B_c_592_n N_A_2096_417#_M1031_g 0.0544346f $X=11.62 $Y=1.23 $X2=0
+ $Y2=0
cc_586 N_RESET_B_c_594_n N_A_2096_417#_M1031_g 0.0135357f $X=11.65 $Y=1.065
+ $X2=0 $Y2=0
cc_587 N_RESET_B_c_697_p N_A_1875_543#_M1023_g 0.00298948f $X=11.62 $Y=1.23
+ $X2=0 $Y2=0
cc_588 N_RESET_B_c_594_n N_A_1875_543#_M1023_g 0.0480303f $X=11.65 $Y=1.065
+ $X2=0 $Y2=0
cc_589 N_RESET_B_M1005_g N_A_1875_543#_c_1326_n 0.058805f $X=11.615 $Y=2.925
+ $X2=0 $Y2=0
cc_590 N_RESET_B_c_592_n N_A_1875_543#_c_1326_n 0.0480303f $X=11.62 $Y=1.23
+ $X2=0 $Y2=0
cc_591 N_RESET_B_c_584_n N_A_1875_543#_c_1364_n 0.0211392f $X=10.78 $Y=0.35
+ $X2=0 $Y2=0
cc_592 N_RESET_B_c_584_n N_A_1875_543#_c_1351_n 0.0511362f $X=10.78 $Y=0.35
+ $X2=0 $Y2=0
cc_593 N_RESET_B_c_622_n N_A_1875_543#_c_1351_n 0.00568401f $X=10.865 $Y=1.095
+ $X2=0 $Y2=0
cc_594 N_RESET_B_c_622_n N_A_1875_543#_c_1329_n 0.0150257f $X=10.865 $Y=1.095
+ $X2=0 $Y2=0
cc_595 N_RESET_B_c_696_p N_A_1875_543#_c_1329_n 0.0130055f $X=10.95 $Y=1.18
+ $X2=0 $Y2=0
cc_596 N_RESET_B_M1005_g N_A_1875_543#_c_1342_n 0.0381274f $X=11.615 $Y=2.925
+ $X2=0 $Y2=0
cc_597 N_RESET_B_M1024_g N_VPWR_c_1510_n 0.00576304f $X=2.795 $Y=3.37 $X2=0
+ $Y2=0
cc_598 N_RESET_B_M1006_g N_VPWR_c_1513_n 0.00343208f $X=6.705 $Y=3.37 $X2=0
+ $Y2=0
cc_599 N_RESET_B_M1005_g N_VPWR_c_1519_n 0.0317984f $X=11.615 $Y=2.925 $X2=0
+ $Y2=0
cc_600 N_RESET_B_M1005_g N_VPWR_c_1522_n 6.04648e-19 $X=11.615 $Y=2.925 $X2=0
+ $Y2=0
cc_601 N_RESET_B_M1024_g N_VPWR_c_1528_n 0.00861444f $X=2.795 $Y=3.37 $X2=0
+ $Y2=0
cc_602 N_RESET_B_M1006_g N_VPWR_c_1528_n 0.0150028f $X=6.705 $Y=3.37 $X2=0 $Y2=0
cc_603 N_RESET_B_M1005_g N_VPWR_c_1528_n 0.0135073f $X=11.615 $Y=2.925 $X2=0
+ $Y2=0
cc_604 N_RESET_B_M1024_g N_A_452_632#_c_1634_n 0.012368f $X=2.795 $Y=3.37 $X2=0
+ $Y2=0
cc_605 N_RESET_B_M1024_g N_A_452_632#_c_1635_n 0.0299996f $X=2.795 $Y=3.37 $X2=0
+ $Y2=0
cc_606 N_RESET_B_c_590_n N_A_452_632#_c_1635_n 6.32641e-19 $X=2.86 $Y=1.785
+ $X2=0 $Y2=0
cc_607 RESET_B N_A_452_632#_c_1635_n 0.0395447f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_608 N_RESET_B_c_576_n N_A_452_632#_c_1631_n 0.0178153f $X=5.84 $Y=0.545 $X2=0
+ $Y2=0
cc_609 RESET_B N_A_452_632#_c_1640_n 0.0049369f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_610 N_RESET_B_c_581_n N_VGND_M1029_d 0.0218147f $X=8.29 $Y=1.21 $X2=0 $Y2=0
cc_611 N_RESET_B_c_578_n N_VGND_c_1710_n 0.00792736f $X=3.235 $Y=0.545 $X2=0
+ $Y2=0
cc_612 N_RESET_B_c_589_n N_VGND_c_1710_n 0.00414707f $X=2.86 $Y=1.785 $X2=0
+ $Y2=0
cc_613 N_RESET_B_c_590_n N_VGND_c_1710_n 0.00551305f $X=2.86 $Y=1.785 $X2=0
+ $Y2=0
cc_614 N_RESET_B_c_591_n N_VGND_c_1710_n 0.0322297f $X=2.965 $Y=1.62 $X2=0 $Y2=0
cc_615 N_RESET_B_c_593_n N_VGND_c_1710_n 0.0221614f $X=2.865 $Y=1.395 $X2=0
+ $Y2=0
cc_616 N_RESET_B_M1029_g N_VGND_c_1712_n 0.00881572f $X=6.65 $Y=1.075 $X2=0
+ $Y2=0
cc_617 N_RESET_B_c_581_n N_VGND_c_1712_n 0.0699268f $X=8.29 $Y=1.21 $X2=0 $Y2=0
cc_618 N_RESET_B_c_631_p N_VGND_c_1712_n 0.0212201f $X=8.375 $Y=1.125 $X2=0
+ $Y2=0
cc_619 N_RESET_B_c_586_n N_VGND_c_1712_n 0.00473621f $X=8.46 $Y=0.35 $X2=0 $Y2=0
cc_620 N_RESET_B_c_584_n N_VGND_c_1714_n 0.00461601f $X=10.78 $Y=0.35 $X2=0
+ $Y2=0
cc_621 N_RESET_B_c_622_n N_VGND_c_1714_n 0.0327013f $X=10.865 $Y=1.095 $X2=0
+ $Y2=0
cc_622 N_RESET_B_c_588_n N_VGND_c_1714_n 0.0188137f $X=11.455 $Y=1.18 $X2=0
+ $Y2=0
cc_623 N_RESET_B_c_697_p N_VGND_c_1714_n 0.0245795f $X=11.62 $Y=1.23 $X2=0 $Y2=0
cc_624 N_RESET_B_c_592_n N_VGND_c_1714_n 0.00176966f $X=11.62 $Y=1.23 $X2=0
+ $Y2=0
cc_625 N_RESET_B_c_594_n N_VGND_c_1714_n 0.0486062f $X=11.65 $Y=1.065 $X2=0
+ $Y2=0
cc_626 N_RESET_B_M1029_g N_VGND_c_1718_n 0.016332f $X=6.65 $Y=1.075 $X2=0 $Y2=0
cc_627 N_RESET_B_c_576_n N_VGND_c_1718_n 0.147599f $X=5.84 $Y=0.545 $X2=0 $Y2=0
cc_628 N_RESET_B_c_578_n N_VGND_c_1718_n 0.0141563f $X=3.235 $Y=0.545 $X2=0
+ $Y2=0
cc_629 N_RESET_B_c_581_n N_VGND_c_1718_n 0.0489825f $X=8.29 $Y=1.21 $X2=0 $Y2=0
cc_630 N_RESET_B_c_631_p N_VGND_c_1718_n 0.0199533f $X=8.375 $Y=1.125 $X2=0
+ $Y2=0
cc_631 N_RESET_B_c_584_n N_VGND_c_1718_n 0.0857538f $X=10.78 $Y=0.35 $X2=0 $Y2=0
cc_632 N_RESET_B_c_586_n N_VGND_c_1718_n 0.00776561f $X=8.46 $Y=0.35 $X2=0 $Y2=0
cc_633 N_RESET_B_c_622_n N_VGND_c_1718_n 0.0199528f $X=10.865 $Y=1.095 $X2=0
+ $Y2=0
cc_634 N_RESET_B_c_588_n N_VGND_c_1718_n 0.00669854f $X=11.455 $Y=1.18 $X2=0
+ $Y2=0
cc_635 N_RESET_B_c_697_p N_VGND_c_1718_n 0.00135575f $X=11.62 $Y=1.23 $X2=0
+ $Y2=0
cc_636 N_RESET_B_c_593_n N_VGND_c_1718_n 0.00903327f $X=2.865 $Y=1.395 $X2=0
+ $Y2=0
cc_637 N_RESET_B_c_581_n A_1233_173# 0.00223175f $X=8.29 $Y=1.21 $X2=0 $Y2=0
cc_638 N_D_c_767_n N_A_339_537#_c_815_n 2.5842e-19 $X=3.61 $Y=3.05 $X2=0 $Y2=0
cc_639 N_D_c_767_n N_A_339_537#_c_816_n 0.040362f $X=3.61 $Y=3.05 $X2=0 $Y2=0
cc_640 N_D_M1014_g N_A_339_537#_c_818_n 0.00111565f $X=3.645 $Y=1.075 $X2=0
+ $Y2=0
cc_641 N_D_c_767_n N_A_339_537#_c_820_n 0.00165925f $X=3.61 $Y=3.05 $X2=0 $Y2=0
cc_642 D N_A_339_537#_c_820_n 0.0279247f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_643 N_D_M1014_g N_A_339_537#_c_820_n 0.0157014f $X=3.645 $Y=1.075 $X2=0 $Y2=0
cc_644 N_D_c_767_n N_VPWR_c_1510_n 0.00576304f $X=3.61 $Y=3.05 $X2=0 $Y2=0
cc_645 N_D_c_767_n N_VPWR_c_1528_n 0.00853934f $X=3.61 $Y=3.05 $X2=0 $Y2=0
cc_646 N_D_c_767_n N_A_452_632#_c_1635_n 0.0337593f $X=3.61 $Y=3.05 $X2=0 $Y2=0
cc_647 D N_A_452_632#_c_1635_n 0.00444654f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_648 N_D_c_767_n N_A_452_632#_c_1637_n 0.00725092f $X=3.61 $Y=3.05 $X2=15.12
+ $Y2=0
cc_649 N_D_M1014_g N_A_452_632#_c_1637_n 0.00350467f $X=3.645 $Y=1.075 $X2=15.12
+ $Y2=0
cc_650 N_D_c_767_n N_A_452_632#_c_1638_n 0.0106687f $X=3.61 $Y=3.05 $X2=0 $Y2=0
cc_651 D N_A_452_632#_c_1631_n 0.0742844f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_652 N_D_M1014_g N_A_452_632#_c_1631_n 0.0131439f $X=3.645 $Y=1.075 $X2=0
+ $Y2=0
cc_653 N_D_M1014_g N_A_452_632#_c_1640_n 0.00656151f $X=3.645 $Y=1.075 $X2=0
+ $Y2=0
cc_654 N_D_c_767_n N_A_452_632#_c_1641_n 0.00122231f $X=3.61 $Y=3.05 $X2=0 $Y2=0
cc_655 D N_VGND_c_1718_n 0.00254029f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_656 N_A_339_537#_c_850_n N_A_1119_506#_c_1002_n 2.40057e-19 $X=5.14 $Y=1.57
+ $X2=15.12 $Y2=0
cc_657 N_A_339_537#_M1020_g N_A_1119_506#_c_1003_n 0.0884754f $X=5.205 $Y=1.075
+ $X2=0 $Y2=0
cc_658 N_A_339_537#_c_822_n N_A_1119_506#_c_1042_n 0.0195049f $X=9.695 $Y=2.035
+ $X2=7.68 $Y2=0
cc_659 N_A_339_537#_c_822_n N_A_1119_506#_c_1004_n 0.00614569f $X=9.695 $Y=2.035
+ $X2=0 $Y2=0
cc_660 N_A_339_537#_c_822_n N_A_1119_506#_c_1012_n 0.0681002f $X=9.695 $Y=2.035
+ $X2=0 $Y2=0
cc_661 N_A_339_537#_c_804_n N_A_1119_506#_c_1048_n 0.0153829f $X=9.195 $Y=1.395
+ $X2=0 $Y2=0
cc_662 N_A_339_537#_c_804_n N_A_1119_506#_c_1005_n 0.0078944f $X=9.195 $Y=1.395
+ $X2=0 $Y2=0
cc_663 N_A_339_537#_c_822_n N_A_1119_506#_c_1005_n 0.0364434f $X=9.695 $Y=2.035
+ $X2=0 $Y2=0
cc_664 N_A_339_537#_c_811_n N_A_1119_506#_c_1005_n 4.20779e-19 $X=9.905 $Y=2.085
+ $X2=0 $Y2=0
cc_665 N_A_339_537#_c_822_n N_A_1119_506#_c_1030_n 0.00389023f $X=9.695 $Y=2.035
+ $X2=0 $Y2=0
cc_666 N_A_339_537#_c_804_n N_A_1119_506#_c_1006_n 0.00534901f $X=9.195 $Y=1.395
+ $X2=0 $Y2=0
cc_667 N_A_339_537#_c_822_n N_A_921_632#_M1022_g 0.0126067f $X=9.695 $Y=2.035
+ $X2=0 $Y2=0
cc_668 N_A_339_537#_c_804_n N_A_921_632#_c_1097_n 0.0131667f $X=9.195 $Y=1.395
+ $X2=0 $Y2=0
cc_669 N_A_339_537#_c_819_n N_A_921_632#_c_1108_n 0.034714f $X=4.975 $Y=2.035
+ $X2=0 $Y2=0
cc_670 N_A_339_537#_c_822_n N_A_921_632#_c_1108_n 0.0108728f $X=9.695 $Y=2.035
+ $X2=0 $Y2=0
cc_671 N_A_339_537#_M1020_g N_A_921_632#_c_1108_n 0.00291112f $X=5.205 $Y=1.075
+ $X2=0 $Y2=0
cc_672 N_A_339_537#_c_818_n N_A_921_632#_c_1109_n 0.0127006f $X=4.34 $Y=2.67
+ $X2=0 $Y2=0
cc_673 N_A_339_537#_c_819_n N_A_921_632#_c_1109_n 0.0112822f $X=4.975 $Y=2.035
+ $X2=0 $Y2=0
cc_674 N_A_339_537#_c_822_n N_A_921_632#_c_1109_n 6.81135e-19 $X=9.695 $Y=2.035
+ $X2=0 $Y2=0
cc_675 N_A_339_537#_c_823_n N_A_921_632#_c_1109_n 0.00179568f $X=4.705 $Y=2.035
+ $X2=0 $Y2=0
cc_676 N_A_339_537#_c_850_n N_A_921_632#_c_1154_n 0.0235686f $X=5.14 $Y=1.57
+ $X2=7.68 $Y2=0
cc_677 N_A_339_537#_M1020_g N_A_921_632#_c_1154_n 0.0294605f $X=5.205 $Y=1.075
+ $X2=7.68 $Y2=0
cc_678 N_A_339_537#_c_850_n N_A_921_632#_c_1099_n 0.00348991f $X=5.14 $Y=1.57
+ $X2=0 $Y2=0
cc_679 N_A_339_537#_M1020_g N_A_921_632#_c_1099_n 0.00397359f $X=5.205 $Y=1.075
+ $X2=0 $Y2=0
cc_680 N_A_339_537#_c_850_n N_A_921_632#_c_1100_n 0.0193189f $X=5.14 $Y=1.57
+ $X2=0 $Y2=0
cc_681 N_A_339_537#_c_819_n N_A_921_632#_c_1100_n 0.0158435f $X=4.975 $Y=2.035
+ $X2=0 $Y2=0
cc_682 N_A_339_537#_c_822_n N_A_921_632#_c_1100_n 0.0219382f $X=9.695 $Y=2.035
+ $X2=0 $Y2=0
cc_683 N_A_339_537#_M1020_g N_A_921_632#_c_1100_n 0.00309961f $X=5.205 $Y=1.075
+ $X2=0 $Y2=0
cc_684 N_A_339_537#_c_822_n N_A_921_632#_c_1101_n 0.0255245f $X=9.695 $Y=2.035
+ $X2=0 $Y2=0
cc_685 N_A_339_537#_c_822_n N_A_921_632#_c_1111_n 0.00787454f $X=9.695 $Y=2.035
+ $X2=0 $Y2=0
cc_686 N_A_339_537#_c_816_n N_A_921_632#_c_1132_n 0.00756007f $X=4.34 $Y=2.835
+ $X2=0 $Y2=0
cc_687 N_A_339_537#_c_816_n N_A_921_632#_c_1113_n 0.00525464f $X=4.34 $Y=2.835
+ $X2=0 $Y2=0
cc_688 N_A_339_537#_c_818_n N_A_921_632#_c_1113_n 0.0352617f $X=4.34 $Y=2.67
+ $X2=0 $Y2=0
cc_689 N_A_339_537#_c_819_n N_A_921_632#_c_1102_n 0.00725412f $X=4.975 $Y=2.035
+ $X2=0 $Y2=0
cc_690 N_A_339_537#_M1020_g N_A_921_632#_c_1102_n 0.00839629f $X=5.205 $Y=1.075
+ $X2=0 $Y2=0
cc_691 N_A_339_537#_c_850_n N_A_921_632#_c_1103_n 0.0134501f $X=5.14 $Y=1.57
+ $X2=0 $Y2=0
cc_692 N_A_339_537#_M1020_g N_A_921_632#_c_1103_n 0.00150062f $X=5.205 $Y=1.075
+ $X2=0 $Y2=0
cc_693 N_A_339_537#_c_805_n N_A_921_632#_c_1104_n 0.0131667f $X=9.647 $Y=1.525
+ $X2=0 $Y2=0
cc_694 N_A_339_537#_c_822_n N_A_921_632#_c_1104_n 0.00135956f $X=9.695 $Y=2.035
+ $X2=0 $Y2=0
cc_695 N_A_339_537#_M1027_g N_A_2096_417#_M1021_g 0.0400147f $X=10.02 $Y=2.925
+ $X2=0 $Y2=0
cc_696 N_A_339_537#_c_826_n N_A_2096_417#_c_1242_n 2.23203e-19 $X=9.84 $Y=2.035
+ $X2=0 $Y2=0
cc_697 N_A_339_537#_c_828_n N_A_2096_417#_c_1242_n 0.0400147f $X=9.79 $Y=2.27
+ $X2=0 $Y2=0
cc_698 N_A_339_537#_c_804_n N_A_1875_543#_c_1364_n 0.00452157f $X=9.195 $Y=1.395
+ $X2=0 $Y2=0
cc_699 N_A_339_537#_c_804_n N_A_1875_543#_c_1328_n 0.0156863f $X=9.195 $Y=1.395
+ $X2=0 $Y2=0
cc_700 N_A_339_537#_c_805_n N_A_1875_543#_c_1328_n 0.0095296f $X=9.647 $Y=1.525
+ $X2=0 $Y2=0
cc_701 N_A_339_537#_c_822_n N_A_1875_543#_c_1334_n 0.00703926f $X=9.695 $Y=2.035
+ $X2=0 $Y2=0
cc_702 N_A_339_537#_c_826_n N_A_1875_543#_c_1334_n 0.00338612f $X=9.84 $Y=2.035
+ $X2=0 $Y2=0
cc_703 N_A_339_537#_c_828_n N_A_1875_543#_c_1334_n 0.00426537f $X=9.79 $Y=2.27
+ $X2=0 $Y2=0
cc_704 N_A_339_537#_M1027_g N_A_1875_543#_c_1335_n 0.0115771f $X=10.02 $Y=2.925
+ $X2=0 $Y2=0
cc_705 N_A_339_537#_M1027_g N_A_1875_543#_c_1338_n 0.0321274f $X=10.02 $Y=2.925
+ $X2=0 $Y2=0
cc_706 N_A_339_537#_c_825_n N_A_1875_543#_c_1338_n 0.00185975f $X=9.84 $Y=2.035
+ $X2=0 $Y2=0
cc_707 N_A_339_537#_c_826_n N_A_1875_543#_c_1338_n 0.0147007f $X=9.84 $Y=2.035
+ $X2=0 $Y2=0
cc_708 N_A_339_537#_c_828_n N_A_1875_543#_c_1338_n 5.81569e-19 $X=9.79 $Y=2.27
+ $X2=0 $Y2=0
cc_709 N_A_339_537#_M1027_g N_A_1875_543#_c_1339_n 0.0132244f $X=10.02 $Y=2.925
+ $X2=0 $Y2=0
cc_710 N_A_339_537#_c_826_n N_A_1875_543#_c_1339_n 0.00545705f $X=9.84 $Y=2.035
+ $X2=0 $Y2=0
cc_711 N_A_339_537#_c_828_n N_A_1875_543#_c_1339_n 0.00311909f $X=9.79 $Y=2.27
+ $X2=0 $Y2=0
cc_712 N_A_339_537#_c_825_n N_A_1875_543#_c_1329_n 0.00602337f $X=9.84 $Y=2.035
+ $X2=0 $Y2=0
cc_713 N_A_339_537#_c_826_n N_A_1875_543#_c_1329_n 0.00592974f $X=9.84 $Y=2.035
+ $X2=0 $Y2=0
cc_714 N_A_339_537#_c_828_n N_A_1875_543#_c_1329_n 9.28046e-19 $X=9.79 $Y=2.27
+ $X2=0 $Y2=0
cc_715 N_A_339_537#_c_811_n N_A_1875_543#_c_1329_n 0.00397771f $X=9.905 $Y=2.085
+ $X2=0 $Y2=0
cc_716 N_A_339_537#_c_826_n N_A_1875_543#_c_1341_n 0.0128062f $X=9.84 $Y=2.035
+ $X2=0 $Y2=0
cc_717 N_A_339_537#_c_828_n N_A_1875_543#_c_1341_n 0.00839426f $X=9.79 $Y=2.27
+ $X2=0 $Y2=0
cc_718 N_A_339_537#_M1027_g N_VPWR_c_1519_n 0.00323622f $X=10.02 $Y=2.925 $X2=0
+ $Y2=0
cc_719 N_A_339_537#_M1027_g N_VPWR_c_1528_n 0.0156697f $X=10.02 $Y=2.925 $X2=0
+ $Y2=0
cc_720 N_A_339_537#_c_814_n N_VPWR_c_1528_n 0.0174343f $X=1.835 $Y=2.83 $X2=0
+ $Y2=0
cc_721 N_A_339_537#_c_815_n N_VPWR_c_1528_n 0.00500435f $X=4.34 $Y=2.835 $X2=0
+ $Y2=0
cc_722 N_A_339_537#_c_816_n N_VPWR_c_1528_n 0.0176075f $X=4.34 $Y=2.835 $X2=0
+ $Y2=0
cc_723 N_A_339_537#_c_814_n N_A_452_632#_c_1634_n 0.0384542f $X=1.835 $Y=2.83
+ $X2=0 $Y2=0
cc_724 N_A_339_537#_c_820_n N_A_452_632#_c_1635_n 0.0176538f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_725 N_A_339_537#_c_814_n N_A_452_632#_c_1636_n 0.0115781f $X=1.835 $Y=2.83
+ $X2=0 $Y2=0
cc_726 N_A_339_537#_c_820_n N_A_452_632#_c_1636_n 0.0066903f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_727 N_A_339_537#_c_821_n N_A_452_632#_c_1636_n 0.00199723f $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_728 N_A_339_537#_c_824_n N_A_452_632#_c_1636_n 8.19979e-19 $X=2.16 $Y=2.035
+ $X2=0 $Y2=0
cc_729 N_A_339_537#_c_818_n N_A_452_632#_c_1637_n 0.010882f $X=4.34 $Y=2.67
+ $X2=15.12 $Y2=0
cc_730 N_A_339_537#_c_815_n N_A_452_632#_c_1638_n 0.0111344f $X=4.34 $Y=2.835
+ $X2=0 $Y2=0
cc_731 N_A_339_537#_c_816_n N_A_452_632#_c_1638_n 0.00326424f $X=4.34 $Y=2.835
+ $X2=0 $Y2=0
cc_732 N_A_339_537#_c_818_n N_A_452_632#_c_1632_n 0.0235843f $X=4.34 $Y=2.67
+ $X2=0 $Y2=0
cc_733 N_A_339_537#_c_860_n N_A_452_632#_c_1632_n 0.0154442f $X=4.45 $Y=2.035
+ $X2=0 $Y2=0
cc_734 N_A_339_537#_c_820_n N_A_452_632#_c_1632_n 0.0233075f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_735 N_A_339_537#_c_823_n N_A_452_632#_c_1632_n 4.87179e-19 $X=4.705 $Y=2.035
+ $X2=0 $Y2=0
cc_736 N_A_339_537#_c_820_n N_A_452_632#_c_1640_n 0.0023597f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_737 N_A_339_537#_c_815_n N_A_452_632#_c_1641_n 0.0133613f $X=4.34 $Y=2.835
+ $X2=0 $Y2=0
cc_738 N_A_339_537#_c_816_n N_A_452_632#_c_1641_n 0.00142073f $X=4.34 $Y=2.835
+ $X2=0 $Y2=0
cc_739 N_A_339_537#_c_806_n N_VGND_c_1708_n 0.0360269f $X=1.855 $Y=0.745 $X2=0
+ $Y2=0
cc_740 N_A_339_537#_c_806_n N_VGND_c_1710_n 0.0604113f $X=1.855 $Y=0.745 $X2=0
+ $Y2=0
cc_741 N_A_339_537#_c_824_n N_VGND_c_1710_n 0.00184466f $X=2.16 $Y=2.035 $X2=0
+ $Y2=0
cc_742 N_A_339_537#_c_804_n N_VGND_c_1718_n 0.0234259f $X=9.195 $Y=1.395 $X2=0
+ $Y2=0
cc_743 N_A_339_537#_c_806_n N_VGND_c_1718_n 0.0309537f $X=1.855 $Y=0.745 $X2=0
+ $Y2=0
cc_744 N_A_1119_506#_c_1012_n N_A_921_632#_M1022_g 0.0390936f $X=8.57 $Y=2.26
+ $X2=0 $Y2=0
cc_745 N_A_1119_506#_c_1023_n N_A_921_632#_M1022_g 0.0319393f $X=8.735 $Y=2.84
+ $X2=0 $Y2=0
cc_746 N_A_1119_506#_c_1005_n N_A_921_632#_M1022_g 0.00518457f $X=8.77 $Y=2.175
+ $X2=0 $Y2=0
cc_747 N_A_1119_506#_c_1030_n N_A_921_632#_M1022_g 0.00284694f $X=8.735 $Y=2.26
+ $X2=0 $Y2=0
cc_748 N_A_1119_506#_c_1048_n N_A_921_632#_c_1097_n 0.0100123f $X=8.805 $Y=0.7
+ $X2=0 $Y2=0
cc_749 N_A_1119_506#_c_1005_n N_A_921_632#_c_1097_n 0.00175914f $X=8.77 $Y=2.175
+ $X2=0 $Y2=0
cc_750 N_A_1119_506#_c_1006_n N_A_921_632#_c_1097_n 0.00319898f $X=8.805
+ $Y=1.325 $X2=0 $Y2=0
cc_751 N_A_1119_506#_c_1003_n N_A_921_632#_c_1099_n 0.00484224f $X=5.927
+ $Y=1.395 $X2=0 $Y2=0
cc_752 N_A_1119_506#_c_1002_n N_A_921_632#_c_1100_n 0.00901906f $X=5.927
+ $Y=1.657 $X2=0 $Y2=0
cc_753 N_A_1119_506#_c_1042_n N_A_921_632#_c_1100_n 0.0240295f $X=6.005 $Y=1.915
+ $X2=0 $Y2=0
cc_754 N_A_1119_506#_c_1074_p N_A_921_632#_c_1100_n 0.012969f $X=6.17 $Y=2.26
+ $X2=0 $Y2=0
cc_755 N_A_1119_506#_c_1002_n N_A_921_632#_c_1101_n 0.031622f $X=5.927 $Y=1.657
+ $X2=0 $Y2=0
cc_756 N_A_1119_506#_c_1042_n N_A_921_632#_c_1101_n 0.0218043f $X=6.005 $Y=1.915
+ $X2=0 $Y2=0
cc_757 N_A_1119_506#_c_1012_n N_A_921_632#_c_1101_n 0.00575138f $X=8.57 $Y=2.26
+ $X2=0 $Y2=0
cc_758 N_A_1119_506#_c_1010_n N_A_921_632#_c_1111_n 0.0177094f $X=5.892 $Y=3.03
+ $X2=0 $Y2=0
cc_759 N_A_1119_506#_c_1004_n N_A_921_632#_c_1111_n 0.00856422f $X=6.005
+ $Y=1.915 $X2=0 $Y2=0
cc_760 N_A_1119_506#_c_1012_n N_A_921_632#_c_1111_n 0.0730271f $X=8.57 $Y=2.26
+ $X2=0 $Y2=0
cc_761 N_A_1119_506#_c_1074_p N_A_921_632#_c_1111_n 0.0223051f $X=6.17 $Y=2.26
+ $X2=0 $Y2=0
cc_762 N_A_1119_506#_c_1003_n N_A_921_632#_c_1102_n 7.66324e-19 $X=5.927
+ $Y=1.395 $X2=0 $Y2=0
cc_763 N_A_1119_506#_c_1010_n N_A_921_632#_c_1114_n 0.00481137f $X=5.892 $Y=3.03
+ $X2=0 $Y2=0
cc_764 N_A_1119_506#_c_1004_n N_A_921_632#_c_1114_n 0.00901906f $X=6.005
+ $Y=1.915 $X2=0 $Y2=0
cc_765 N_A_1119_506#_c_1012_n N_A_921_632#_c_1104_n 0.00180572f $X=8.57 $Y=2.26
+ $X2=0 $Y2=0
cc_766 N_A_1119_506#_c_1005_n N_A_921_632#_c_1104_n 0.0155852f $X=8.77 $Y=2.175
+ $X2=0 $Y2=0
cc_767 N_A_1119_506#_c_1030_n N_A_921_632#_c_1104_n 0.00193547f $X=8.735 $Y=2.26
+ $X2=0 $Y2=0
cc_768 N_A_1119_506#_c_1048_n N_A_1875_543#_c_1364_n 0.00586146f $X=8.805 $Y=0.7
+ $X2=0 $Y2=0
cc_769 N_A_1119_506#_c_1048_n N_A_1875_543#_c_1328_n 0.0180396f $X=8.805 $Y=0.7
+ $X2=0 $Y2=0
cc_770 N_A_1119_506#_M1026_g N_VPWR_c_1513_n 0.0353437f $X=5.845 $Y=3.37 $X2=0
+ $Y2=0
cc_771 N_A_1119_506#_c_1010_n N_VPWR_c_1513_n 5.24152e-19 $X=5.892 $Y=3.03 $X2=0
+ $Y2=0
cc_772 N_A_1119_506#_M1022_d N_VPWR_c_1516_n 0.00487614f $X=8.595 $Y=2.715 $X2=0
+ $Y2=0
cc_773 N_A_1119_506#_M1022_d N_VPWR_c_1528_n 0.00242411f $X=8.595 $Y=2.715 $X2=0
+ $Y2=0
cc_774 N_A_1119_506#_M1026_g N_VPWR_c_1528_n 0.00499575f $X=5.845 $Y=3.37 $X2=0
+ $Y2=0
cc_775 N_A_1119_506#_c_1003_n N_VGND_c_1718_n 0.00509893f $X=5.927 $Y=1.395
+ $X2=0 $Y2=0
cc_776 N_A_1119_506#_c_1048_n N_VGND_c_1718_n 0.0228585f $X=8.805 $Y=0.7 $X2=0
+ $Y2=0
cc_777 N_A_921_632#_M1022_g N_VPWR_c_1516_n 0.0232236f $X=8.345 $Y=3.215 $X2=0
+ $Y2=0
cc_778 N_A_921_632#_M1022_g N_VPWR_c_1528_n 0.00752887f $X=8.345 $Y=3.215 $X2=0
+ $Y2=0
cc_779 N_A_921_632#_c_1112_n N_VPWR_c_1528_n 0.0227758f $X=7.095 $Y=3.325 $X2=0
+ $Y2=0
cc_780 N_A_921_632#_c_1132_n N_VPWR_c_1528_n 0.0215818f $X=4.745 $Y=3.325 $X2=0
+ $Y2=0
cc_781 N_A_921_632#_c_1132_n N_A_452_632#_c_1638_n 0.00374485f $X=4.745 $Y=3.325
+ $X2=0 $Y2=0
cc_782 N_A_921_632#_c_1113_n N_A_452_632#_c_1638_n 0.00502812f $X=4.745 $Y=3.2
+ $X2=0 $Y2=0
cc_783 N_A_921_632#_c_1102_n N_A_452_632#_c_1631_n 0.01409f $X=4.815 $Y=1.075
+ $X2=0 $Y2=0
cc_784 N_A_921_632#_c_1097_n N_VGND_c_1712_n 0.0127791f $X=8.415 $Y=1.395 $X2=0
+ $Y2=0
cc_785 N_A_921_632#_c_1097_n N_VGND_c_1718_n 0.0156107f $X=8.415 $Y=1.395 $X2=0
+ $Y2=0
cc_786 N_A_921_632#_c_1154_n N_VGND_c_1718_n 0.00428084f $X=5.49 $Y=1.16 $X2=0
+ $Y2=0
cc_787 N_A_921_632#_c_1102_n N_VGND_c_1718_n 0.00255615f $X=4.815 $Y=1.075 $X2=0
+ $Y2=0
cc_788 N_A_921_632#_c_1154_n A_1091_173# 0.00161044f $X=5.49 $Y=1.16 $X2=0 $Y2=0
cc_789 N_A_2096_417#_c_1235_n N_A_1875_543#_M1023_g 0.00880415f $X=12.785
+ $Y=0.745 $X2=0 $Y2=0
cc_790 N_A_2096_417#_c_1237_n N_A_1875_543#_M1023_g 0.0245645f $X=12.732
+ $Y=1.835 $X2=0 $Y2=0
cc_791 N_A_2096_417#_c_1238_n N_A_1875_543#_M1023_g 0.00510414f $X=12.785
+ $Y=0.995 $X2=0 $Y2=0
cc_792 N_A_2096_417#_c_1237_n N_A_1875_543#_c_1324_n 0.013597f $X=12.732
+ $Y=1.835 $X2=0.24 $Y2=0
cc_793 N_A_2096_417#_c_1247_n N_A_1875_543#_c_1324_n 0.00907295f $X=12.76
+ $Y=2.535 $X2=0.24 $Y2=0
cc_794 N_A_2096_417#_c_1238_n N_A_1875_543#_c_1324_n 0.00299261f $X=12.785
+ $Y=0.995 $X2=0.24 $Y2=0
cc_795 N_A_2096_417#_c_1282_p N_A_1875_543#_c_1324_n 0.00837999f $X=12.732
+ $Y=1.92 $X2=0.24 $Y2=0
cc_796 N_A_2096_417#_c_1237_n N_A_1875_543#_M1015_g 0.00155468f $X=12.732
+ $Y=1.835 $X2=0 $Y2=0
cc_797 N_A_2096_417#_c_1238_n N_A_1875_543#_M1015_g 0.00249326f $X=12.785
+ $Y=0.995 $X2=0 $Y2=0
cc_798 N_A_2096_417#_c_1234_n N_A_1875_543#_c_1326_n 0.0384835f $X=12.62 $Y=1.92
+ $X2=0 $Y2=0
cc_799 N_A_2096_417#_c_1237_n N_A_1875_543#_c_1326_n 0.00754828f $X=12.732
+ $Y=1.835 $X2=0 $Y2=0
cc_800 N_A_2096_417#_c_1282_p N_A_1875_543#_c_1326_n 9.9512e-19 $X=12.732
+ $Y=1.92 $X2=0 $Y2=0
cc_801 N_A_2096_417#_M1021_g N_A_1875_543#_c_1338_n 6.95068e-19 $X=10.73
+ $Y=2.925 $X2=0 $Y2=0
cc_802 N_A_2096_417#_M1031_g N_A_1875_543#_c_1351_n 7.33647e-19 $X=10.905
+ $Y=0.745 $X2=0 $Y2=0
cc_803 N_A_2096_417#_c_1242_n N_A_1875_543#_c_1339_n 0.00662553f $X=10.817
+ $Y=2.585 $X2=0 $Y2=0
cc_804 N_A_2096_417#_c_1242_n N_A_1875_543#_c_1329_n 0.00898266f $X=10.817
+ $Y=2.585 $X2=0 $Y2=0
cc_805 N_A_2096_417#_c_1249_n N_A_1875_543#_c_1329_n 0.0254288f $X=10.97
+ $Y=1.555 $X2=0 $Y2=0
cc_806 N_A_2096_417#_c_1293_p N_A_1875_543#_c_1329_n 0.0117859f $X=11.135
+ $Y=1.92 $X2=0 $Y2=0
cc_807 N_A_2096_417#_M1031_g N_A_1875_543#_c_1329_n 0.0198821f $X=10.905
+ $Y=0.745 $X2=0 $Y2=0
cc_808 N_A_2096_417#_c_1242_n N_A_1875_543#_c_1341_n 0.00625697f $X=10.817
+ $Y=2.585 $X2=0 $Y2=0
cc_809 N_A_2096_417#_c_1242_n N_A_1875_543#_c_1342_n 0.0337751f $X=10.817
+ $Y=2.585 $X2=0 $Y2=0
cc_810 N_A_2096_417#_c_1234_n N_A_1875_543#_c_1342_n 0.0917351f $X=12.62 $Y=1.92
+ $X2=0 $Y2=0
cc_811 N_A_2096_417#_c_1293_p N_A_1875_543#_c_1342_n 0.0236209f $X=11.135
+ $Y=1.92 $X2=0 $Y2=0
cc_812 N_A_2096_417#_c_1245_n N_A_1875_543#_c_1342_n 0.0266022f $X=12.675
+ $Y=2.62 $X2=0 $Y2=0
cc_813 N_A_2096_417#_c_1246_n N_A_1875_543#_c_1342_n 0.0199673f $X=12.09 $Y=2.62
+ $X2=0 $Y2=0
cc_814 N_A_2096_417#_c_1247_n N_A_1875_543#_c_1342_n 0.0128523f $X=12.76
+ $Y=2.535 $X2=0 $Y2=0
cc_815 N_A_2096_417#_c_1244_n N_A_1875_543#_c_1343_n 7.39752e-19 $X=12.005
+ $Y=2.925 $X2=0 $Y2=0
cc_816 N_A_2096_417#_c_1245_n N_A_1875_543#_c_1343_n 0.0322257f $X=12.675
+ $Y=2.62 $X2=0 $Y2=0
cc_817 N_A_2096_417#_c_1247_n N_A_1875_543#_c_1343_n 0.0178294f $X=12.76
+ $Y=2.535 $X2=0 $Y2=0
cc_818 N_A_2096_417#_c_1237_n N_A_2649_207#_c_1457_n 0.0231612f $X=12.732
+ $Y=1.835 $X2=15.12 $Y2=0
cc_819 N_A_2096_417#_c_1237_n N_A_2649_207#_c_1458_n 0.0059307f $X=12.732
+ $Y=1.835 $X2=0 $Y2=0
cc_820 N_A_2096_417#_c_1245_n N_A_2649_207#_c_1465_n 0.0066962f $X=12.675
+ $Y=2.62 $X2=7.68 $Y2=0.057
cc_821 N_A_2096_417#_c_1247_n N_A_2649_207#_c_1465_n 0.0183025f $X=12.76
+ $Y=2.535 $X2=7.68 $Y2=0.057
cc_822 N_A_2096_417#_c_1237_n N_A_2649_207#_c_1472_n 0.00512676f $X=12.732
+ $Y=1.835 $X2=0 $Y2=0
cc_823 N_A_2096_417#_c_1282_p N_A_2649_207#_c_1472_n 0.00593551f $X=12.732
+ $Y=1.92 $X2=0 $Y2=0
cc_824 N_A_2096_417#_M1021_g N_VPWR_c_1519_n 0.0581985f $X=10.73 $Y=2.925 $X2=0
+ $Y2=0
cc_825 N_A_2096_417#_c_1242_n N_VPWR_c_1519_n 0.00572618f $X=10.817 $Y=2.585
+ $X2=0 $Y2=0
cc_826 N_A_2096_417#_c_1244_n N_VPWR_c_1519_n 0.018164f $X=12.005 $Y=2.925 $X2=0
+ $Y2=0
cc_827 N_A_2096_417#_c_1246_n N_VPWR_c_1519_n 0.00125202f $X=12.09 $Y=2.62 $X2=0
+ $Y2=0
cc_828 N_A_2096_417#_c_1244_n N_VPWR_c_1522_n 0.0131078f $X=12.005 $Y=2.925
+ $X2=0 $Y2=0
cc_829 N_A_2096_417#_c_1245_n N_VPWR_c_1522_n 0.0420395f $X=12.675 $Y=2.62 $X2=0
+ $Y2=0
cc_830 N_A_2096_417#_c_1244_n N_VPWR_c_1528_n 0.0126975f $X=12.005 $Y=2.925
+ $X2=0 $Y2=0
cc_831 N_A_2096_417#_c_1235_n N_VGND_c_1714_n 0.0117406f $X=12.785 $Y=0.745
+ $X2=0 $Y2=0
cc_832 N_A_2096_417#_M1031_g N_VGND_c_1714_n 0.00955903f $X=10.905 $Y=0.745
+ $X2=0 $Y2=0
cc_833 N_A_2096_417#_c_1235_n N_VGND_c_1718_n 0.0352665f $X=12.785 $Y=0.745
+ $X2=0 $Y2=0
cc_834 N_A_2096_417#_M1031_g N_VGND_c_1718_n 0.0110498f $X=10.905 $Y=0.745 $X2=0
+ $Y2=0
cc_835 N_A_1875_543#_M1015_g N_A_2649_207#_M1002_g 0.0145305f $X=13.78 $Y=1.245
+ $X2=0 $Y2=0
cc_836 N_A_1875_543#_M1019_g N_A_2649_207#_M1010_g 0.019729f $X=13.82 $Y=2.59
+ $X2=0 $Y2=0
cc_837 N_A_1875_543#_M1023_g N_A_2649_207#_c_1457_n 0.0022681f $X=12.395
+ $Y=0.745 $X2=15.12 $Y2=0
cc_838 N_A_1875_543#_M1015_g N_A_2649_207#_c_1457_n 0.00715068f $X=13.78
+ $Y=1.245 $X2=15.12 $Y2=0
cc_839 N_A_1875_543#_c_1324_n N_A_2649_207#_c_1458_n 0.00594043f $X=13.53
+ $Y=1.835 $X2=0 $Y2=0
cc_840 N_A_1875_543#_M1015_g N_A_2649_207#_c_1458_n 0.00553556f $X=13.78
+ $Y=1.245 $X2=0 $Y2=0
cc_841 N_A_1875_543#_c_1327_n N_A_2649_207#_c_1458_n 0.00401739f $X=13.8
+ $Y=1.835 $X2=0 $Y2=0
cc_842 N_A_1875_543#_c_1324_n N_A_2649_207#_c_1465_n 0.0066977f $X=13.53
+ $Y=1.835 $X2=7.68 $Y2=0.057
cc_843 N_A_1875_543#_M1019_g N_A_2649_207#_c_1465_n 0.0240803f $X=13.82 $Y=2.59
+ $X2=7.68 $Y2=0.057
cc_844 N_A_1875_543#_c_1327_n N_A_2649_207#_c_1465_n 0.00390596f $X=13.8
+ $Y=1.835 $X2=7.68 $Y2=0.057
cc_845 N_A_1875_543#_c_1327_n N_A_2649_207#_c_1459_n 0.0430166f $X=13.8 $Y=1.835
+ $X2=0 $Y2=0
cc_846 N_A_1875_543#_c_1327_n N_A_2649_207#_c_1460_n 0.0239562f $X=13.8 $Y=1.835
+ $X2=0 $Y2=0
cc_847 N_A_1875_543#_c_1324_n N_A_2649_207#_c_1461_n 0.00578003f $X=13.53
+ $Y=1.835 $X2=0 $Y2=0
cc_848 N_A_1875_543#_M1015_g N_A_2649_207#_c_1461_n 0.00386717f $X=13.78
+ $Y=1.245 $X2=0 $Y2=0
cc_849 N_A_1875_543#_c_1324_n N_A_2649_207#_c_1472_n 0.0144101f $X=13.53
+ $Y=1.835 $X2=0 $Y2=0
cc_850 N_A_1875_543#_c_1327_n N_A_2649_207#_c_1472_n 0.00409644f $X=13.8
+ $Y=1.835 $X2=0 $Y2=0
cc_851 N_A_1875_543#_c_1338_n N_VPWR_c_1519_n 0.00858473f $X=10.135 $Y=2.76
+ $X2=0 $Y2=0
cc_852 N_A_1875_543#_c_1341_n N_VPWR_c_1519_n 0.0459993f $X=10.6 $Y=2.27 $X2=0
+ $Y2=0
cc_853 N_A_1875_543#_M1019_g N_VPWR_c_1522_n 0.00246615f $X=13.82 $Y=2.59 $X2=0
+ $Y2=0
cc_854 N_A_1875_543#_c_1343_n N_VPWR_c_1522_n 0.0340077f $X=12.33 $Y=2.27 $X2=0
+ $Y2=0
cc_855 N_A_1875_543#_M1019_g N_VPWR_c_1525_n 0.0637647f $X=13.82 $Y=2.59 $X2=0
+ $Y2=0
cc_856 N_A_1875_543#_M1007_d N_VPWR_c_1528_n 0.00221032f $X=9.375 $Y=2.715 $X2=0
+ $Y2=0
cc_857 N_A_1875_543#_M1019_g N_VPWR_c_1528_n 0.00584154f $X=13.82 $Y=2.59 $X2=0
+ $Y2=0
cc_858 N_A_1875_543#_c_1335_n N_VPWR_c_1528_n 0.0454876f $X=9.515 $Y=3.215 $X2=0
+ $Y2=0
cc_859 N_A_1875_543#_c_1338_n N_VPWR_c_1528_n 0.0197014f $X=10.135 $Y=2.76 $X2=0
+ $Y2=0
cc_860 N_A_1875_543#_c_1343_n N_VPWR_c_1528_n 0.00394878f $X=12.33 $Y=2.27 $X2=0
+ $Y2=0
cc_861 N_A_1875_543#_M1023_g N_VGND_c_1714_n 0.00760888f $X=12.395 $Y=0.745
+ $X2=0 $Y2=0
cc_862 N_A_1875_543#_M1015_g N_VGND_c_1716_n 0.0481833f $X=13.78 $Y=1.245 $X2=0
+ $Y2=0
cc_863 N_A_1875_543#_c_1327_n N_VGND_c_1716_n 0.00120691f $X=13.8 $Y=1.835 $X2=0
+ $Y2=0
cc_864 N_A_1875_543#_M1023_g N_VGND_c_1718_n 0.0326394f $X=12.395 $Y=0.745 $X2=0
+ $Y2=0
cc_865 N_A_1875_543#_M1015_g N_VGND_c_1718_n 0.00608654f $X=13.78 $Y=1.245 $X2=0
+ $Y2=0
cc_866 N_A_1875_543#_c_1364_n N_VGND_c_1718_n 0.0228821f $X=9.595 $Y=0.785 $X2=0
+ $Y2=0
cc_867 N_A_1875_543#_c_1351_n N_VGND_c_1718_n 0.0423573f $X=10.43 $Y=0.7 $X2=0
+ $Y2=0
cc_868 N_A_1875_543#_c_1351_n A_2089_107# 4.80934e-19 $X=10.43 $Y=0.7 $X2=0
+ $Y2=0
cc_869 N_A_2649_207#_c_1465_n N_VPWR_c_1522_n 0.00983841f $X=13.43 $Y=2.34 $X2=0
+ $Y2=0
cc_870 N_A_2649_207#_M1010_g N_VPWR_c_1525_n 0.0677668f $X=14.695 $Y=2.965 $X2=0
+ $Y2=0
cc_871 N_A_2649_207#_c_1465_n N_VPWR_c_1525_n 0.0602601f $X=13.43 $Y=2.34 $X2=0
+ $Y2=0
cc_872 N_A_2649_207#_c_1459_n N_VPWR_c_1525_n 0.0718006f $X=14.555 $Y=1.84 $X2=0
+ $Y2=0
cc_873 N_A_2649_207#_c_1460_n N_VPWR_c_1525_n 0.00210918f $X=14.555 $Y=1.84
+ $X2=0 $Y2=0
cc_874 N_A_2649_207#_M1010_g N_VPWR_c_1528_n 0.0117682f $X=14.695 $Y=2.965 $X2=0
+ $Y2=0
cc_875 N_A_2649_207#_c_1465_n N_VPWR_c_1528_n 0.0108564f $X=13.43 $Y=2.34 $X2=0
+ $Y2=0
cc_876 N_A_2649_207#_M1002_g N_Q_c_1696_n 0.0252289f $X=14.675 $Y=1.08 $X2=0
+ $Y2=0
cc_877 N_A_2649_207#_M1010_g N_Q_c_1696_n 0.0360118f $X=14.695 $Y=2.965 $X2=0
+ $Y2=0
cc_878 N_A_2649_207#_c_1459_n N_Q_c_1696_n 0.0250299f $X=14.555 $Y=1.84 $X2=0
+ $Y2=0
cc_879 N_A_2649_207#_c_1460_n N_Q_c_1696_n 0.0250892f $X=14.555 $Y=1.84 $X2=0
+ $Y2=0
cc_880 N_A_2649_207#_M1002_g N_VGND_c_1716_n 0.0529832f $X=14.675 $Y=1.08 $X2=0
+ $Y2=0
cc_881 N_A_2649_207#_c_1457_n N_VGND_c_1716_n 0.0379082f $X=13.39 $Y=1.245 $X2=0
+ $Y2=0
cc_882 N_A_2649_207#_c_1459_n N_VGND_c_1716_n 0.0753111f $X=14.555 $Y=1.84 $X2=0
+ $Y2=0
cc_883 N_A_2649_207#_c_1460_n N_VGND_c_1716_n 0.00154364f $X=14.555 $Y=1.84
+ $X2=0 $Y2=0
cc_884 N_A_2649_207#_M1002_g N_VGND_c_1718_n 0.0140081f $X=14.675 $Y=1.08 $X2=0
+ $Y2=0
cc_885 N_A_2649_207#_c_1457_n N_VGND_c_1718_n 0.0151966f $X=13.39 $Y=1.245 $X2=0
+ $Y2=0
cc_886 N_VPWR_c_1528_n N_A_452_632#_M1024_s 7.65036e-19 $X=14.605 $Y=3.59 $X2=0
+ $Y2=0
cc_887 N_VPWR_c_1528_n N_A_452_632#_M1009_d 0.00297536f $X=14.605 $Y=3.59 $X2=0
+ $Y2=0
cc_888 N_VPWR_c_1528_n N_A_452_632#_c_1634_n 0.0172954f $X=14.605 $Y=3.59
+ $X2=0.24 $Y2=4.07
cc_889 N_VPWR_c_1528_n N_A_452_632#_c_1635_n 0.0113657f $X=14.605 $Y=3.59
+ $X2=15.12 $Y2=4.07
cc_890 N_VPWR_c_1528_n N_A_452_632#_c_1638_n 0.0114742f $X=14.605 $Y=3.59
+ $X2=7.68 $Y2=4.013
cc_891 N_VPWR_c_1513_n A_1077_632# 0.00356654f $X=6.285 $Y=3.59 $X2=0 $Y2=3.985
cc_892 N_VPWR_c_1528_n A_1077_632# 7.4516e-19 $X=14.605 $Y=3.59 $X2=0 $Y2=3.985
cc_893 N_VPWR_c_1525_n N_Q_c_1696_n 0.112775f $X=14.305 $Y=2.36 $X2=7.68
+ $Y2=4.07
cc_894 N_VPWR_c_1528_n N_Q_c_1696_n 0.0424118f $X=14.605 $Y=3.59 $X2=7.68
+ $Y2=4.07
cc_895 N_A_452_632#_c_1631_n N_VGND_c_1718_n 0.00217159f $X=4.035 $Y=1.075 $X2=0
+ $Y2=0
cc_896 N_Q_c_1696_n N_VGND_c_1716_n 0.0547104f $X=15.065 $Y=0.83 $X2=0 $Y2=0
cc_897 N_Q_c_1696_n N_VGND_c_1718_n 0.0148422f $X=15.065 $Y=0.83 $X2=0 $Y2=0
cc_898 N_VGND_c_1718_n A_2089_107# 0.00225203f $X=14.57 $Y=0.48 $X2=0 $Y2=0
cc_899 N_VGND_c_1714_n A_2387_107# 0.00891833f $X=11.965 $Y=0.48 $X2=0 $Y2=0
cc_900 N_VGND_c_1718_n A_2387_107# 0.00271077f $X=14.57 $Y=0.48 $X2=0 $Y2=0
