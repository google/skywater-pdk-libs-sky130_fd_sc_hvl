* File: sky130_fd_sc_hvl__buf_4.pxi.spice
* Created: Wed Sep  2 09:04:20 2020
* 
x_PM_SKY130_FD_SC_HVL__BUF_4%VNB N_VNB_M1000_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__BUF_4%VNB
x_PM_SKY130_FD_SC_HVL__BUF_4%VPB N_VPB_M1004_b VPB N_VPB_c_35_p VPB
+ PM_SKY130_FD_SC_HVL__BUF_4%VPB
x_PM_SKY130_FD_SC_HVL__BUF_4%A_149_81# N_A_149_81#_M1007_d N_A_149_81#_M1001_d
+ N_A_149_81#_M1000_g N_A_149_81#_M1004_g N_A_149_81#_M1002_g
+ N_A_149_81#_M1006_g N_A_149_81#_M1003_g N_A_149_81#_M1008_g
+ N_A_149_81#_M1005_g N_A_149_81#_M1009_g N_A_149_81#_c_121_p N_A_149_81#_c_79_n
+ N_A_149_81#_c_80_n N_A_149_81#_c_82_n N_A_149_81#_c_106_p N_A_149_81#_c_83_n
+ N_A_149_81#_c_84_n PM_SKY130_FD_SC_HVL__BUF_4%A_149_81#
x_PM_SKY130_FD_SC_HVL__BUF_4%A A N_A_M1007_g N_A_c_187_n N_A_M1001_g
+ PM_SKY130_FD_SC_HVL__BUF_4%A
x_PM_SKY130_FD_SC_HVL__BUF_4%VPWR N_VPWR_M1004_d N_VPWR_M1006_d N_VPWR_M1009_d
+ VPWR N_VPWR_c_196_n N_VPWR_c_199_n N_VPWR_c_202_n N_VPWR_c_205_n
+ PM_SKY130_FD_SC_HVL__BUF_4%VPWR
x_PM_SKY130_FD_SC_HVL__BUF_4%X N_X_M1000_s N_X_M1003_s N_X_M1004_s N_X_M1008_s
+ N_X_c_237_n N_X_c_239_n N_X_c_257_n N_X_c_245_n N_X_c_240_n N_X_c_248_n
+ N_X_c_241_n N_X_c_249_n N_X_c_243_n N_X_c_244_n X X
+ PM_SKY130_FD_SC_HVL__BUF_4%X
x_PM_SKY130_FD_SC_HVL__BUF_4%VGND N_VGND_M1000_d N_VGND_M1002_d N_VGND_M1005_d
+ VGND N_VGND_c_301_n N_VGND_c_303_n N_VGND_c_305_n N_VGND_c_307_n
+ PM_SKY130_FD_SC_HVL__BUF_4%VGND
cc_1 N_VNB_M1000_b N_A_149_81#_M1000_g 0.0480486f $X=-0.33 $Y=-0.265 $X2=0.995
+ $Y2=0.91
cc_2 N_VNB_c_2_p N_A_149_81#_M1000_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.995 $Y2=0.91
cc_3 N_VNB_M1000_b N_A_149_81#_M1002_g 0.0405519f $X=-0.33 $Y=-0.265 $X2=1.775
+ $Y2=0.91
cc_4 N_VNB_c_2_p N_A_149_81#_M1002_g 5.86481e-19 $X=0.24 $Y=0 $X2=1.775 $Y2=0.91
cc_5 N_VNB_M1000_b N_A_149_81#_M1003_g 0.0422505f $X=-0.33 $Y=-0.265 $X2=2.555
+ $Y2=0.91
cc_6 N_VNB_c_2_p N_A_149_81#_M1003_g 9.58849e-19 $X=0.24 $Y=0 $X2=2.555 $Y2=0.91
cc_7 N_VNB_M1000_b N_A_149_81#_M1005_g 0.0416851f $X=-0.33 $Y=-0.265 $X2=3.335
+ $Y2=0.91
cc_8 N_VNB_c_2_p N_A_149_81#_M1005_g 5.86481e-19 $X=0.24 $Y=0 $X2=3.335 $Y2=0.91
cc_9 N_VNB_M1000_b N_A_149_81#_c_79_n 0.0107068f $X=-0.33 $Y=-0.265 $X2=4.34
+ $Y2=1.51
cc_10 N_VNB_M1000_b N_A_149_81#_c_80_n 0.0440426f $X=-0.33 $Y=-0.265 $X2=4.505
+ $Y2=0.66
cc_11 N_VNB_c_2_p N_A_149_81#_c_80_n 8.20017e-19 $X=0.24 $Y=0 $X2=4.505 $Y2=0.66
cc_12 N_VNB_M1000_b N_A_149_81#_c_82_n 0.0146238f $X=-0.33 $Y=-0.265 $X2=4.505
+ $Y2=2.34
cc_13 N_VNB_M1000_b N_A_149_81#_c_83_n 0.179178f $X=-0.33 $Y=-0.265 $X2=3.435
+ $Y2=1.64
cc_14 N_VNB_M1000_b N_A_149_81#_c_84_n 0.00994965f $X=-0.33 $Y=-0.265 $X2=4.505
+ $Y2=1.51
cc_15 N_VNB_M1000_b N_A_M1007_g 0.0918746f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_16 N_VNB_c_2_p N_A_M1007_g 9.58849e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_17 N_VNB_M1000_b N_X_c_237_n 0.00864253f $X=-0.33 $Y=-0.265 $X2=1.775
+ $Y2=1.415
cc_18 N_VNB_c_2_p N_X_c_237_n 6.32535e-19 $X=0.24 $Y=0 $X2=1.775 $Y2=1.415
cc_19 N_VNB_M1000_b N_X_c_239_n 3.66238e-19 $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_20 N_VNB_M1000_b N_X_c_240_n 0.00588496f $X=-0.33 $Y=-0.265 $X2=2.555
+ $Y2=0.91
cc_21 N_VNB_M1000_b N_X_c_241_n 0.00864253f $X=-0.33 $Y=-0.265 $X2=3.335
+ $Y2=1.415
cc_22 N_VNB_c_2_p N_X_c_241_n 6.32535e-19 $X=0.24 $Y=0 $X2=3.335 $Y2=1.415
cc_23 N_VNB_M1000_b N_X_c_243_n 7.98126e-19 $X=-0.33 $Y=-0.265 $X2=3.43 $Y2=1.64
cc_24 N_VNB_M1000_b N_X_c_244_n 0.0273739f $X=-0.33 $Y=-0.265 $X2=1.735 $Y2=1.64
cc_25 N_VNB_M1000_b N_VGND_c_301_n 0.0999516f $X=-0.33 $Y=-0.265 $X2=0.995
+ $Y2=2.965
cc_26 N_VNB_c_2_p N_VGND_c_301_n 0.00269049f $X=0.24 $Y=0 $X2=0.995 $Y2=2.965
cc_27 N_VNB_M1000_b N_VGND_c_303_n 0.0466622f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_28 N_VNB_c_2_p N_VGND_c_303_n 0.00269176f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_29 N_VNB_M1000_b N_VGND_c_305_n 0.0468473f $X=-0.33 $Y=-0.265 $X2=3.335
+ $Y2=1.415
cc_30 N_VNB_c_2_p N_VGND_c_305_n 0.00269049f $X=0.24 $Y=0 $X2=3.335 $Y2=1.415
cc_31 N_VNB_M1000_b N_VGND_c_307_n 0.0841239f $X=-0.33 $Y=-0.265 $X2=3.335
+ $Y2=1.915
cc_32 N_VNB_c_2_p N_VGND_c_307_n 0.51328f $X=0.24 $Y=0 $X2=3.335 $Y2=1.915
cc_33 N_VPB_M1004_b N_A_149_81#_M1004_g 0.0610236f $X=-0.33 $Y=1.885 $X2=0.995
+ $Y2=2.965
cc_34 VPB N_A_149_81#_M1004_g 0.00970178f $X=0 $Y=3.955 $X2=0.995 $Y2=2.965
cc_35 N_VPB_c_35_p N_A_149_81#_M1004_g 0.0158814f $X=4.56 $Y=4.07 $X2=0.995
+ $Y2=2.965
cc_36 N_VPB_M1004_b N_A_149_81#_M1006_g 0.0483801f $X=-0.33 $Y=1.885 $X2=1.775
+ $Y2=2.965
cc_37 VPB N_A_149_81#_M1006_g 0.00970178f $X=0 $Y=3.955 $X2=1.775 $Y2=2.965
cc_38 N_VPB_c_35_p N_A_149_81#_M1006_g 0.0152133f $X=4.56 $Y=4.07 $X2=1.775
+ $Y2=2.965
cc_39 N_VPB_M1004_b N_A_149_81#_M1008_g 0.04781f $X=-0.33 $Y=1.885 $X2=2.555
+ $Y2=2.965
cc_40 VPB N_A_149_81#_M1008_g 0.00970178f $X=0 $Y=3.955 $X2=2.555 $Y2=2.965
cc_41 N_VPB_c_35_p N_A_149_81#_M1008_g 0.0158814f $X=4.56 $Y=4.07 $X2=2.555
+ $Y2=2.965
cc_42 N_VPB_M1004_b N_A_149_81#_M1009_g 0.0492445f $X=-0.33 $Y=1.885 $X2=3.335
+ $Y2=2.965
cc_43 VPB N_A_149_81#_M1009_g 0.00970178f $X=0 $Y=3.955 $X2=3.335 $Y2=2.965
cc_44 N_VPB_c_35_p N_A_149_81#_M1009_g 0.0158814f $X=4.56 $Y=4.07 $X2=3.335
+ $Y2=2.965
cc_45 N_VPB_M1004_b N_A_149_81#_c_82_n 0.0682168f $X=-0.33 $Y=1.885 $X2=4.505
+ $Y2=2.34
cc_46 VPB N_A_149_81#_c_82_n 7.60114e-19 $X=0 $Y=3.955 $X2=4.505 $Y2=2.34
cc_47 N_VPB_c_35_p N_A_149_81#_c_82_n 0.0131049f $X=4.56 $Y=4.07 $X2=4.505
+ $Y2=2.34
cc_48 N_VPB_M1004_b N_A_149_81#_c_83_n 0.020961f $X=-0.33 $Y=1.885 $X2=3.435
+ $Y2=1.64
cc_49 N_VPB_M1004_b N_A_M1007_g 0.05863f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_50 VPB N_A_M1007_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_51 N_VPB_c_35_p N_A_M1007_g 0.0152133f $X=4.56 $Y=4.07 $X2=0 $Y2=0
cc_52 N_VPB_M1004_b N_VPWR_c_196_n 0.0901534f $X=-0.33 $Y=1.885 $X2=0.995
+ $Y2=2.965
cc_53 VPB N_VPWR_c_196_n 0.00341542f $X=0 $Y=3.955 $X2=0.995 $Y2=2.965
cc_54 N_VPB_c_35_p N_VPWR_c_196_n 0.0489311f $X=4.56 $Y=4.07 $X2=0.995 $Y2=2.965
cc_55 N_VPB_M1004_b N_VPWR_c_199_n 0.00125033f $X=-0.33 $Y=1.885 $X2=2.555
+ $Y2=1.415
cc_56 VPB N_VPWR_c_199_n 0.00406397f $X=0 $Y=3.955 $X2=2.555 $Y2=1.415
cc_57 N_VPB_c_35_p N_VPWR_c_199_n 0.047451f $X=4.56 $Y=4.07 $X2=2.555 $Y2=1.415
cc_58 N_VPB_M1004_b N_VPWR_c_202_n 0.00125033f $X=-0.33 $Y=1.885 $X2=3.335
+ $Y2=0.91
cc_59 VPB N_VPWR_c_202_n 0.00406397f $X=0 $Y=3.955 $X2=3.335 $Y2=0.91
cc_60 N_VPB_c_35_p N_VPWR_c_202_n 0.047451f $X=4.56 $Y=4.07 $X2=3.335 $Y2=0.91
cc_61 N_VPB_M1004_b N_VPWR_c_205_n 0.0469352f $X=-0.33 $Y=1.885 $X2=1.735
+ $Y2=1.64
cc_62 VPB N_VPWR_c_205_n 0.509005f $X=0 $Y=3.955 $X2=1.735 $Y2=1.64
cc_63 N_VPB_c_35_p N_VPWR_c_205_n 0.0209143f $X=4.56 $Y=4.07 $X2=1.735 $Y2=1.64
cc_64 N_VPB_M1004_b N_X_c_245_n 0.00251996f $X=-0.33 $Y=1.885 $X2=1.775
+ $Y2=2.965
cc_65 VPB N_X_c_245_n 8.01732e-19 $X=0 $Y=3.955 $X2=1.775 $Y2=2.965
cc_66 N_VPB_c_35_p N_X_c_245_n 0.0130099f $X=4.56 $Y=4.07 $X2=1.775 $Y2=2.965
cc_67 N_VPB_M1004_b N_X_c_248_n 0.00447242f $X=-0.33 $Y=1.885 $X2=2.555
+ $Y2=1.915
cc_68 N_VPB_M1004_b N_X_c_249_n 0.00125033f $X=-0.33 $Y=1.885 $X2=3.335
+ $Y2=1.915
cc_69 VPB N_X_c_249_n 0.00108855f $X=0 $Y=3.955 $X2=3.335 $Y2=1.915
cc_70 N_VPB_c_35_p N_X_c_249_n 0.0171423f $X=4.56 $Y=4.07 $X2=3.335 $Y2=1.915
cc_71 N_A_149_81#_M1005_g N_A_M1007_g 0.0188315f $X=3.335 $Y=0.91 $X2=0 $Y2=0
cc_72 N_A_149_81#_M1009_g N_A_M1007_g 0.0251156f $X=3.335 $Y=2.965 $X2=0 $Y2=0
cc_73 N_A_149_81#_c_79_n N_A_M1007_g 0.0324363f $X=4.34 $Y=1.51 $X2=0 $Y2=0
cc_74 N_A_149_81#_c_80_n N_A_M1007_g 0.0260752f $X=4.505 $Y=0.66 $X2=0 $Y2=0
cc_75 N_A_149_81#_c_82_n N_A_M1007_g 0.0259732f $X=4.505 $Y=2.34 $X2=0 $Y2=0
cc_76 N_A_149_81#_c_106_p N_A_M1007_g 0.00101702f $X=3.515 $Y=1.51 $X2=0 $Y2=0
cc_77 N_A_149_81#_c_83_n N_A_M1007_g 0.030513f $X=3.435 $Y=1.64 $X2=0 $Y2=0
cc_78 N_A_149_81#_c_84_n N_A_M1007_g 0.00513266f $X=4.505 $Y=1.51 $X2=0 $Y2=0
cc_79 N_A_149_81#_M1009_g N_A_c_187_n 0.00139641f $X=3.335 $Y=2.965 $X2=0 $Y2=0
cc_80 N_A_149_81#_c_79_n N_A_c_187_n 0.0225651f $X=4.34 $Y=1.51 $X2=0 $Y2=0
cc_81 N_A_149_81#_c_82_n N_A_c_187_n 0.0232095f $X=4.505 $Y=2.34 $X2=0 $Y2=0
cc_82 N_A_149_81#_c_83_n N_A_c_187_n 0.00101103f $X=3.435 $Y=1.64 $X2=0 $Y2=0
cc_83 N_A_149_81#_M1004_g N_VPWR_c_196_n 0.07598f $X=0.995 $Y=2.965 $X2=0 $Y2=0
cc_84 N_A_149_81#_M1004_g N_VPWR_c_199_n 6.30116e-19 $X=0.995 $Y=2.965 $X2=2.4
+ $Y2=0.057
cc_85 N_A_149_81#_M1006_g N_VPWR_c_199_n 0.0726059f $X=1.775 $Y=2.965 $X2=2.4
+ $Y2=0.057
cc_86 N_A_149_81#_M1008_g N_VPWR_c_199_n 0.0679112f $X=2.555 $Y=2.965 $X2=2.4
+ $Y2=0.057
cc_87 N_A_149_81#_M1009_g N_VPWR_c_199_n 5.13552e-19 $X=3.335 $Y=2.965 $X2=2.4
+ $Y2=0.057
cc_88 N_A_149_81#_c_83_n N_VPWR_c_199_n 5.3984e-19 $X=3.435 $Y=1.64 $X2=2.4
+ $Y2=0.057
cc_89 N_A_149_81#_M1008_g N_VPWR_c_202_n 5.02847e-19 $X=2.555 $Y=2.965 $X2=0
+ $Y2=0
cc_90 N_A_149_81#_M1009_g N_VPWR_c_202_n 0.0694068f $X=3.335 $Y=2.965 $X2=0
+ $Y2=0
cc_91 N_A_149_81#_c_121_p N_VPWR_c_202_n 0.00386707f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_92 N_A_149_81#_c_82_n N_VPWR_c_202_n 0.0612867f $X=4.505 $Y=2.34 $X2=0 $Y2=0
cc_93 N_A_149_81#_c_106_p N_VPWR_c_202_n 0.00464317f $X=3.515 $Y=1.51 $X2=0
+ $Y2=0
cc_94 N_A_149_81#_M1001_d N_VPWR_c_205_n 0.00221032f $X=4.365 $Y=2.215 $X2=0
+ $Y2=0
cc_95 N_A_149_81#_M1004_g N_VPWR_c_205_n 0.0107323f $X=0.995 $Y=2.965 $X2=0
+ $Y2=0
cc_96 N_A_149_81#_M1006_g N_VPWR_c_205_n 0.00778801f $X=1.775 $Y=2.965 $X2=0
+ $Y2=0
cc_97 N_A_149_81#_M1008_g N_VPWR_c_205_n 0.0101061f $X=2.555 $Y=2.965 $X2=0
+ $Y2=0
cc_98 N_A_149_81#_M1009_g N_VPWR_c_205_n 0.0101228f $X=3.335 $Y=2.965 $X2=0
+ $Y2=0
cc_99 N_A_149_81#_c_82_n N_VPWR_c_205_n 0.0354327f $X=4.505 $Y=2.34 $X2=0 $Y2=0
cc_100 N_A_149_81#_M1000_g N_X_c_237_n 0.0124286f $X=0.995 $Y=0.91 $X2=0 $Y2=0
cc_101 N_A_149_81#_M1002_g N_X_c_237_n 9.97785e-19 $X=1.775 $Y=0.91 $X2=0 $Y2=0
cc_102 N_A_149_81#_M1000_g N_X_c_239_n 0.00194238f $X=0.995 $Y=0.91 $X2=0 $Y2=0
cc_103 N_A_149_81#_M1002_g N_X_c_239_n 8.86045e-19 $X=1.775 $Y=0.91 $X2=0 $Y2=0
cc_104 N_A_149_81#_c_83_n N_X_c_239_n 0.0149627f $X=3.435 $Y=1.64 $X2=0 $Y2=0
cc_105 N_A_149_81#_M1004_g N_X_c_257_n 0.0100021f $X=0.995 $Y=2.965 $X2=0 $Y2=0
cc_106 N_A_149_81#_c_121_p N_X_c_257_n 0.0135767f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_107 N_A_149_81#_c_83_n N_X_c_257_n 0.0272595f $X=3.435 $Y=1.64 $X2=0 $Y2=0
cc_108 N_A_149_81#_M1004_g N_X_c_245_n 0.0310842f $X=0.995 $Y=2.965 $X2=2.4
+ $Y2=0
cc_109 N_A_149_81#_M1006_g N_X_c_245_n 0.00480667f $X=1.775 $Y=2.965 $X2=2.4
+ $Y2=0
cc_110 N_A_149_81#_M1002_g N_X_c_240_n 0.0267003f $X=1.775 $Y=0.91 $X2=2.4
+ $Y2=0.058
cc_111 N_A_149_81#_M1003_g N_X_c_240_n 0.0261559f $X=2.555 $Y=0.91 $X2=2.4
+ $Y2=0.058
cc_112 N_A_149_81#_M1005_g N_X_c_240_n 0.00294046f $X=3.335 $Y=0.91 $X2=2.4
+ $Y2=0.058
cc_113 N_A_149_81#_c_121_p N_X_c_240_n 0.0985774f $X=3.43 $Y=1.64 $X2=2.4
+ $Y2=0.058
cc_114 N_A_149_81#_c_83_n N_X_c_240_n 0.00585093f $X=3.435 $Y=1.64 $X2=2.4
+ $Y2=0.058
cc_115 N_A_149_81#_M1006_g N_X_c_248_n 0.0220433f $X=1.775 $Y=2.965 $X2=0 $Y2=0
cc_116 N_A_149_81#_M1008_g N_X_c_248_n 0.0233066f $X=2.555 $Y=2.965 $X2=0 $Y2=0
cc_117 N_A_149_81#_M1009_g N_X_c_248_n 0.0100021f $X=3.335 $Y=2.965 $X2=0 $Y2=0
cc_118 N_A_149_81#_c_121_p N_X_c_248_n 0.102313f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_119 N_A_149_81#_c_83_n N_X_c_248_n 0.0305803f $X=3.435 $Y=1.64 $X2=0 $Y2=0
cc_120 N_A_149_81#_M1003_g N_X_c_241_n 0.0176338f $X=2.555 $Y=0.91 $X2=0 $Y2=0
cc_121 N_A_149_81#_M1005_g N_X_c_241_n 9.97785e-19 $X=3.335 $Y=0.91 $X2=0 $Y2=0
cc_122 N_A_149_81#_M1008_g N_X_c_249_n 0.0346038f $X=2.555 $Y=2.965 $X2=0 $Y2=0
cc_123 N_A_149_81#_M1009_g N_X_c_249_n 0.0359664f $X=3.335 $Y=2.965 $X2=0 $Y2=0
cc_124 N_A_149_81#_M1000_g N_X_c_243_n 0.00567795f $X=0.995 $Y=0.91 $X2=0 $Y2=0
cc_125 N_A_149_81#_c_83_n N_X_c_243_n 0.0016314f $X=3.435 $Y=1.64 $X2=0 $Y2=0
cc_126 N_A_149_81#_c_83_n N_X_c_244_n 0.0431855f $X=3.435 $Y=1.64 $X2=0 $Y2=0
cc_127 N_A_149_81#_M1000_g N_VGND_c_301_n 0.0534576f $X=0.995 $Y=0.91 $X2=0
+ $Y2=0
cc_128 N_A_149_81#_M1002_g N_VGND_c_301_n 5.45818e-19 $X=1.775 $Y=0.91 $X2=0
+ $Y2=0
cc_129 N_A_149_81#_M1000_g N_VGND_c_303_n 6.27378e-19 $X=0.995 $Y=0.91 $X2=0
+ $Y2=0
cc_130 N_A_149_81#_M1002_g N_VGND_c_303_n 0.0406305f $X=1.775 $Y=0.91 $X2=0
+ $Y2=0
cc_131 N_A_149_81#_M1003_g N_VGND_c_303_n 0.0365587f $X=2.555 $Y=0.91 $X2=0
+ $Y2=0
cc_132 N_A_149_81#_M1005_g N_VGND_c_303_n 4.60243e-19 $X=3.335 $Y=0.91 $X2=0
+ $Y2=0
cc_133 N_A_149_81#_M1003_g N_VGND_c_305_n 6.9169e-19 $X=2.555 $Y=0.91 $X2=0
+ $Y2=0
cc_134 N_A_149_81#_M1005_g N_VGND_c_305_n 0.0513588f $X=3.335 $Y=0.91 $X2=0
+ $Y2=0
cc_135 N_A_149_81#_c_121_p N_VGND_c_305_n 0.0102941f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_136 N_A_149_81#_c_79_n N_VGND_c_305_n 0.0380299f $X=4.34 $Y=1.51 $X2=0 $Y2=0
cc_137 N_A_149_81#_c_80_n N_VGND_c_305_n 0.0550348f $X=4.505 $Y=0.66 $X2=0 $Y2=0
cc_138 N_A_149_81#_c_106_p N_VGND_c_305_n 0.0121758f $X=3.515 $Y=1.51 $X2=0
+ $Y2=0
cc_139 N_A_149_81#_M1000_g N_VGND_c_307_n 0.0109133f $X=0.995 $Y=0.91 $X2=0
+ $Y2=0
cc_140 N_A_149_81#_M1002_g N_VGND_c_307_n 0.0041077f $X=1.775 $Y=0.91 $X2=0
+ $Y2=0
cc_141 N_A_149_81#_M1003_g N_VGND_c_307_n 0.00559592f $X=2.555 $Y=0.91 $X2=0
+ $Y2=0
cc_142 N_A_149_81#_M1005_g N_VGND_c_307_n 0.00774885f $X=3.335 $Y=0.91 $X2=0
+ $Y2=0
cc_143 N_A_149_81#_c_80_n N_VGND_c_307_n 0.0332558f $X=4.505 $Y=0.66 $X2=0 $Y2=0
cc_144 N_A_M1007_g N_VPWR_c_202_n 0.0724223f $X=4.115 $Y=0.91 $X2=0 $Y2=0
cc_145 N_A_c_187_n N_VPWR_c_202_n 0.0252067f $X=4.05 $Y=1.89 $X2=0 $Y2=0
cc_146 N_A_M1007_g N_VPWR_c_205_n 0.00854631f $X=4.115 $Y=0.91 $X2=0 $Y2=0
cc_147 N_A_M1007_g N_VGND_c_305_n 0.0469268f $X=4.115 $Y=0.91 $X2=0 $Y2=0
cc_148 N_A_M1007_g N_VGND_c_307_n 0.0115807f $X=4.115 $Y=0.91 $X2=0 $Y2=0
cc_149 N_VPWR_c_205_n N_X_M1004_s 0.00221032f $X=4.125 $Y=3.59 $X2=0 $Y2=0
cc_150 N_VPWR_c_196_n N_X_c_245_n 0.113499f $X=0.605 $Y=2.34 $X2=2.4 $Y2=4.013
cc_151 N_VPWR_c_199_n N_X_c_245_n 0.0630887f $X=2.165 $Y=2.34 $X2=2.4 $Y2=4.013
cc_152 N_VPWR_c_205_n N_X_c_245_n 0.0305382f $X=4.125 $Y=3.59 $X2=2.4 $Y2=4.013
cc_153 N_VPWR_c_199_n N_X_c_248_n 0.0658158f $X=2.165 $Y=2.34 $X2=0 $Y2=0
cc_154 N_VPWR_c_199_n N_X_c_249_n 0.109346f $X=2.165 $Y=2.34 $X2=0 $Y2=0
cc_155 N_VPWR_c_202_n N_X_c_249_n 0.105931f $X=3.725 $Y=2.385 $X2=0 $Y2=0
cc_156 N_VPWR_c_205_n N_X_c_249_n 0.0381262f $X=4.125 $Y=3.59 $X2=0 $Y2=0
cc_157 N_VPWR_c_196_n N_X_c_244_n 0.0413608f $X=0.605 $Y=2.34 $X2=0 $Y2=0
cc_158 N_X_c_240_n N_VGND_M1002_d 0.00177996f $X=2.78 $Y=1.29 $X2=0 $Y2=0
cc_159 N_X_c_237_n N_VGND_c_301_n 0.0510899f $X=1.385 $Y=0.66 $X2=0 $Y2=0
cc_160 N_X_c_243_n N_VGND_c_301_n 0.00965422f $X=1.345 $Y=1.29 $X2=0 $Y2=0
cc_161 N_X_c_244_n N_VGND_c_301_n 0.0621648f $X=1.22 $Y=1.665 $X2=0 $Y2=0
cc_162 N_X_c_237_n N_VGND_c_303_n 0.0228725f $X=1.385 $Y=0.66 $X2=0 $Y2=0
cc_163 N_X_c_240_n N_VGND_c_303_n 0.0597017f $X=2.78 $Y=1.29 $X2=0 $Y2=0
cc_164 N_X_c_241_n N_VGND_c_303_n 0.0377331f $X=2.945 $Y=0.66 $X2=0 $Y2=0
cc_165 N_X_c_241_n N_VGND_c_305_n 0.0300809f $X=2.945 $Y=0.66 $X2=0 $Y2=0
cc_166 N_X_M1000_s N_VGND_c_307_n 7.45741e-19 $X=1.245 $Y=0.535 $X2=0 $Y2=0
cc_167 N_X_M1003_s N_VGND_c_307_n 0.00221032f $X=2.805 $Y=0.535 $X2=0 $Y2=0
cc_168 N_X_c_237_n N_VGND_c_307_n 0.0243085f $X=1.385 $Y=0.66 $X2=0 $Y2=0
cc_169 N_X_c_240_n N_VGND_c_307_n 0.0130199f $X=2.78 $Y=1.29 $X2=0 $Y2=0
cc_170 N_X_c_241_n N_VGND_c_307_n 0.0243085f $X=2.945 $Y=0.66 $X2=0 $Y2=0
