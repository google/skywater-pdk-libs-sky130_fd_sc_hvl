* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
X0 VPWR a_30_131# a_340_593# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X1 a_2553_203# a_1787_137# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 VPWR a_2553_203# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X3 VGND a_798_107# a_1645_137# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_958_107# a_1000_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 a_1989_203# a_2031_177# a_2131_203# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X6 a_1268_251# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X7 a_982_529# a_1000_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X8 VPWR a_798_107# a_1000_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X9 a_1653_515# a_30_131# a_1787_137# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X10 VGND a_1787_137# a_2031_177# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X11 a_1787_137# a_340_593# a_1989_515# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X12 a_642_107# a_340_593# a_798_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X13 a_2553_203# a_1787_137# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X14 a_798_107# a_30_131# a_982_529# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X15 VPWR SET_B a_1787_137# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X16 a_642_107# a_30_131# a_798_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 a_1645_137# a_340_593# a_1787_137# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 VGND a_2553_203# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X19 a_2031_177# a_1787_137# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X20 a_1000_81# a_798_107# a_1268_251# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X21 a_30_131# CLK VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X22 VGND D a_642_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X23 a_2131_203# SET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X24 a_1989_515# a_2031_177# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X25 a_1000_81# SET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X26 VGND a_30_131# a_340_593# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X27 VPWR D a_642_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X28 VPWR a_798_107# a_1653_515# VPB sky130_fd_pr__pfet_g5v0d10v5 w=1e+06u l=500000u
X29 a_30_131# CLK VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X30 a_798_107# a_340_593# a_958_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X31 a_1787_137# a_30_131# a_1989_203# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends
