* NGSPICE file created from sky130_fd_sc_hvl__sdlxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__sdlxtp_1 D GATE SCD SCE VGND VNB VPB VPWR Q
M1000 a_1724_593# a_1214_107# a_1480_107# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=2.5995e+11p ps=2.29e+06u
M1001 VPWR a_1678_81# a_1724_593# VPB phv w=420000u l=500000u
+  ad=1.2621e+12p pd=1.158e+07u as=0p ps=0u
M1002 a_1480_107# a_1214_107# a_489_107# VNB nhv w=420000u l=500000u
+  ad=1.176e+11p pd=1.4e+06u as=2.289e+11p ps=2.77e+06u
M1003 a_660_587# a_30_587# a_489_107# VPB phv w=750000u l=500000u
+  ad=1.575e+11p pd=1.92e+06u as=4.2375e+11p ps=4.13e+06u
M1004 VGND SCE a_30_587# VNB nhv w=420000u l=500000u
+  ad=7.1325e+11p pd=7.84e+06u as=1.197e+11p ps=1.41e+06u
M1005 a_1214_107# a_944_107# VGND VNB nhv w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1006 a_944_107# GATE VGND VNB nhv w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 a_1480_107# a_944_107# a_489_107# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_645_107# SCE a_489_107# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1009 VGND SCD a_645_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_362_587# SCE VPWR VPB phv w=750000u l=500000u
+  ad=1.575e+11p pd=1.92e+06u as=0p ps=0u
M1011 VPWR a_1480_107# a_1678_81# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1012 VPWR SCD a_660_587# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_1480_107# a_1678_81# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1014 a_1214_107# a_944_107# VPWR VPB phv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
M1015 a_347_107# D VGND VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1016 a_489_107# a_30_587# a_347_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_489_107# D a_362_587# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR SCE a_30_587# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1019 a_1636_107# a_944_107# a_1480_107# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1020 Q a_1480_107# VGND VNB nhv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
M1021 Q a_1480_107# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=0p ps=0u
M1022 VGND a_1678_81# a_1636_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_944_107# GATE VPWR VPB phv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
.ends

