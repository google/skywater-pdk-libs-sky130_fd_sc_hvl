* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1569_126# a_1290_126# VGND VNB nhv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=1.1909e+12p ps=1.226e+07u
M1001 a_496_655# D a_339_655# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=3.738e+11p ps=4.3e+06u
M1002 a_1290_126# CLK VPWR VPB phv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=2.188e+12p ps=2.015e+07u
M1003 a_2014_537# a_1816_659# VPWR VPB phv w=1e+06u l=500000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1004 a_1999_126# a_1569_126# a_1816_659# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1005 a_2141_126# a_2014_537# a_1999_126# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1006 a_339_655# a_222_131# a_794_655# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1007 VGND RESET_B a_361_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=3.0115e+11p ps=3.2e+06u
M1008 VGND RESET_B a_2141_126# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_2624_107# a_3613_443# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1010 Q a_3613_443# VGND VNB nhv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
M1011 a_2871_543# a_1569_126# a_2624_107# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=3.312e+11p ps=2.79e+06u
M1012 VPWR RESET_B a_339_655# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1816_659# RESET_B VPWR VPB phv w=420000u l=500000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1014 a_3098_107# RESET_B VGND VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1015 a_2841_81# a_2624_107# a_3098_107# VNB nhv w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1016 VPWR SCE a_496_655# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1816_659# a_1569_126# a_339_655# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_222_131# SCE VPWR VPB phv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1019 a_1569_126# a_1290_126# VPWR VPB phv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
M1020 a_2799_107# a_1290_126# a_2624_107# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=2.4495e+11p ps=2.25e+06u
M1021 VPWR a_2624_107# a_2841_81# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1022 Q a_3613_443# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=0p ps=0u
M1023 Q_N a_2624_107# VGND VNB nhv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
M1024 a_2624_107# a_1290_126# a_2014_537# VPB phv w=1e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_2841_81# a_2871_543# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1290_126# CLK VGND VNB nhv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1027 a_1816_659# a_1290_126# a_339_655# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=2.373e+11p ps=2.81e+06u
M1028 a_2624_107# a_1569_126# a_2014_537# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=2.1e+11p ps=2.06e+06u
M1029 a_222_131# SCE VGND VNB nhv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1030 VGND a_2841_81# a_2799_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_816_107# SCE a_339_655# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1032 Q_N a_2624_107# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=3.975e+11p pd=3.53e+06u as=0p ps=0u
M1033 a_794_655# SCD VPWR VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2841_81# RESET_B VPWR VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_361_107# SCD a_816_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR a_2624_107# a_3613_443# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u
M1037 a_1972_659# a_1290_126# a_1816_659# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1038 VPWR a_2014_537# a_1972_659# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2014_537# a_1816_659# VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_518_107# D a_361_107# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1041 a_339_655# a_222_131# a_518_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
