# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
SITE unithvdbl
    SYMMETRY y  ;
    CLASS CORE  ;
    SIZE  0.480 BY 8.140 ;
END unithvdbl
MACRO sky130_fd_sc_hvl__sdfstp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  18.72000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.845000 2.275000 2.355000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.478750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.260000 0.495000 18.610000 3.395000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.420000 1.175000 3.750000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.495000 2.890000 1.665000 ;
        RECT 0.565000 1.665000 0.895000 2.165000 ;
        RECT 2.525000 1.095000 2.890000 1.495000 ;
        RECT 2.525000 1.665000 2.890000 1.780000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.535000 1.175000 11.635000 1.345000 ;
        RECT 11.465000 0.265000 14.215000 0.435000 ;
        RECT 11.465000 0.435000 11.635000 1.175000 ;
        RECT 14.045000 0.435000 14.215000 0.810000 ;
        RECT 14.045000 0.810000 14.520000 1.760000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.175000 4.525000 2.150000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.620000 0.365000 1.570000 0.915000 ;
    END
    PORT
      LAYER li1 ;
        RECT 10.335000 0.365000 11.285000 0.995000 ;
    END
    PORT
      LAYER li1 ;
        RECT 14.700000 0.365000 15.590000 1.325000 ;
    END
    PORT
      LAYER li1 ;
        RECT 17.095000 0.365000 18.045000 1.325000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.420000 0.365000 4.370000 0.995000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.200000 0.365000 5.450000 1.055000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.200000 0.365000 9.150000 0.925000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 18.720000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 18.720000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 18.720000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 18.720000 4.155000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 18.720000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.620000 2.885000 1.570000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 10.835000 3.285000 11.785000 3.755000 ;
    END
    PORT
      LAYER li1 ;
        RECT 13.265000 2.675000 14.215000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 15.815000 3.045000 16.405000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 17.135000 2.355000 18.080000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.420000 2.805000 4.315000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.545000 2.625000 5.725000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.495000 2.925000 9.445000 3.705000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 18.720000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.110000 0.515000  0.440000 1.095000 ;
      RECT  0.110000 1.095000  2.255000 1.315000 ;
      RECT  0.110000 1.315000  0.280000 2.535000 ;
      RECT  0.110000 2.535000  2.890000 2.705000 ;
      RECT  0.110000 2.705000  0.440000 3.285000 ;
      RECT  2.380000 0.495000  2.710000 0.745000 ;
      RECT  2.380000 0.745000  3.240000 0.915000 ;
      RECT  2.380000 2.885000  3.240000 3.055000 ;
      RECT  2.380000 3.055000  2.710000 3.305000 ;
      RECT  2.635000 2.015000  2.890000 2.535000 ;
      RECT  3.070000 0.915000  3.240000 2.455000 ;
      RECT  3.070000 2.455000  4.665000 2.625000 ;
      RECT  3.070000 2.625000  3.240000 2.885000 ;
      RECT  4.495000 2.625000  4.665000 3.635000 ;
      RECT  4.495000 3.635000  5.365000 3.805000 ;
      RECT  4.650000 0.515000  5.015000 0.975000 ;
      RECT  4.845000 0.975000  5.015000 1.735000 ;
      RECT  4.845000 1.735000  5.835000 1.905000 ;
      RECT  4.845000 1.905000  5.015000 3.455000 ;
      RECT  5.195000 2.275000  6.075000 2.445000 ;
      RECT  5.195000 2.445000  5.365000 3.635000 ;
      RECT  5.505000 1.235000  5.835000 1.735000 ;
      RECT  5.630000 0.265000  7.230000 0.435000 ;
      RECT  5.630000 0.435000  5.800000 1.235000 ;
      RECT  5.905000 2.445000  6.075000 3.635000 ;
      RECT  5.905000 3.635000  7.095000 3.805000 ;
      RECT  5.980000 0.675000  6.310000 1.055000 ;
      RECT  6.140000 1.055000  6.310000 1.425000 ;
      RECT  6.140000 1.425000  6.530000 2.095000 ;
      RECT  6.255000 2.095000  6.530000 3.455000 ;
      RECT  6.550000 0.615000  6.880000 1.025000 ;
      RECT  6.710000 1.025000  6.880000 2.675000 ;
      RECT  6.710000 2.675000  7.095000 3.635000 ;
      RECT  7.060000 0.435000  7.230000 1.605000 ;
      RECT  7.060000 1.605000  7.445000 1.775000 ;
      RECT  7.275000 1.775000  7.445000 3.355000 ;
      RECT  7.275000 3.355000  8.305000 3.525000 ;
      RECT  7.410000 0.525000  7.795000 1.025000 ;
      RECT  7.625000 1.025000  7.795000 1.355000 ;
      RECT  7.625000 1.355000  8.655000 1.525000 ;
      RECT  7.625000 1.525000  7.795000 2.675000 ;
      RECT  7.625000 2.675000  7.955000 3.175000 ;
      RECT  7.975000 1.705000  8.305000 1.875000 ;
      RECT  7.975000 1.875000 12.220000 2.045000 ;
      RECT  8.135000 2.225000  8.410000 2.575000 ;
      RECT  8.135000 2.575000  9.795000 2.745000 ;
      RECT  8.135000 2.745000  8.305000 3.355000 ;
      RECT  8.485000 1.525000 11.525000 1.695000 ;
      RECT  8.790000 2.225000 10.305000 2.395000 ;
      RECT  8.835000 1.105000  9.700000 1.275000 ;
      RECT  8.835000 1.275000  9.165000 1.345000 ;
      RECT  9.370000 0.515000  9.700000 1.105000 ;
      RECT  9.520000 1.455000  9.850000 1.525000 ;
      RECT  9.625000 2.745000  9.795000 3.105000 ;
      RECT  9.625000 3.105000 10.655000 3.275000 ;
      RECT  9.975000 2.395000 10.305000 2.925000 ;
      RECT 10.485000 2.935000 12.180000 3.105000 ;
      RECT 11.905000 2.225000 12.570000 2.395000 ;
      RECT 11.905000 2.395000 12.180000 2.935000 ;
      RECT 11.970000 1.685000 12.220000 1.875000 ;
      RECT 12.095000 0.615000 13.350000 0.785000 ;
      RECT 12.095000 0.785000 12.265000 1.335000 ;
      RECT 12.095000 1.335000 12.570000 1.505000 ;
      RECT 12.360000 2.675000 12.920000 2.845000 ;
      RECT 12.360000 2.845000 12.690000 3.755000 ;
      RECT 12.400000 1.505000 12.570000 2.225000 ;
      RECT 12.445000 0.965000 12.920000 1.155000 ;
      RECT 12.750000 1.155000 12.920000 1.940000 ;
      RECT 12.750000 1.940000 15.585000 2.110000 ;
      RECT 12.750000 2.110000 12.920000 2.675000 ;
      RECT 13.100000 0.785000 13.350000 1.745000 ;
      RECT 13.710000 2.290000 14.565000 2.495000 ;
      RECT 14.395000 2.495000 14.565000 3.335000 ;
      RECT 14.395000 3.335000 15.625000 3.505000 ;
      RECT 14.745000 2.110000 15.585000 2.175000 ;
      RECT 14.745000 2.175000 15.075000 3.155000 ;
      RECT 15.255000 1.505000 15.585000 1.940000 ;
      RECT 15.295000 2.695000 16.020000 2.865000 ;
      RECT 15.295000 2.865000 15.625000 3.335000 ;
      RECT 15.770000 0.825000 16.020000 2.695000 ;
      RECT 16.585000 0.825000 16.915000 1.505000 ;
      RECT 16.585000 1.505000 18.080000 1.675000 ;
      RECT 16.585000 1.675000 16.915000 2.355000 ;
      RECT 16.585000 2.355000 16.955000 3.145000 ;
      RECT 17.750000 1.675000 18.080000 2.175000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.650000  0.395000  0.820000 0.565000 ;
      RECT  0.650000  3.505000  0.820000 3.675000 ;
      RECT  1.010000  0.395000  1.180000 0.565000 ;
      RECT  1.010000  3.505000  1.180000 3.675000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.370000  0.395000  1.540000 0.565000 ;
      RECT  1.370000  3.505000  1.540000 3.675000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.420000  3.505000  3.590000 3.675000 ;
      RECT  3.450000  0.395000  3.620000 0.565000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.780000  3.505000  3.950000 3.675000 ;
      RECT  3.810000  0.395000  3.980000 0.565000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.140000  3.505000  4.310000 3.675000 ;
      RECT  4.170000  0.395000  4.340000 0.565000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.230000  0.395000  5.400000 0.565000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.550000  3.505000  5.720000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.230000  0.395000  8.400000 0.565000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.525000  3.505000  8.695000 3.675000 ;
      RECT  8.590000  0.395000  8.760000 0.565000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.885000  3.505000  9.055000 3.675000 ;
      RECT  8.950000  0.395000  9.120000 0.565000 ;
      RECT  9.245000  3.505000  9.415000 3.675000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.365000  0.395000 10.535000 0.565000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.725000  0.395000 10.895000 0.565000 ;
      RECT 10.865000  3.505000 11.035000 3.675000 ;
      RECT 11.085000  0.395000 11.255000 0.565000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.225000  3.505000 11.395000 3.675000 ;
      RECT 11.585000  3.505000 11.755000 3.675000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.295000  3.505000 13.465000 3.675000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.655000  3.505000 13.825000 3.675000 ;
      RECT 14.015000  3.505000 14.185000 3.675000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.700000  0.395000 14.870000 0.565000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.060000  0.395000 15.230000 0.565000 ;
      RECT 15.420000  0.395000 15.590000 0.565000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.845000  3.505000 16.015000 3.675000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.205000  3.505000 16.375000 3.675000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 17.125000  0.395000 17.295000 0.565000 ;
      RECT 17.160000  3.505000 17.330000 3.675000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
      RECT 17.485000  0.395000 17.655000 0.565000 ;
      RECT 17.520000  3.505000 17.690000 3.675000 ;
      RECT 17.845000  0.395000 18.015000 0.565000 ;
      RECT 17.880000  3.505000 18.050000 3.675000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.985000 18.085000 4.155000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.985000 18.565000 4.155000 ;
  END
END sky130_fd_sc_hvl__sdfstp_1
END LIBRARY
