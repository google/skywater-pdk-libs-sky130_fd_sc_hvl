* File: sky130_fd_sc_hvl__sdfrtp_1.pex.spice
* Created: Wed Sep  2 09:10:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%VNB 5 7 11
c130 5 0 5.08179e-19 $X=-0.33 $Y=-0.265
r131 7 11 0.000371094 $w=1.92e-05 $l=5.7e-08 $layer=MET1_cond $X=9.6 $Y=0.057
+ $X2=9.6 $Y2=0
r132 5 11 0.465 $w=1.7e-07 $l=3.4e-06 $layer=mcon $count=20 $X=18.96 $Y=0
+ $X2=18.96 $Y2=0
r133 5 11 0.465 $w=1.7e-07 $l=3.4e-06 $layer=mcon $count=20 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%VPB 4 6 14
r208 10 14 0.465 $w=1.7e-07 $l=3.4e-06 $layer=mcon $count=20 $X=18.96 $Y=4.07
+ $X2=18.96 $Y2=4.07
r209 9 14 1221.3 $w=1.68e-07 $l=1.872e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=18.96 $Y2=4.07
r210 9 10 0.465 $w=1.7e-07 $l=3.4e-06 $layer=mcon $count=20 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r211 6 10 0.000371094 $w=1.92e-05 $l=5.7e-08 $layer=MET1_cond $X=9.6 $Y=4.013
+ $X2=9.6 $Y2=4.07
r212 4 14 9.1 $w=1.7e-07 $l=1.90025e-05 $layer=licon1_NTAP_notbjt $count=20 $X=0
+ $Y=3.985 $X2=18.96 $Y2=4.07
r213 4 9 9.1 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=20 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%A_116_451# 1 2 7 9 11 13 17 20 21 23 24 25
+ 26 29 30 31 32 35 36 37 40 44 46 47
c161 47 0 1.50894e-19 $X=2.645 $Y=1.18
r162 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=1.57 $X2=2.645 $Y2=1.57
r163 49 51 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.645 $Y=1.26
+ $X2=2.645 $Y2=1.57
r164 47 49 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.645 $Y=1.18
+ $X2=2.645 $Y2=1.26
r165 42 44 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.41 $Y=1.175
+ $X2=5.41 $Y2=0.84
r166 38 40 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.32 $Y=2.875
+ $X2=5.32 $Y2=3.37
r167 36 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.155 $Y=2.79
+ $X2=5.32 $Y2=2.875
r168 36 37 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=5.155 $Y=2.79
+ $X2=3.555 $Y2=2.79
r169 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.47 $Y=2.705
+ $X2=3.555 $Y2=2.79
r170 34 35 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.47 $Y=2.48
+ $X2=3.47 $Y2=2.705
r171 33 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.81 $Y=1.26
+ $X2=2.645 $Y2=1.26
r172 32 42 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.285 $Y=1.26
+ $X2=5.41 $Y2=1.175
r173 32 33 161.471 $w=1.68e-07 $l=2.475e-06 $layer=LI1_cond $X=5.285 $Y=1.26
+ $X2=2.81 $Y2=1.26
r174 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.385 $Y=2.395
+ $X2=3.47 $Y2=2.48
r175 30 31 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.385 $Y=2.395
+ $X2=2.73 $Y2=2.395
r176 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.645 $Y=2.48
+ $X2=2.73 $Y2=2.395
r177 28 29 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.645 $Y=2.48
+ $X2=2.645 $Y2=2.755
r178 27 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.815 $Y=2.84
+ $X2=1.73 $Y2=2.84
r179 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.56 $Y=2.84
+ $X2=2.645 $Y2=2.755
r180 26 27 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.56 $Y=2.84
+ $X2=1.815 $Y2=2.84
r181 24 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=1.18
+ $X2=2.645 $Y2=1.18
r182 24 25 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.48 $Y=1.18
+ $X2=1.815 $Y2=1.18
r183 23 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=2.755
+ $X2=1.73 $Y2=2.84
r184 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.73 $Y=1.265
+ $X2=1.815 $Y2=1.18
r185 22 23 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=1.73 $Y=1.265
+ $X2=1.73 $Y2=2.755
r186 20 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=2.84
+ $X2=1.73 $Y2=2.84
r187 20 21 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.645 $Y=2.84
+ $X2=1.06 $Y2=2.84
r188 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.895
+ $Y=2.42 $X2=0.895 $Y2=2.42
r189 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.895 $Y=2.755
+ $X2=1.06 $Y2=2.84
r190 15 17 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.895 $Y=2.755
+ $X2=0.895 $Y2=2.42
r191 11 52 25.3258 $w=5e-07 $l=2.55e-07 $layer=POLY_cond $X=2.71 $Y=1.315
+ $X2=2.71 $Y2=1.57
r192 11 13 50.8278 $w=5e-07 $l=4.75e-07 $layer=POLY_cond $X=2.71 $Y=1.315
+ $X2=2.71 $Y2=0.84
r193 7 18 65.8134 $w=5.09e-07 $l=7.0246e-07 $layer=POLY_cond $X=0.86 $Y=3.115
+ $X2=0.845 $Y2=2.42
r194 7 9 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.86 $Y=3.115 $X2=0.86
+ $Y2=3.455
r195 2 40 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=5.18
+ $Y=3.245 $X2=5.32 $Y2=3.37
r196 1 44 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.23
+ $Y=0.63 $X2=5.37 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%SCD 1 3 5 8 10 11 14 15 24
c51 5 0 1.36627e-19 $X=1.22 $Y=1.985
r52 23 24 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.345 $X2=0.95 $Y2=1.345
r53 19 23 93.3789 $w=4.05e-07 $l=6.8e-07 $layer=POLY_cond $X=0.27 $Y=1.362
+ $X2=0.95 $Y2=1.362
r54 15 24 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.72 $Y=1.345
+ $X2=0.95 $Y2=1.345
r55 14 15 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.345
+ $X2=0.72 $Y2=1.345
r56 14 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.345 $X2=0.27 $Y2=1.345
r57 10 23 2.74644 $w=4.05e-07 $l=2e-08 $layer=POLY_cond $X=0.97 $Y=1.362
+ $X2=0.95 $Y2=1.362
r58 10 11 8.34116 $w=4.05e-07 $l=2.5e-07 $layer=POLY_cond $X=0.97 $Y=1.362
+ $X2=1.22 $Y2=1.362
r59 6 8 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=1.57 $Y=2.405 $X2=1.57
+ $Y2=3.455
r60 5 6 57.774 $w=2.92e-07 $l=4.42719e-07 $layer=POLY_cond $X=1.22 $Y=1.985
+ $X2=1.57 $Y2=2.195
r61 4 11 17.0691 $w=5e-07 $l=2.03e-07 $layer=POLY_cond $X=1.22 $Y=1.565 $X2=1.22
+ $Y2=1.362
r62 4 5 44.9425 $w=5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.22 $Y=1.565 $X2=1.22
+ $Y2=1.985
r63 1 11 17.0691 $w=5e-07 $l=2.02e-07 $layer=POLY_cond $X=1.22 $Y=1.16 $X2=1.22
+ $Y2=1.362
r64 1 3 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.22 $Y=1.16 $X2=1.22
+ $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%SCE 3 5 7 11 15 18 19 23 26 28 29 30 31 32
+ 33 43 52
c129 43 0 1.34856e-19 $X=4.98 $Y=0.84
c130 33 0 5.7967e-21 $X=5.52 $Y=1.665
c131 28 0 1.36627e-19 $X=2.187 $Y=1.92
c132 23 0 1.21896e-19 $X=2.215 $Y=2.15
c133 19 0 9.7103e-20 $X=2.08 $Y=1.61
c134 3 0 1.50894e-19 $X=1.93 $Y=0.84
r135 53 65 14.8749 $w=1.68e-07 $l=2.28e-07 $layer=LI1_cond $X=3.09 $Y=1.692
+ $X2=3.09 $Y2=1.92
r136 47 52 5.19621 $w=7.53e-07 $l=3.28e-07 $layer=LI1_cond $X=5.257 $Y=2.02
+ $X2=5.257 $Y2=1.692
r137 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.045
+ $Y=2.02 $X2=5.045 $Y2=2.02
r138 43 46 126.267 $w=5e-07 $l=1.18e-06 $layer=POLY_cond $X=4.98 $Y=0.84
+ $X2=4.98 $Y2=2.02
r139 33 52 0.427737 $w=7.53e-07 $l=2.7e-08 $layer=LI1_cond $X=5.257 $Y=1.665
+ $X2=5.257 $Y2=1.692
r140 32 52 12.9397 $w=2.83e-07 $l=3.2e-07 $layer=LI1_cond $X=4.56 $Y=1.692
+ $X2=4.88 $Y2=1.692
r141 31 32 19.4096 $w=2.83e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.692
+ $X2=4.56 $Y2=1.692
r142 30 31 19.4096 $w=2.83e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.692
+ $X2=4.08 $Y2=1.692
r143 29 53 1.7615 $w=1.68e-07 $l=2.7e-08 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=1.692
r144 29 30 16.579 $w=2.83e-07 $l=4.1e-07 $layer=LI1_cond $X=3.19 $Y=1.692
+ $X2=3.6 $Y2=1.692
r145 29 53 0.606549 $w=2.83e-07 $l=1.5e-08 $layer=LI1_cond $X=3.19 $Y=1.692
+ $X2=3.175 $Y2=1.692
r146 27 28 3.66292 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.38 $Y=1.92
+ $X2=2.187 $Y2=1.92
r147 26 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.005 $Y=1.92
+ $X2=3.09 $Y2=1.92
r148 26 27 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.005 $Y=1.92
+ $X2=2.38 $Y2=1.92
r149 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.215
+ $Y=2.15 $X2=2.215 $Y2=2.15
r150 21 28 2.99104 $w=3.17e-07 $l=8.5e-08 $layer=LI1_cond $X=2.187 $Y=2.005
+ $X2=2.187 $Y2=1.92
r151 21 23 4.34037 $w=3.83e-07 $l=1.45e-07 $layer=LI1_cond $X=2.187 $Y=2.005
+ $X2=2.187 $Y2=2.15
r152 19 49 32.3893 $w=5.7e-07 $l=3.35e-07 $layer=POLY_cond $X=1.965 $Y=1.61
+ $X2=1.965 $Y2=1.275
r153 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.61 $X2=2.08 $Y2=1.61
r154 16 28 2.99104 $w=3.17e-07 $l=1.13666e-07 $layer=LI1_cond $X=2.12 $Y=1.835
+ $X2=2.187 $Y2=1.92
r155 16 18 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=2.12 $Y=1.835
+ $X2=2.12 $Y2=1.61
r156 14 46 2.67515 $w=5e-07 $l=2.5e-08 $layer=POLY_cond $X=4.98 $Y=2.045
+ $X2=4.98 $Y2=2.02
r157 14 15 48.639 $w=5.5e-07 $l=5e-07 $layer=POLY_cond $X=4.955 $Y=2.045
+ $X2=4.955 $Y2=2.545
r158 11 15 97.3754 $w=5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.93 $Y=3.455
+ $X2=4.93 $Y2=2.545
r159 5 24 48.034 $w=5.29e-07 $l=5.47037e-07 $layer=POLY_cond $X=2.37 $Y=2.675
+ $X2=2.325 $Y2=2.15
r160 5 7 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.37 $Y=2.675 $X2=2.37
+ $Y2=3.455
r161 3 49 46.5476 $w=5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.84 $X2=1.93
+ $Y2=1.275
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%D 1 3 10 11 15 18
c57 15 0 4.66067e-19 $X=3.06 $Y=2.825
c58 10 0 1.36153e-20 $X=3.12 $Y=2.775
r59 15 18 67.4137 $w=5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.08 $Y=2.825 $X2=3.08
+ $Y2=3.455
r60 10 11 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=3.057 $Y=2.775
+ $X2=3.057 $Y2=3.145
r61 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.06
+ $Y=2.825 $X2=3.06 $Y2=2.825
r62 6 15 55.6431 $w=5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.08 $Y=2.305 $X2=3.08
+ $Y2=2.825
r63 1 6 126.062 $w=1.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.42 $Y=2.24 $X2=3.08
+ $Y2=2.24
r64 1 3 142.853 $w=5e-07 $l=1.335e-06 $layer=POLY_cond $X=3.42 $Y=2.175 $X2=3.42
+ $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%A_1212_471# 1 2 7 9 13 14 15 16 17 18 20
+ 23 27 28 29 30 33 34 35 38 41 42 46 50 51 55 56 58 60 64 67 69 73 76 83
c239 58 0 1.33662e-19 $X=7.15 $Y=1.26
c240 30 0 7.88029e-20 $X=9.305 $Y=1.26
r241 65 67 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=11.395 $Y=2.37
+ $X2=11.705 $Y2=2.37
r242 60 62 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=9.47 $Y=1.115
+ $X2=9.47 $Y2=1.26
r243 56 83 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=12.62 $Y=2.39
+ $X2=12.62 $Y2=2.925
r244 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.645
+ $Y=2.39 $X2=12.645 $Y2=2.39
r245 53 55 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=12.645 $Y=3.135
+ $X2=12.645 $Y2=2.39
r246 52 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.79 $Y=3.22
+ $X2=11.705 $Y2=3.22
r247 51 53 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.48 $Y=3.22
+ $X2=12.645 $Y2=3.135
r248 51 52 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.48 $Y=3.22
+ $X2=11.79 $Y2=3.22
r249 50 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.705 $Y=3.135
+ $X2=11.705 $Y2=3.22
r250 49 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.705 $Y=2.455
+ $X2=11.705 $Y2=2.37
r251 49 50 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=11.705 $Y=2.455
+ $X2=11.705 $Y2=3.135
r252 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.395
+ $Y=1.63 $X2=11.395 $Y2=1.63
r253 44 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.395 $Y=2.285
+ $X2=11.395 $Y2=2.37
r254 44 46 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=11.395 $Y=2.285
+ $X2=11.395 $Y2=1.63
r255 43 64 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.785 $Y=3.22
+ $X2=9.62 $Y2=3.22
r256 42 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.62 $Y=3.22
+ $X2=11.705 $Y2=3.22
r257 42 43 119.717 $w=1.68e-07 $l=1.835e-06 $layer=LI1_cond $X=11.62 $Y=3.22
+ $X2=9.785 $Y2=3.22
r258 40 64 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.62 $Y=3.305
+ $X2=9.62 $Y2=3.22
r259 40 41 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=9.62 $Y=3.305
+ $X2=9.62 $Y2=3.635
r260 36 64 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.62 $Y=3.135
+ $X2=9.62 $Y2=3.22
r261 36 38 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.62 $Y=3.135
+ $X2=9.62 $Y2=2.86
r262 34 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.455 $Y=3.72
+ $X2=9.62 $Y2=3.635
r263 34 35 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=9.455 $Y=3.72
+ $X2=8.705 $Y2=3.72
r264 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.62 $Y=3.635
+ $X2=8.705 $Y2=3.72
r265 32 33 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=8.62 $Y=3.235
+ $X2=8.62 $Y2=3.635
r266 31 58 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.255 $Y=1.26
+ $X2=7.15 $Y2=1.26
r267 30 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.305 $Y=1.26
+ $X2=9.47 $Y2=1.26
r268 30 31 133.743 $w=1.68e-07 $l=2.05e-06 $layer=LI1_cond $X=9.305 $Y=1.26
+ $X2=7.255 $Y2=1.26
r269 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.535 $Y=3.15
+ $X2=8.62 $Y2=3.235
r270 28 29 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=8.535 $Y=3.15
+ $X2=7.215 $Y2=3.15
r271 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.13 $Y=3.235
+ $X2=7.215 $Y2=3.15
r272 26 27 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.13 $Y=3.235
+ $X2=7.13 $Y2=3.635
r273 24 76 78.1143 $w=5e-07 $l=7.3e-07 $layer=POLY_cond $X=7.09 $Y=1.57 $X2=7.09
+ $Y2=0.84
r274 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.15
+ $Y=1.57 $X2=7.15 $Y2=1.57
r275 21 58 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.15 $Y=1.345
+ $X2=7.15 $Y2=1.26
r276 21 23 11.8831 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=7.15 $Y=1.345
+ $X2=7.15 $Y2=1.57
r277 20 58 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.15 $Y=1.175
+ $X2=7.15 $Y2=1.26
r278 19 20 39.0823 $w=2.08e-07 $l=7.4e-07 $layer=LI1_cond $X=7.15 $Y=0.435
+ $X2=7.15 $Y2=1.175
r279 17 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.045 $Y=3.72
+ $X2=7.13 $Y2=3.635
r280 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.045 $Y=3.72
+ $X2=6.355 $Y2=3.72
r281 15 19 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.045 $Y=0.35
+ $X2=7.15 $Y2=0.435
r282 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.045 $Y=0.35
+ $X2=6.355 $Y2=0.35
r283 14 73 93.6302 $w=5e-07 $l=8.75e-07 $layer=POLY_cond $X=6.31 $Y=2.54
+ $X2=6.31 $Y2=3.415
r284 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.27
+ $Y=2.54 $X2=6.27 $Y2=2.54
r285 11 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.27 $Y=3.635
+ $X2=6.355 $Y2=3.72
r286 11 13 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=6.27 $Y=3.635
+ $X2=6.27 $Y2=2.54
r287 10 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.27 $Y=0.435
+ $X2=6.355 $Y2=0.35
r288 10 13 137.332 $w=1.68e-07 $l=2.105e-06 $layer=LI1_cond $X=6.27 $Y=0.435
+ $X2=6.27 $Y2=2.54
r289 7 47 17.5532 $w=5.08e-07 $l=2.01742e-07 $layer=POLY_cond $X=11.55 $Y=1.445
+ $X2=11.515 $Y2=1.63
r290 7 9 47.718 $w=5e-07 $l=4.95e-07 $layer=POLY_cond $X=11.55 $Y=1.445
+ $X2=11.55 $Y2=0.95
r291 2 38 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=9.495
+ $Y=2.715 $X2=9.62 $Y2=2.86
r292 1 60 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.345
+ $Y=0.905 $X2=9.47 $Y2=1.115
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%A_1212_100# 1 2 9 11 12 13 15 17 19 20 22
+ 24 26 28 31 35 39 40 41 46 47 48 49 55 56 59 60 61 65 66 67 70 72 73 75 78 83
+ 84
c269 56 0 1.30422e-19 $X=14.225 $Y=1.63
c270 46 0 1.47605e-19 $X=10.695 $Y=1.525
c271 17 0 4.60399e-20 $X=9.86 $Y=1.435
c272 13 0 8.84733e-20 $X=7.09 $Y=2.635
c273 9 0 1.33662e-19 $X=6.31 $Y=0.84
r274 82 84 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=12.855 $Y=1.65
+ $X2=13.02 $Y2=1.65
r275 82 83 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.855
+ $Y=1.65 $X2=12.855 $Y2=1.65
r276 80 82 25.6147 $w=2.08e-07 $l=4.85e-07 $layer=LI1_cond $X=12.37 $Y=1.65
+ $X2=12.855 $Y2=1.65
r277 74 75 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=17.115 $Y=1.425
+ $X2=17.115 $Y2=1.955
r278 72 75 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=17.03 $Y=2.04
+ $X2=17.115 $Y2=1.955
r279 72 73 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=17.03 $Y=2.04
+ $X2=16.595 $Y2=2.04
r280 68 73 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=16.47 $Y=2.125
+ $X2=16.595 $Y2=2.04
r281 68 70 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=16.47 $Y=2.125
+ $X2=16.47 $Y2=2.84
r282 66 74 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=17.03 $Y=1.34
+ $X2=17.115 $Y2=1.425
r283 66 67 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=17.03 $Y=1.34
+ $X2=16.085 $Y2=1.34
r284 63 67 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=15.92 $Y=1.255
+ $X2=16.085 $Y2=1.34
r285 63 65 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=15.92 $Y=1.255
+ $X2=15.92 $Y2=0.765
r286 62 65 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=15.92 $Y=0.705
+ $X2=15.92 $Y2=0.765
r287 60 62 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=15.755 $Y=0.62
+ $X2=15.92 $Y2=0.705
r288 60 61 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=15.755 $Y=0.62
+ $X2=14.395 $Y2=0.62
r289 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.31 $Y=0.705
+ $X2=14.395 $Y2=0.62
r290 58 59 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=14.31 $Y=0.705
+ $X2=14.31 $Y2=1.545
r291 56 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.225 $Y=1.63
+ $X2=14.31 $Y2=1.545
r292 56 84 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=14.225 $Y=1.63
+ $X2=13.02 $Y2=1.63
r293 55 80 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=12.37 $Y=1.545
+ $X2=12.37 $Y2=1.65
r294 54 55 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=12.37 $Y=0.435
+ $X2=12.37 $Y2=1.545
r295 52 88 13.1721 $w=3.8e-07 $l=9e-08 $layer=POLY_cond $X=12.175 $Y=1.645
+ $X2=12.085 $Y2=1.645
r296 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.175
+ $Y=1.65 $X2=12.175 $Y2=1.65
r297 49 80 4.48918 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=12.285 $Y=1.65
+ $X2=12.37 $Y2=1.65
r298 49 51 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=12.285 $Y=1.65
+ $X2=12.175 $Y2=1.65
r299 47 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.285 $Y=0.35
+ $X2=12.37 $Y2=0.435
r300 47 48 98.1872 $w=1.68e-07 $l=1.505e-06 $layer=LI1_cond $X=12.285 $Y=0.35
+ $X2=10.78 $Y2=0.35
r301 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.695 $Y=0.435
+ $X2=10.78 $Y2=0.35
r302 45 46 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=10.695 $Y=0.435
+ $X2=10.695 $Y2=1.525
r303 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.925
+ $Y=1.61 $X2=9.925 $Y2=1.61
r304 41 43 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=7.605 $Y=1.61
+ $X2=9.925 $Y2=1.61
r305 40 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.61 $Y=1.61
+ $X2=10.695 $Y2=1.525
r306 40 43 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=10.61 $Y=1.61
+ $X2=9.925 $Y2=1.61
r307 39 78 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.52 $Y=1.915
+ $X2=7.52 $Y2=2
r308 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.52 $Y=1.695
+ $X2=7.605 $Y2=1.61
r309 38 39 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=7.52 $Y=1.695
+ $X2=7.52 $Y2=1.915
r310 36 85 7.30303 $w=5.28e-07 $l=8e-08 $layer=POLY_cond $X=7.07 $Y=2.11
+ $X2=7.07 $Y2=2.03
r311 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.115
+ $Y=2.11 $X2=7.115 $Y2=2.11
r312 33 78 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.115 $Y=2
+ $X2=7.52 $Y2=2
r313 33 35 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=7.115 $Y=2.085
+ $X2=7.115 $Y2=2.11
r314 29 83 60.0061 $w=3.8e-07 $l=4.1e-07 $layer=POLY_cond $X=12.445 $Y=1.645
+ $X2=12.855 $Y2=1.645
r315 29 52 39.5162 $w=3.8e-07 $l=2.7e-07 $layer=POLY_cond $X=12.445 $Y=1.645
+ $X2=12.175 $Y2=1.645
r316 29 31 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=12.445 $Y=1.455
+ $X2=12.445 $Y2=1.115
r317 27 88 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=12.085 $Y=1.835
+ $X2=12.085 $Y2=1.645
r318 27 28 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=12.085 $Y=1.835
+ $X2=12.085 $Y2=2.155
r319 24 28 40.618 $w=5.34e-07 $l=6.257e-07 $layer=POLY_cond $X=11.665 $Y=2.605
+ $X2=12.085 $Y2=2.155
r320 24 26 58.804 $w=5e-07 $l=6.1e-07 $layer=POLY_cond $X=11.665 $Y=2.605
+ $X2=11.665 $Y2=3.215
r321 20 44 60.3609 $w=9.45e-07 $l=1.09955e-06 $layer=POLY_cond $X=10.01 $Y=2.585
+ $X2=9.745 $Y2=1.61
r322 20 22 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=10.01 $Y=2.585
+ $X2=10.01 $Y2=3.09
r323 17 44 19.5567 $w=9.45e-07 $l=2.25278e-07 $layer=POLY_cond $X=9.86 $Y=1.435
+ $X2=9.745 $Y2=1.61
r324 17 19 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.86 $Y=1.435 $X2=9.86
+ $Y2=1.115
r325 13 36 48.1131 $w=5.28e-07 $l=5.34907e-07 $layer=POLY_cond $X=7.09 $Y=2.635
+ $X2=7.07 $Y2=2.11
r326 13 15 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.09 $Y=2.635
+ $X2=7.09 $Y2=3.415
r327 11 85 29.6317 $w=1.7e-07 $l=2.7e-07 $layer=POLY_cond $X=6.8 $Y=2.03
+ $X2=7.07 $Y2=2.03
r328 11 12 101.474 $w=1.7e-07 $l=2.4e-07 $layer=POLY_cond $X=6.8 $Y=2.03
+ $X2=6.56 $Y2=2.03
r329 7 12 36.4687 $w=1.7e-07 $l=2.89396e-07 $layer=POLY_cond $X=6.31 $Y=1.945
+ $X2=6.56 $Y2=2.03
r330 7 9 118.242 $w=5e-07 $l=1.105e-06 $layer=POLY_cond $X=6.31 $Y=1.945
+ $X2=6.31 $Y2=0.84
r331 2 70 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=16.29
+ $Y=2.715 $X2=16.43 $Y2=2.84
r332 1 65 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=15.795
+ $Y=0.555 $X2=15.92 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%A_1510_100# 1 2 9 13 17 21 24 26 28 29 30
+ 31 35
c106 31 0 6.08432e-20 $X=11.045 $Y=1.96
c107 28 0 5.57103e-20 $X=7.95 $Y=2.035
r108 32 35 9.4665 $w=2.78e-07 $l=2.3e-07 $layer=LI1_cond $X=11.045 $Y=2.815
+ $X2=11.275 $Y2=2.815
r109 29 39 49.2965 $w=5.85e-07 $l=5.25e-07 $layer=POLY_cond $X=7.842 $Y=2.035
+ $X2=7.842 $Y2=2.56
r110 29 38 18.2007 $w=5.85e-07 $l=1.85e-07 $layer=POLY_cond $X=7.842 $Y=2.035
+ $X2=7.842 $Y2=1.85
r111 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.95
+ $Y=2.035 $X2=7.95 $Y2=2.035
r112 26 32 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=11.045 $Y=2.675
+ $X2=11.045 $Y2=2.815
r113 25 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.045 $Y=2.045
+ $X2=11.045 $Y2=1.96
r114 25 26 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=11.045 $Y=2.045
+ $X2=11.045 $Y2=2.675
r115 24 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.045 $Y=1.875
+ $X2=11.045 $Y2=1.96
r116 24 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.045 $Y=1.875
+ $X2=11.045 $Y2=1.285
r117 19 30 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=11.142 $Y=1.103
+ $X2=11.142 $Y2=1.285
r118 19 21 12.7242 $w=3.63e-07 $l=4.03e-07 $layer=LI1_cond $X=11.142 $Y=1.103
+ $X2=11.142 $Y2=0.7
r119 18 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.115 $Y=1.96
+ $X2=7.95 $Y2=1.96
r120 17 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.96 $Y=1.96
+ $X2=11.045 $Y2=1.96
r121 17 18 185.61 $w=1.68e-07 $l=2.845e-06 $layer=LI1_cond $X=10.96 $Y=1.96
+ $X2=8.115 $Y2=1.96
r122 13 39 91.49 $w=5e-07 $l=8.55e-07 $layer=POLY_cond $X=7.8 $Y=3.415 $X2=7.8
+ $Y2=2.56
r123 9 38 108.076 $w=5e-07 $l=1.01e-06 $layer=POLY_cond $X=7.8 $Y=0.84 $X2=7.8
+ $Y2=1.85
r124 2 35 600 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_PDIFF $count=1 $X=11.135
+ $Y=2.715 $X2=11.275 $Y2=2.855
r125 1 21 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=11.02
+ $Y=0.575 $X2=11.16 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%RESET_B 3 8 9 10 14 17 19 22 23 25 26 27
+ 28 31 37 41 42 44 45 47 50 54 56
c209 42 0 3.32014e-19 $X=4.135 $Y=2.1
c210 19 0 5.7967e-21 $X=4.2 $Y=1.565
c211 3 0 1.36153e-20 $X=3.86 $Y=3.455
r212 58 73 2.83207 $w=2.35e-07 $l=1.68e-07 $layer=LI1_cond $X=4.3 $Y=2.407
+ $X2=4.132 $Y2=2.407
r213 53 56 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=14.27 $Y=2.025
+ $X2=14.27 $Y2=2.925
r214 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.205
+ $Y=2.025 $X2=14.205 $Y2=2.025
r215 50 53 97.3754 $w=5e-07 $l=9.1e-07 $layer=POLY_cond $X=14.27 $Y=1.115
+ $X2=14.27 $Y2=2.025
r216 44 47 110.751 $w=5e-07 $l=1.035e-06 $layer=POLY_cond $X=8.66 $Y=2.38
+ $X2=8.66 $Y2=3.415
r217 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.595
+ $Y=2.38 $X2=8.595 $Y2=2.38
r218 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.135
+ $Y=2.1 $X2=4.135 $Y2=2.1
r219 38 54 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=14.205 $Y=2.405
+ $X2=14.205 $Y2=2.025
r220 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=2.405
+ $X2=14.16 $Y2=2.405
r221 35 45 7.24924 $w=3.08e-07 $l=1.95e-07 $layer=LI1_cond $X=8.4 $Y=2.38
+ $X2=8.595 $Y2=2.38
r222 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.405
+ $X2=8.4 $Y2=2.405
r223 31 58 12.7504 $w=2.33e-07 $l=2.6e-07 $layer=LI1_cond $X=4.56 $Y=2.407
+ $X2=4.3 $Y2=2.407
r224 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=2.405
+ $X2=4.56 $Y2=2.405
r225 28 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.545 $Y=2.405
+ $X2=8.4 $Y2=2.405
r226 27 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.015 $Y=2.405
+ $X2=14.16 $Y2=2.405
r227 27 28 6.76979 $w=1.4e-07 $l=5.47e-06 $layer=MET1_cond $X=14.015 $Y=2.405
+ $X2=8.545 $Y2=2.405
r228 26 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=2.405
+ $X2=4.56 $Y2=2.405
r229 25 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=2.405
+ $X2=8.4 $Y2=2.405
r230 25 26 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=8.255 $Y=2.405
+ $X2=4.705 $Y2=2.405
r231 23 73 0.0688026 $w=3.33e-07 $l=2e-09 $layer=LI1_cond $X=4.132 $Y=2.405
+ $X2=4.132 $Y2=2.407
r232 23 42 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=4.132 $Y=2.405
+ $X2=4.132 $Y2=2.1
r233 22 44 85.0697 $w=5e-07 $l=7.95e-07 $layer=POLY_cond $X=8.66 $Y=1.585
+ $X2=8.66 $Y2=2.38
r234 21 22 37.8636 $w=6.5e-07 $l=4.6e-07 $layer=POLY_cond $X=8.585 $Y=1.125
+ $X2=8.585 $Y2=1.585
r235 19 41 83.4372 $w=3.7e-07 $l=5.35e-07 $layer=POLY_cond $X=4.135 $Y=1.565
+ $X2=4.135 $Y2=2.1
r236 16 41 69.401 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=4.135 $Y=2.545
+ $X2=4.135 $Y2=2.1
r237 16 17 64.7199 $w=5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.965 $Y=2.545
+ $X2=3.965 $Y2=3.115
r238 14 21 30.4967 $w=5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.51 $Y=0.84
+ $X2=8.51 $Y2=1.125
r239 11 14 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=8.51 $Y=0.29 $X2=8.51
+ $Y2=0.84
r240 9 11 38.6381 $w=1.5e-07 $l=2.85044e-07 $layer=POLY_cond $X=8.26 $Y=0.215
+ $X2=8.51 $Y2=0.29
r241 9 10 1953.64 $w=1.5e-07 $l=3.81e-06 $layer=POLY_cond $X=8.26 $Y=0.215
+ $X2=4.45 $Y2=0.215
r242 6 19 30.478 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.2 $Y=1.315 $X2=4.2
+ $Y2=1.565
r243 6 8 50.8278 $w=5e-07 $l=4.75e-07 $layer=POLY_cond $X=4.2 $Y=1.315 $X2=4.2
+ $Y2=0.84
r244 5 10 38.6381 $w=1.5e-07 $l=2.85044e-07 $layer=POLY_cond $X=4.2 $Y=0.29
+ $X2=4.45 $Y2=0.215
r245 5 8 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.2 $Y=0.29 $X2=4.2
+ $Y2=0.84
r246 3 17 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.86 $Y=3.455 $X2=3.86
+ $Y2=3.115
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%A_1312_126# 1 2 3 12 14 16 18 21 23 27 30
+ 31 32 36 38 39 40
r129 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.655
+ $Y=2.39 $X2=10.655 $Y2=2.39
r130 40 43 3.17915 $w=2.88e-07 $l=8e-08 $layer=LI1_cond $X=10.635 $Y=2.31
+ $X2=10.635 $Y2=2.39
r131 33 36 2.4262 $w=3.78e-07 $l=8e-08 $layer=LI1_cond $X=6.62 $Y=0.805 $X2=6.7
+ $Y2=0.805
r132 31 40 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=10.49 $Y=2.31
+ $X2=10.635 $Y2=2.31
r133 31 32 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=10.49 $Y=2.31
+ $X2=9.215 $Y2=2.31
r134 30 39 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=9.13 $Y=2.715
+ $X2=9.05 $Y2=2.8
r135 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.13 $Y=2.395
+ $X2=9.215 $Y2=2.31
r136 29 30 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.13 $Y=2.395
+ $X2=9.13 $Y2=2.715
r137 25 39 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.05 $Y=2.885
+ $X2=9.05 $Y2=2.8
r138 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.05 $Y=2.885
+ $X2=9.05 $Y2=3.35
r139 24 38 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.865 $Y=2.8
+ $X2=6.7 $Y2=2.8
r140 23 39 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.885 $Y=2.8
+ $X2=9.05 $Y2=2.8
r141 23 24 131.786 $w=1.68e-07 $l=2.02e-06 $layer=LI1_cond $X=8.885 $Y=2.8
+ $X2=6.865 $Y2=2.8
r142 19 38 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.7 $Y=2.885 $X2=6.7
+ $Y2=2.8
r143 19 21 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.7 $Y=2.885
+ $X2=6.7 $Y2=3.35
r144 18 38 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.62 $Y=2.715
+ $X2=6.7 $Y2=2.8
r145 17 33 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.62 $Y=0.995
+ $X2=6.62 $Y2=0.805
r146 17 18 112.214 $w=1.68e-07 $l=1.72e-06 $layer=LI1_cond $X=6.62 $Y=0.995
+ $X2=6.62 $Y2=2.715
r147 14 44 19.5756 $w=5.38e-07 $l=2.53121e-07 $layer=POLY_cond $X=10.885
+ $Y=2.605 $X2=10.802 $Y2=2.39
r148 14 16 58.804 $w=5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.885 $Y=2.605
+ $X2=10.885 $Y2=3.215
r149 10 44 61.6834 $w=5.38e-07 $l=7.00817e-07 $layer=POLY_cond $X=10.77 $Y=1.705
+ $X2=10.802 $Y2=2.39
r150 10 12 80.7895 $w=5e-07 $l=7.55e-07 $layer=POLY_cond $X=10.77 $Y=1.705
+ $X2=10.77 $Y2=0.95
r151 3 27 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.91
+ $Y=3.205 $X2=9.05 $Y2=3.35
r152 2 21 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.56
+ $Y=3.205 $X2=6.7 $Y2=3.35
r153 1 36 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=6.56
+ $Y=0.63 $X2=6.7 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%A_2616_417# 1 2 9 13 16 19 20 23 26 27 28
+ 29 31 36
c92 28 0 1.08219e-19 $X=14.745 $Y=1.26
r93 31 33 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=15.37 $Y=1.115
+ $X2=15.37 $Y2=1.26
r94 27 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.205 $Y=1.26
+ $X2=15.37 $Y2=1.26
r95 27 28 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=15.205 $Y=1.26
+ $X2=14.745 $Y2=1.26
r96 26 29 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=14.66 $Y=2.67
+ $X2=14.62 $Y2=2.755
r97 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.66 $Y=1.345
+ $X2=14.745 $Y2=1.26
r98 25 26 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=14.66 $Y=1.345
+ $X2=14.66 $Y2=2.67
r99 21 29 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=14.62 $Y=2.84
+ $X2=14.62 $Y2=2.755
r100 21 23 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=14.62 $Y=2.84
+ $X2=14.62 $Y2=2.925
r101 19 29 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.495 $Y=2.755
+ $X2=14.62 $Y2=2.755
r102 19 20 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=14.495 $Y=2.755
+ $X2=13.71 $Y2=2.755
r103 17 36 100.051 $w=5e-07 $l=9.35e-07 $layer=POLY_cond $X=13.48 $Y=2.05
+ $X2=13.48 $Y2=1.115
r104 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.545
+ $Y=2.05 $X2=13.545 $Y2=2.05
r105 14 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.545 $Y=2.67
+ $X2=13.71 $Y2=2.755
r106 14 16 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=13.545 $Y=2.67
+ $X2=13.545 $Y2=2.05
r107 12 17 3.74521 $w=5e-07 $l=3.5e-08 $layer=POLY_cond $X=13.48 $Y=2.085
+ $X2=13.48 $Y2=2.05
r108 12 13 41.1561 $w=6.5e-07 $l=5e-07 $layer=POLY_cond $X=13.405 $Y=2.085
+ $X2=13.405 $Y2=2.585
r109 9 13 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=13.33 $Y=2.925
+ $X2=13.33 $Y2=2.585
r110 2 23 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=14.52
+ $Y=2.715 $X2=14.66 $Y2=2.925
r111 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=15.23
+ $Y=0.905 $X2=15.37 $Y2=1.115
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%A_2360_115# 1 2 9 13 17 21 23 24 27 30 33
+ 35 36 38 39 40 42 43 44 45 46 48 51 55 62
c177 62 0 1.30422e-19 $X=15.09 $Y=1.77
c178 23 0 9.71226e-20 $X=17.37 $Y=1.795
r179 62 68 50.2236 $w=5.7e-07 $l=5.25e-07 $layer=POLY_cond $X=15.015 $Y=1.77
+ $X2=15.015 $Y2=2.295
r180 62 67 30.512 $w=5.7e-07 $l=3.15e-07 $layer=POLY_cond $X=15.015 $Y=1.77
+ $X2=15.015 $Y2=1.455
r181 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=15.09
+ $Y=1.77 $X2=15.09 $Y2=1.77
r182 55 56 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=11.882 $Y=1.2
+ $X2=11.882 $Y2=1.365
r183 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.685
+ $Y=1.69 $X2=16.685 $Y2=1.69
r184 49 61 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.255 $Y=1.69
+ $X2=15.09 $Y2=1.69
r185 49 51 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=15.255 $Y=1.69
+ $X2=16.685 $Y2=1.69
r186 48 63 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=15.01 $Y=3.355
+ $X2=15.01 $Y2=2.275
r187 46 63 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=15.09 $Y=2.11
+ $X2=15.09 $Y2=2.275
r188 45 61 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.09 $Y=1.775
+ $X2=15.09 $Y2=1.69
r189 45 46 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=15.09 $Y=1.775
+ $X2=15.09 $Y2=2.11
r190 43 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.925 $Y=3.44
+ $X2=15.01 $Y2=3.355
r191 43 44 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=14.925 $Y=3.44
+ $X2=14.315 $Y2=3.44
r192 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.23 $Y=3.355
+ $X2=14.315 $Y2=3.44
r193 41 42 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=14.23 $Y=3.19
+ $X2=14.23 $Y2=3.355
r194 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.145 $Y=3.105
+ $X2=14.23 $Y2=3.19
r195 39 40 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=14.145 $Y=3.105
+ $X2=13.2 $Y2=3.105
r196 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.115 $Y=3.02
+ $X2=13.2 $Y2=3.105
r197 37 38 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=13.115 $Y=2.105
+ $X2=13.115 $Y2=3.02
r198 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.03 $Y=2.02
+ $X2=13.115 $Y2=2.105
r199 35 36 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=13.03 $Y=2.02
+ $X2=12.3 $Y2=2.02
r200 31 36 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=12.135 $Y=2.02
+ $X2=12.3 $Y2=2.02
r201 31 57 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=12.135 $Y=2.02
+ $X2=11.745 $Y2=2.02
r202 31 33 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=12.135 $Y=2.105
+ $X2=12.135 $Y2=2.865
r203 30 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.745 $Y=1.935
+ $X2=11.745 $Y2=2.02
r204 30 56 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=11.745 $Y=1.935
+ $X2=11.745 $Y2=1.365
r205 25 55 1.47616 $w=4.43e-07 $l=5.7e-08 $layer=LI1_cond $X=11.882 $Y=1.143
+ $X2=11.882 $Y2=1.2
r206 25 27 11.4726 $w=4.43e-07 $l=4.43e-07 $layer=LI1_cond $X=11.882 $Y=1.143
+ $X2=11.882 $Y2=0.7
r207 23 52 63.1888 $w=5.8e-07 $l=6.85e-07 $layer=POLY_cond $X=17.37 $Y=1.795
+ $X2=16.685 $Y2=1.795
r208 23 24 3.21582 $w=5.8e-07 $l=2.7e-07 $layer=POLY_cond $X=17.37 $Y=1.795
+ $X2=17.64 $Y2=1.795
r209 19 24 23.051 $w=5e-07 $l=2.99833e-07 $layer=POLY_cond $X=17.66 $Y=1.505
+ $X2=17.64 $Y2=1.795
r210 19 21 46.0125 $w=5e-07 $l=4.3e-07 $layer=POLY_cond $X=17.66 $Y=1.505
+ $X2=17.66 $Y2=1.075
r211 15 24 23.051 $w=5e-07 $l=2.99833e-07 $layer=POLY_cond $X=17.62 $Y=2.085
+ $X2=17.64 $Y2=1.795
r212 15 17 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=17.62 $Y=2.085
+ $X2=17.62 $Y2=2.59
r213 13 68 67.4137 $w=5e-07 $l=6.3e-07 $layer=POLY_cond $X=15.05 $Y=2.925
+ $X2=15.05 $Y2=2.295
r214 9 67 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=14.98 $Y=1.115
+ $X2=14.98 $Y2=1.455
r215 2 33 600 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_PDIFF $count=1 $X=11.915
+ $Y=2.715 $X2=12.135 $Y2=2.865
r216 1 55 182 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_NDIFF $count=1 $X=11.8
+ $Y=0.575 $X2=11.94 $Y2=1.2
r217 1 27 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=11.8
+ $Y=0.575 $X2=11.94 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%CLK 1 3 9 12 13 15
c37 13 0 9.71226e-20 $X=15.975 $Y=2.05
r38 12 15 111.286 $w=5e-07 $l=1.04e-06 $layer=POLY_cond $X=16.04 $Y=2.05
+ $X2=16.04 $Y2=3.09
r39 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=15.975
+ $Y=2.05 $X2=15.975 $Y2=2.05
r40 9 13 8.3061 $w=5.38e-07 $l=3.75e-07 $layer=LI1_cond $X=15.6 $Y=2.225
+ $X2=15.975 $Y2=2.225
r41 5 12 83.9996 $w=5e-07 $l=7.85e-07 $layer=POLY_cond $X=16.04 $Y=1.265
+ $X2=16.04 $Y2=2.05
r42 1 5 114.158 $w=1.7e-07 $l=2.7e-07 $layer=POLY_cond $X=16.31 $Y=1.18
+ $X2=16.04 $Y2=1.18
r43 1 3 31.812 $w=5e-07 $l=3.3e-07 $layer=POLY_cond $X=16.31 $Y=1.095 $X2=16.31
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%A_3417_443# 1 2 9 13 15 20 25 26 29 30 32
c51 32 0 1.91511e-19 $X=17.465 $Y=1.65
r52 29 30 7.45324 $w=4.83e-07 $l=8.5e-08 $layer=LI1_cond $X=17.307 $Y=2.39
+ $X2=17.307 $Y2=2.305
r53 26 35 44.7573 $w=5.2e-07 $l=4.35e-07 $layer=POLY_cond $X=18.525 $Y=1.65
+ $X2=18.525 $Y2=2.085
r54 26 34 24.1792 $w=5.2e-07 $l=2.35e-07 $layer=POLY_cond $X=18.525 $Y=1.65
+ $X2=18.525 $Y2=1.415
r55 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=18.45
+ $Y=1.65 $X2=18.45 $Y2=1.65
r56 23 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=17.55 $Y=1.65
+ $X2=17.465 $Y2=1.65
r57 23 25 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=17.55 $Y=1.65
+ $X2=18.45 $Y2=1.65
r58 21 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.465 $Y=1.815
+ $X2=17.465 $Y2=1.65
r59 21 30 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=17.465 $Y=1.815
+ $X2=17.465 $Y2=2.305
r60 20 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.465 $Y=1.485
+ $X2=17.465 $Y2=1.65
r61 19 20 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=17.465 $Y=1.075
+ $X2=17.465 $Y2=1.485
r62 15 19 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=17.38 $Y=0.95
+ $X2=17.465 $Y2=1.075
r63 15 17 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=17.38 $Y=0.95
+ $X2=17.27 $Y2=0.95
r64 13 34 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=18.535 $Y=0.91
+ $X2=18.535 $Y2=1.415
r65 9 35 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=18.515 $Y=2.965
+ $X2=18.515 $Y2=2.085
r66 2 29 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=17.085
+ $Y=2.215 $X2=17.23 $Y2=2.39
r67 1 17 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=17.125
+ $Y=0.865 $X2=17.27 $Y2=0.99
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%A_65_649# 1 2 3 4 5 17 20 22 23 24 27 28
+ 30 33 34 35 39 40 41 43 44 45 46 49 52 55 56 57
c151 22 0 9.7103e-20 $X=1.295 $Y=1.775
r152 56 57 140.92 $w=1.68e-07 $l=2.16e-06 $layer=LI1_cond $X=5.92 $Y=1.005
+ $X2=5.92 $Y2=3.165
r153 50 52 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=5.88 $Y=3.635
+ $X2=5.88 $Y2=3.415
r154 49 57 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.88 $Y=3.29
+ $X2=5.88 $Y2=3.165
r155 49 52 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.88 $Y=3.29
+ $X2=5.88 $Y2=3.415
r156 46 56 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.88 $Y=0.88
+ $X2=5.88 $Y2=1.005
r157 46 48 1.952 $w=2.5e-07 $l=4e-08 $layer=LI1_cond $X=5.88 $Y=0.88 $X2=5.88
+ $Y2=0.84
r158 44 50 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.755 $Y=3.72
+ $X2=5.88 $Y2=3.635
r159 44 45 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.755 $Y=3.72
+ $X2=4.975 $Y2=3.72
r160 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.89 $Y=3.635
+ $X2=4.975 $Y2=3.72
r161 42 43 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.89 $Y=3.225
+ $X2=4.89 $Y2=3.635
r162 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.805 $Y=3.14
+ $X2=4.89 $Y2=3.225
r163 40 41 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=4.805 $Y=3.14
+ $X2=3.555 $Y2=3.14
r164 37 39 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.47 $Y=3.535
+ $X2=3.47 $Y2=3.455
r165 36 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.47 $Y=3.225
+ $X2=3.555 $Y2=3.14
r166 36 39 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.47 $Y=3.225
+ $X2=3.47 $Y2=3.455
r167 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.385 $Y=3.62
+ $X2=3.47 $Y2=3.535
r168 34 35 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.385 $Y=3.62
+ $X2=2.73 $Y2=3.62
r169 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.645 $Y=3.535
+ $X2=2.73 $Y2=3.62
r170 32 33 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.645 $Y=3.275
+ $X2=2.645 $Y2=3.535
r171 28 30 32.8446 $w=2.98e-07 $l=8.55e-07 $layer=LI1_cond $X=1.465 $Y=0.765
+ $X2=2.32 $Y2=0.765
r172 26 28 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.38 $Y=0.915
+ $X2=1.465 $Y2=0.765
r173 26 27 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.38 $Y=0.915
+ $X2=1.38 $Y2=1.69
r174 25 55 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=3.19
+ $X2=0.47 $Y2=3.19
r175 24 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.56 $Y=3.19
+ $X2=2.645 $Y2=3.275
r176 24 25 125.588 $w=1.68e-07 $l=1.925e-06 $layer=LI1_cond $X=2.56 $Y=3.19
+ $X2=0.635 $Y2=3.19
r177 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.295 $Y=1.775
+ $X2=1.38 $Y2=1.69
r178 22 23 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.295 $Y=1.775
+ $X2=0.475 $Y2=1.775
r179 18 55 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.47 $Y=3.275
+ $X2=0.47 $Y2=3.19
r180 18 20 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.47 $Y=3.275
+ $X2=0.47 $Y2=3.455
r181 17 55 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.39 $Y=3.105
+ $X2=0.47 $Y2=3.19
r182 16 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.39 $Y=1.86
+ $X2=0.475 $Y2=1.775
r183 16 17 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=0.39 $Y=1.86
+ $X2=0.39 $Y2=3.105
r184 5 52 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.775
+ $Y=3.205 $X2=5.92 $Y2=3.415
r185 4 39 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.33
+ $Y=3.245 $X2=3.47 $Y2=3.455
r186 3 20 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=3.245 $X2=0.47 $Y2=3.455
r187 2 48 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.795
+ $Y=0.63 $X2=5.92 $Y2=0.84
r188 1 30 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=2.18
+ $Y=0.63 $X2=2.32 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%VPWR 1 2 3 4 5 6 7 22 31 41 49 60 68 73 84
+ 92
c144 41 0 1.47013e-19 $X=4.54 $Y=3.59
r145 90 92 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=17.825 $Y=3.63
+ $X2=18.545 $Y2=3.63
r146 89 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=18.545 $Y=3.59
+ $X2=18.545 $Y2=3.59
r147 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.825 $Y=3.59
+ $X2=17.825 $Y2=3.59
r148 87 89 5.56374 $w=9.08e-07 $l=4.15e-07 $layer=LI1_cond $X=18.185 $Y=3.175
+ $X2=18.185 $Y2=3.59
r149 84 87 11.1945 $w=9.08e-07 $l=8.35e-07 $layer=LI1_cond $X=18.185 $Y=2.34
+ $X2=18.185 $Y2=3.175
r150 81 90 0.669915 $w=3.7e-07 $l=1.745e-06 $layer=MET1_cond $X=16.08 $Y=3.63
+ $X2=17.825 $Y2=3.63
r151 79 81 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=15.36 $Y=3.63
+ $X2=16.08 $Y2=3.63
r152 78 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.08 $Y=3.59
+ $X2=16.08 $Y2=3.59
r153 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.36 $Y=3.59
+ $X2=15.36 $Y2=3.59
r154 76 78 3.42697 $w=8.88e-07 $l=2.5e-07 $layer=LI1_cond $X=15.72 $Y=3.34
+ $X2=15.72 $Y2=3.59
r155 73 76 6.85393 $w=8.88e-07 $l=5e-07 $layer=LI1_cond $X=15.72 $Y=2.84
+ $X2=15.72 $Y2=3.34
r156 70 79 0.579697 $w=3.7e-07 $l=1.51e-06 $layer=MET1_cond $X=13.85 $Y=3.63
+ $X2=15.36 $Y2=3.63
r157 68 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.85 $Y=3.59
+ $X2=13.85 $Y2=3.59
r158 65 70 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=13.13 $Y=3.63
+ $X2=13.85 $Y2=3.63
r159 64 68 23.0489 $w=3.33e-07 $l=6.7e-07 $layer=LI1_cond $X=13.13 $Y=3.537
+ $X2=13.8 $Y2=3.537
r160 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.13 $Y=3.59
+ $X2=13.13 $Y2=3.59
r161 61 65 0.8945 $w=3.7e-07 $l=2.33e-06 $layer=MET1_cond $X=10.8 $Y=3.63
+ $X2=13.13 $Y2=3.63
r162 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=3.6
+ $X2=10.8 $Y2=3.6
r163 58 60 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=10.495 $Y=3.61
+ $X2=10.8 $Y2=3.61
r164 55 61 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.08 $Y=3.63
+ $X2=10.8 $Y2=3.63
r165 54 58 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=10.08 $Y=3.61
+ $X2=10.495 $Y2=3.61
r166 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.08 $Y=3.6
+ $X2=10.08 $Y2=3.6
r167 49 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.24 $Y=3.59
+ $X2=8.24 $Y2=3.59
r168 46 51 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.52 $Y=3.63
+ $X2=8.24 $Y2=3.63
r169 45 49 26.6254 $w=2.88e-07 $l=6.7e-07 $layer=LI1_cond $X=7.52 $Y=3.56
+ $X2=8.19 $Y2=3.56
r170 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.52 $Y=3.59
+ $X2=7.52 $Y2=3.59
r171 42 46 1.14404 $w=3.7e-07 $l=2.98e-06 $layer=MET1_cond $X=4.54 $Y=3.63
+ $X2=7.52 $Y2=3.63
r172 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.54 $Y=3.59
+ $X2=4.54 $Y2=3.59
r173 39 41 10.9482 $w=2.98e-07 $l=2.85e-07 $layer=LI1_cond $X=4.255 $Y=3.555
+ $X2=4.54 $Y2=3.555
r174 36 42 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.82 $Y=3.63
+ $X2=4.54 $Y2=3.63
r175 35 39 16.7104 $w=2.98e-07 $l=4.35e-07 $layer=LI1_cond $X=3.82 $Y=3.555
+ $X2=4.255 $Y2=3.555
r176 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.82 $Y=3.59
+ $X2=3.82 $Y2=3.59
r177 32 36 0.600812 $w=3.7e-07 $l=1.565e-06 $layer=MET1_cond $X=2.255 $Y=3.63
+ $X2=3.82 $Y2=3.63
r178 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.255 $Y=3.59
+ $X2=2.255 $Y2=3.59
r179 29 31 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.96 $Y=3.58
+ $X2=2.255 $Y2=3.58
r180 26 32 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.535 $Y=3.63
+ $X2=2.255 $Y2=3.63
r181 25 29 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=1.535 $Y=3.58
+ $X2=1.96 $Y2=3.58
r182 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.535 $Y=3.59
+ $X2=1.535 $Y2=3.59
r183 22 55 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=9.6 $Y=3.63
+ $X2=10.08 $Y2=3.63
r184 22 51 0.522111 $w=3.7e-07 $l=1.36e-06 $layer=MET1_cond $X=9.6 $Y=3.63
+ $X2=8.24 $Y2=3.63
r185 7 87 300 $w=1.7e-07 $l=1.08e-06 $layer=licon1_PDIFF $count=2 $X=17.87
+ $Y=2.215 $X2=18.125 $Y2=3.175
r186 7 84 300 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=2 $X=17.87
+ $Y=2.215 $X2=18.125 $Y2=2.34
r187 6 76 600 $w=1.7e-07 $l=7.80625e-07 $layer=licon1_PDIFF $count=1 $X=15.3
+ $Y=2.715 $X2=15.65 $Y2=3.34
r188 6 73 600 $w=1.7e-07 $l=4.07738e-07 $layer=licon1_PDIFF $count=1 $X=15.3
+ $Y=2.715 $X2=15.65 $Y2=2.84
r189 5 68 600 $w=1.7e-07 $l=8.42852e-07 $layer=licon1_PDIFF $count=1 $X=13.58
+ $Y=2.715 $X2=13.8 $Y2=3.455
r190 4 58 600 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=10.26
+ $Y=2.715 $X2=10.495 $Y2=3.57
r191 3 49 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=8.05
+ $Y=3.205 $X2=8.19 $Y2=3.5
r192 2 39 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=4.11
+ $Y=3.245 $X2=4.255 $Y2=3.515
r193 1 29 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.82
+ $Y=3.245 $X2=1.96 $Y2=3.54
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%Q 1 2 7 8 9 10 11 12 13 22
r14 13 40 20.1113 $w=2.53e-07 $l=4.45e-07 $layer=LI1_cond $X=18.947 $Y=3.145
+ $X2=18.947 $Y2=3.59
r15 12 13 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=18.947 $Y=2.775
+ $X2=18.947 $Y2=3.145
r16 11 12 19.6593 $w=2.53e-07 $l=4.35e-07 $layer=LI1_cond $X=18.947 $Y=2.34
+ $X2=18.947 $Y2=2.775
r17 10 11 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=18.947 $Y=2.035
+ $X2=18.947 $Y2=2.34
r18 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=18.947 $Y=1.665
+ $X2=18.947 $Y2=2.035
r19 8 9 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=18.947 $Y=1.295
+ $X2=18.947 $Y2=1.665
r20 7 8 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=18.947 $Y=0.925
+ $X2=18.947 $Y2=1.295
r21 7 22 11.0725 $w=2.53e-07 $l=2.45e-07 $layer=LI1_cond $X=18.947 $Y=0.925
+ $X2=18.947 $Y2=0.68
r22 2 40 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=18.765
+ $Y=2.215 $X2=18.905 $Y2=3.59
r23 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=18.765
+ $Y=2.215 $X2=18.905 $Y2=2.34
r24 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=18.785
+ $Y=0.535 $X2=18.925 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%noxref_23 1 2 9 11 12 15
r31 13 15 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=3.81 $Y=0.435
+ $X2=3.81 $Y2=0.84
r32 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.645 $Y=0.35
+ $X2=3.81 $Y2=0.435
r33 11 12 172.888 $w=1.68e-07 $l=2.65e-06 $layer=LI1_cond $X=3.645 $Y=0.35
+ $X2=0.995 $Y2=0.35
r34 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.83 $Y=0.435
+ $X2=0.995 $Y2=0.35
r35 7 9 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.83 $Y=0.435
+ $X2=0.83 $Y2=0.84
r36 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.63 $X2=3.81 $Y2=0.84
r37 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.685
+ $Y=0.63 $X2=0.83 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFRTP_1%VGND 1 2 3 4 5 6 19 22 31 40 49 58 65 69
r114 71 73 6.16703 $w=9.08e-07 $l=4.6e-07 $layer=LI1_cond $X=18.185 $Y=0.68
+ $X2=18.185 $Y2=1.14
r115 66 69 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=17.825 $Y=0.44
+ $X2=18.545 $Y2=0.44
r116 65 71 2.68132 $w=9.08e-07 $l=2e-07 $layer=LI1_cond $X=18.185 $Y=0.48
+ $X2=18.185 $Y2=0.68
r117 65 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=18.545 $Y=0.48
+ $X2=18.545 $Y2=0.48
r118 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.825 $Y=0.48
+ $X2=17.825 $Y2=0.48
r119 59 66 0.412698 $w=3.7e-07 $l=1.075e-06 $layer=MET1_cond $X=16.75 $Y=0.44
+ $X2=17.825 $Y2=0.44
r120 58 62 5.77767 $w=5.88e-07 $l=2.85e-07 $layer=LI1_cond $X=16.57 $Y=0.48
+ $X2=16.57 $Y2=0.765
r121 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.75 $Y=0.48
+ $X2=16.75 $Y2=0.48
r122 53 59 1.08645 $w=3.7e-07 $l=2.83e-06 $layer=MET1_cond $X=13.92 $Y=0.44
+ $X2=16.75 $Y2=0.44
r123 50 53 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=13.2 $Y=0.44
+ $X2=13.92 $Y2=0.44
r124 49 55 8.15474 $w=9.48e-07 $l=6.35e-07 $layer=LI1_cond $X=13.56 $Y=0.48
+ $X2=13.56 $Y2=1.115
r125 49 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.92 $Y=0.48
+ $X2=13.92 $Y2=0.48
r126 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=0.48
+ $X2=13.2 $Y2=0.48
r127 44 46 9.32536 $w=5.88e-07 $l=4.6e-07 $layer=LI1_cond $X=10.135 $Y=0.72
+ $X2=10.135 $Y2=1.18
r128 41 50 1.10757 $w=3.7e-07 $l=2.885e-06 $layer=MET1_cond $X=10.315 $Y=0.44
+ $X2=13.2 $Y2=0.44
r129 40 44 4.8654 $w=5.88e-07 $l=2.4e-07 $layer=LI1_cond $X=10.135 $Y=0.48
+ $X2=10.135 $Y2=0.72
r130 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.315 $Y=0.48
+ $X2=10.315 $Y2=0.48
r131 32 35 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.23 $Y=0.44
+ $X2=8.95 $Y2=0.44
r132 31 37 4.88 $w=9.48e-07 $l=3.8e-07 $layer=LI1_cond $X=8.59 $Y=0.48 $X2=8.59
+ $Y2=0.86
r133 31 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.95 $Y=0.48
+ $X2=8.95 $Y2=0.48
r134 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.23 $Y=0.48
+ $X2=8.23 $Y2=0.48
r135 26 32 1.24385 $w=3.7e-07 $l=3.24e-06 $layer=MET1_cond $X=4.99 $Y=0.44
+ $X2=8.23 $Y2=0.44
r136 23 26 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=4.27 $Y=0.44
+ $X2=4.99 $Y2=0.44
r137 22 28 4.62316 $w=9.48e-07 $l=3.6e-07 $layer=LI1_cond $X=4.63 $Y=0.48
+ $X2=4.63 $Y2=0.84
r138 22 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.99 $Y=0.48
+ $X2=4.99 $Y2=0.48
r139 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.27 $Y=0.48
+ $X2=4.27 $Y2=0.48
r140 19 41 0.274492 $w=3.7e-07 $l=7.15e-07 $layer=MET1_cond $X=9.6 $Y=0.44
+ $X2=10.315 $Y2=0.44
r141 19 35 0.249539 $w=3.7e-07 $l=6.5e-07 $layer=MET1_cond $X=9.6 $Y=0.44
+ $X2=8.95 $Y2=0.44
r142 6 73 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=17.91
+ $Y=0.865 $X2=18.145 $Y2=1.14
r143 6 71 182 $w=1.7e-07 $l=3.14166e-07 $layer=licon1_NDIFF $count=1 $X=17.91
+ $Y=0.865 $X2=18.145 $Y2=0.68
r144 5 62 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=16.56
+ $Y=0.555 $X2=16.7 $Y2=0.765
r145 4 55 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.73
+ $Y=0.905 $X2=13.87 $Y2=1.115
r146 3 46 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=10.11
+ $Y=0.905 $X2=10.345 $Y2=1.18
r147 3 44 182 $w=1.7e-07 $l=3.14166e-07 $layer=licon1_NDIFF $count=1 $X=10.11
+ $Y=0.905 $X2=10.345 $Y2=0.72
r148 2 37 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=8.76
+ $Y=0.63 $X2=8.9 $Y2=0.86
r149 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.45
+ $Y=0.63 $X2=4.59 $Y2=0.84
.ends

