* File: sky130_fd_sc_hvl__o21a_1.pxi.spice
* Created: Fri Aug 28 09:38:34 2020
* 
x_PM_SKY130_FD_SC_HVL__O21A_1%VNB N_VNB_M1000_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__O21A_1%VNB
x_PM_SKY130_FD_SC_HVL__O21A_1%VPB N_VPB_M1002_b VPB N_VPB_c_36_p VPB
+ PM_SKY130_FD_SC_HVL__O21A_1%VPB
x_PM_SKY130_FD_SC_HVL__O21A_1%A_83_87# N_A_83_87#_M1005_s N_A_83_87#_M1006_d
+ N_A_83_87#_M1000_g N_A_83_87#_M1002_g N_A_83_87#_c_70_n N_A_83_87#_c_71_n
+ N_A_83_87#_c_73_n N_A_83_87#_c_74_n N_A_83_87#_c_104_p N_A_83_87#_c_75_n
+ N_A_83_87#_c_76_n PM_SKY130_FD_SC_HVL__O21A_1%A_83_87#
x_PM_SKY130_FD_SC_HVL__O21A_1%B1 N_B1_M1006_g N_B1_M1005_g B1 B1 N_B1_c_129_n
+ N_B1_c_130_n PM_SKY130_FD_SC_HVL__O21A_1%B1
x_PM_SKY130_FD_SC_HVL__O21A_1%A2 N_A2_M1001_g N_A2_M1003_g A2 A2 A2 A2 A2
+ N_A2_c_165_n PM_SKY130_FD_SC_HVL__O21A_1%A2
x_PM_SKY130_FD_SC_HVL__O21A_1%A1 N_A1_M1007_g N_A1_M1004_g A1 A1 A1 N_A1_c_201_n
+ PM_SKY130_FD_SC_HVL__O21A_1%A1
x_PM_SKY130_FD_SC_HVL__O21A_1%X N_X_M1000_s N_X_M1002_s X X X X X X X
+ N_X_c_224_n N_X_c_227_n X PM_SKY130_FD_SC_HVL__O21A_1%X
x_PM_SKY130_FD_SC_HVL__O21A_1%VPWR N_VPWR_M1002_d N_VPWR_M1007_d VPWR
+ N_VPWR_c_243_n N_VPWR_c_246_n N_VPWR_c_249_n PM_SKY130_FD_SC_HVL__O21A_1%VPWR
x_PM_SKY130_FD_SC_HVL__O21A_1%VGND N_VGND_M1000_d N_VGND_M1003_d VGND
+ N_VGND_c_276_n N_VGND_c_278_n N_VGND_c_280_n PM_SKY130_FD_SC_HVL__O21A_1%VGND
x_PM_SKY130_FD_SC_HVL__O21A_1%A_460_107# N_A_460_107#_M1005_d
+ N_A_460_107#_M1004_d N_A_460_107#_c_306_n N_A_460_107#_c_308_n
+ N_A_460_107#_c_312_n N_A_460_107#_c_309_n
+ PM_SKY130_FD_SC_HVL__O21A_1%A_460_107#
cc_1 N_VNB_M1000_b N_A_83_87#_M1000_g 0.0637428f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=0.94
cc_2 N_VNB_c_2_p N_A_83_87#_M1000_g 6.11322e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=0.94
cc_3 N_VNB_M1000_b N_A_83_87#_c_70_n 0.014005f $X=-0.33 $Y=-0.265 $X2=1.495
+ $Y2=1.54
cc_4 N_VNB_M1000_b N_A_83_87#_c_71_n 0.0200377f $X=-0.33 $Y=-0.265 $X2=1.66
+ $Y2=0.66
cc_5 N_VNB_c_2_p N_A_83_87#_c_71_n 8.20017e-19 $X=0.24 $Y=0 $X2=1.66 $Y2=0.66
cc_6 N_VNB_M1000_b N_A_83_87#_c_73_n 0.00217795f $X=-0.33 $Y=-0.265 $X2=2.205
+ $Y2=1.54
cc_7 N_VNB_M1000_b N_A_83_87#_c_74_n 0.00155995f $X=-0.33 $Y=-0.265 $X2=2.29
+ $Y2=2.34
cc_8 N_VNB_M1000_b N_A_83_87#_c_75_n 0.0450076f $X=-0.33 $Y=-0.265 $X2=0.67
+ $Y2=1.63
cc_9 N_VNB_M1000_b N_A_83_87#_c_76_n 0.00148421f $X=-0.33 $Y=-0.265 $X2=1.66
+ $Y2=1.54
cc_10 N_VNB_M1000_b N_B1_M1005_g 0.0540153f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=1.585
cc_11 N_VNB_c_2_p N_B1_M1005_g 0.0023273f $X=0.24 $Y=0 $X2=0.665 $Y2=1.585
cc_12 N_VNB_M1000_b N_B1_c_129_n 0.0539776f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_13 N_VNB_M1000_b N_B1_c_130_n 0.0051395f $X=-0.33 $Y=-0.265 $X2=1.495
+ $Y2=1.54
cc_14 N_VNB_M1000_b N_A2_M1003_g 0.0439348f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=1.585
cc_15 N_VNB_c_2_p N_A2_M1003_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=1.585
cc_16 N_VNB_M1000_b N_A2_c_165_n 0.0438883f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_17 N_VNB_M1000_b N_A1_M1004_g 0.0496344f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=1.585
cc_18 N_VNB_c_2_p N_A1_M1004_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=1.585
cc_19 N_VNB_M1000_b A1 0.0268399f $X=-0.33 $Y=-0.265 $X2=0.9 $Y2=2.085
cc_20 N_VNB_M1000_b N_A1_c_201_n 0.0545489f $X=-0.33 $Y=-0.265 $X2=0.835
+ $Y2=1.54
cc_21 N_VNB_M1000_b N_X_c_224_n 0.0651504f $X=-0.33 $Y=-0.265 $X2=2.29 $Y2=2.34
cc_22 N_VNB_c_2_p N_X_c_224_n 5.68264e-19 $X=0.24 $Y=0 $X2=2.29 $Y2=2.34
cc_23 N_VNB_M1000_b N_VGND_c_276_n 0.0505892f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_24 N_VNB_c_2_p N_VGND_c_276_n 0.00216545f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_25 N_VNB_M1000_b N_VGND_c_278_n 0.0439761f $X=-0.33 $Y=-0.265 $X2=1.66
+ $Y2=1.455
cc_26 N_VNB_c_2_p N_VGND_c_278_n 0.00252795f $X=0.24 $Y=0 $X2=1.66 $Y2=1.455
cc_27 N_VNB_M1000_b N_VGND_c_280_n 0.0918564f $X=-0.33 $Y=-0.265 $X2=2.205
+ $Y2=1.54
cc_28 N_VNB_c_2_p N_VGND_c_280_n 0.462105f $X=0.24 $Y=0 $X2=2.205 $Y2=1.54
cc_29 N_VNB_M1000_b N_A_460_107#_c_306_n 0.01098f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=0.94
cc_30 N_VNB_c_2_p N_A_460_107#_c_306_n 8.71357e-19 $X=0.24 $Y=0 $X2=0.665
+ $Y2=0.94
cc_31 N_VNB_M1000_b N_A_460_107#_c_308_n 0.0120271f $X=-0.33 $Y=-0.265 $X2=0.9
+ $Y2=2.085
cc_32 N_VNB_M1000_b N_A_460_107#_c_309_n 0.031352f $X=-0.33 $Y=-0.265 $X2=1.495
+ $Y2=1.54
cc_33 N_VNB_c_2_p N_A_460_107#_c_309_n 8.20017e-19 $X=0.24 $Y=0 $X2=1.495
+ $Y2=1.54
cc_34 N_VPB_M1002_b N_A_83_87#_M1002_g 0.040851f $X=-0.33 $Y=1.885 $X2=0.9
+ $Y2=2.965
cc_35 VPB N_A_83_87#_M1002_g 0.00970178f $X=0 $Y=3.955 $X2=0.9 $Y2=2.965
cc_36 N_VPB_c_36_p N_A_83_87#_M1002_g 0.0152133f $X=4.08 $Y=4.07 $X2=0.9
+ $Y2=2.965
cc_37 N_VPB_M1002_b N_A_83_87#_c_74_n 0.00454551f $X=-0.33 $Y=1.885 $X2=2.29
+ $Y2=2.34
cc_38 VPB N_A_83_87#_c_74_n 5.14916e-19 $X=0 $Y=3.955 $X2=2.29 $Y2=2.34
cc_39 N_VPB_c_36_p N_A_83_87#_c_74_n 0.00887752f $X=4.08 $Y=4.07 $X2=2.29
+ $Y2=2.34
cc_40 N_VPB_M1002_b N_A_83_87#_c_75_n 0.0332142f $X=-0.33 $Y=1.885 $X2=0.67
+ $Y2=1.63
cc_41 N_VPB_M1002_b N_B1_M1006_g 0.0379899f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_42 VPB N_B1_M1006_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_43 N_VPB_c_36_p N_B1_M1006_g 0.0152133f $X=4.08 $Y=4.07 $X2=0 $Y2=0
cc_44 N_VPB_M1002_b N_B1_c_129_n 0.0256372f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_45 N_VPB_M1002_b N_B1_c_130_n 0.00593586f $X=-0.33 $Y=1.885 $X2=1.495
+ $Y2=1.54
cc_46 N_VPB_M1002_b N_A2_M1001_g 0.0513105f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_47 VPB N_A2_M1001_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_48 N_VPB_c_36_p N_A2_M1001_g 0.0191501f $X=4.08 $Y=4.07 $X2=0 $Y2=0
cc_49 N_VPB_M1002_b N_A2_c_165_n 0.00477027f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_50 N_VPB_M1002_b N_A1_M1007_g 0.0413428f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_51 VPB N_A1_M1007_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_52 N_VPB_c_36_p N_A1_M1007_g 0.0137101f $X=4.08 $Y=4.07 $X2=0 $Y2=0
cc_53 N_VPB_M1002_b N_A1_c_201_n 0.0295156f $X=-0.33 $Y=1.885 $X2=0.835 $Y2=1.54
cc_54 N_VPB_M1002_b N_X_c_224_n 0.00441854f $X=-0.33 $Y=1.885 $X2=2.29 $Y2=2.34
cc_55 N_VPB_M1002_b N_X_c_227_n 0.0679832f $X=-0.33 $Y=1.885 $X2=1.66 $Y2=1.54
cc_56 VPB N_X_c_227_n 0.00143441f $X=0 $Y=3.955 $X2=1.66 $Y2=1.54
cc_57 N_VPB_c_36_p N_X_c_227_n 0.0247302f $X=4.08 $Y=4.07 $X2=1.66 $Y2=1.54
cc_58 N_VPB_M1002_b X 0.0127472f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_59 N_VPB_M1002_b N_VPWR_c_243_n 0.00243985f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_243_n 0.00512219f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_61 N_VPB_c_36_p N_VPWR_c_243_n 0.0629871f $X=4.08 $Y=4.07 $X2=0 $Y2=0
cc_62 N_VPB_M1002_b N_VPWR_c_246_n 0.077399f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_246_n 0.00481441f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_64 N_VPB_c_36_p N_VPWR_c_246_n 0.0645871f $X=4.08 $Y=4.07 $X2=0 $Y2=0
cc_65 N_VPB_M1002_b N_VPWR_c_249_n 0.0467619f $X=-0.33 $Y=1.885 $X2=2.29
+ $Y2=3.59
cc_66 VPB N_VPWR_c_249_n 0.458533f $X=0 $Y=3.955 $X2=2.29 $Y2=3.59
cc_67 N_VPB_c_36_p N_VPWR_c_249_n 0.0195503f $X=4.08 $Y=4.07 $X2=2.29 $Y2=3.59
cc_68 N_A_83_87#_M1002_g N_B1_M1006_g 0.0181006f $X=0.9 $Y=2.965 $X2=0 $Y2=0
cc_69 N_A_83_87#_c_74_n N_B1_M1006_g 0.00406081f $X=2.29 $Y=2.34 $X2=0 $Y2=0
cc_70 N_A_83_87#_c_71_n N_B1_M1005_g 0.0318362f $X=1.66 $Y=0.66 $X2=0 $Y2=0
cc_71 N_A_83_87#_c_71_n N_B1_c_129_n 0.00595128f $X=1.66 $Y=0.66 $X2=0 $Y2=0
cc_72 N_A_83_87#_c_73_n N_B1_c_129_n 0.0397998f $X=2.205 $Y=1.54 $X2=0 $Y2=0
cc_73 N_A_83_87#_c_74_n N_B1_c_129_n 0.0198607f $X=2.29 $Y=2.34 $X2=0 $Y2=0
cc_74 N_A_83_87#_c_75_n N_B1_c_129_n 0.0181006f $X=0.67 $Y=1.63 $X2=0 $Y2=0
cc_75 N_A_83_87#_c_76_n N_B1_c_129_n 0.00937816f $X=1.66 $Y=1.54 $X2=0 $Y2=0
cc_76 N_A_83_87#_M1002_g N_B1_c_130_n 0.00244858f $X=0.9 $Y=2.965 $X2=0 $Y2=0
cc_77 N_A_83_87#_c_70_n N_B1_c_130_n 0.0305578f $X=1.495 $Y=1.54 $X2=0 $Y2=0
cc_78 N_A_83_87#_c_73_n N_B1_c_130_n 0.0118604f $X=2.205 $Y=1.54 $X2=0 $Y2=0
cc_79 N_A_83_87#_c_74_n N_B1_c_130_n 0.0206019f $X=2.29 $Y=2.34 $X2=0 $Y2=0
cc_80 N_A_83_87#_c_75_n N_B1_c_130_n 0.0189916f $X=0.67 $Y=1.63 $X2=0 $Y2=0
cc_81 N_A_83_87#_c_76_n N_B1_c_130_n 0.0263781f $X=1.66 $Y=1.54 $X2=0 $Y2=0
cc_82 N_A_83_87#_c_73_n A2 0.00591271f $X=2.205 $Y=1.54 $X2=0 $Y2=0
cc_83 N_A_83_87#_c_74_n A2 0.113069f $X=2.29 $Y=2.34 $X2=0 $Y2=0
cc_84 N_A_83_87#_c_73_n N_A2_c_165_n 0.00262132f $X=2.205 $Y=1.54 $X2=0 $Y2=0
cc_85 N_A_83_87#_c_74_n N_A2_c_165_n 0.0180363f $X=2.29 $Y=2.34 $X2=0 $Y2=0
cc_86 N_A_83_87#_c_73_n A1 0.00143297f $X=2.205 $Y=1.54 $X2=0.24 $Y2=0
cc_87 N_A_83_87#_M1000_g N_X_c_224_n 0.0287314f $X=0.665 $Y=0.94 $X2=2.16
+ $Y2=0.058
cc_88 N_A_83_87#_c_104_p N_X_c_224_n 0.0260417f $X=0.692 $Y=1.54 $X2=2.16
+ $Y2=0.058
cc_89 N_A_83_87#_M1002_g X 0.00915757f $X=0.9 $Y=2.965 $X2=0 $Y2=0
cc_90 N_A_83_87#_c_104_p X 0.00330106f $X=0.692 $Y=1.54 $X2=0 $Y2=0
cc_91 N_A_83_87#_c_75_n X 0.0190683f $X=0.67 $Y=1.63 $X2=0 $Y2=0
cc_92 N_A_83_87#_M1002_g N_VPWR_c_243_n 0.0758671f $X=0.9 $Y=2.965 $X2=0.24
+ $Y2=0
cc_93 N_A_83_87#_c_70_n N_VPWR_c_243_n 0.00598865f $X=1.495 $Y=1.54 $X2=0.24
+ $Y2=0
cc_94 N_A_83_87#_c_73_n N_VPWR_c_243_n 5.74911e-19 $X=2.205 $Y=1.54 $X2=0.24
+ $Y2=0
cc_95 N_A_83_87#_c_74_n N_VPWR_c_243_n 0.0612155f $X=2.29 $Y=2.34 $X2=0.24 $Y2=0
cc_96 N_A_83_87#_c_104_p N_VPWR_c_243_n 0.00190697f $X=0.692 $Y=1.54 $X2=0.24
+ $Y2=0
cc_97 N_A_83_87#_c_74_n N_VPWR_c_246_n 0.00951948f $X=2.29 $Y=2.34 $X2=0 $Y2=0
cc_98 N_A_83_87#_M1006_d N_VPWR_c_249_n 0.00788209f $X=2.15 $Y=2.215 $X2=0 $Y2=0
cc_99 N_A_83_87#_M1002_g N_VPWR_c_249_n 0.00885655f $X=0.9 $Y=2.965 $X2=0 $Y2=0
cc_100 N_A_83_87#_c_74_n N_VPWR_c_249_n 0.0269266f $X=2.29 $Y=2.34 $X2=0 $Y2=0
cc_101 N_A_83_87#_M1000_g N_VGND_c_276_n 0.0528502f $X=0.665 $Y=0.94 $X2=0.24
+ $Y2=0
cc_102 N_A_83_87#_c_70_n N_VGND_c_276_n 0.035177f $X=1.495 $Y=1.54 $X2=0.24
+ $Y2=0
cc_103 N_A_83_87#_c_71_n N_VGND_c_276_n 0.0639461f $X=1.66 $Y=0.66 $X2=0.24
+ $Y2=0
cc_104 N_A_83_87#_c_104_p N_VGND_c_276_n 0.0217256f $X=0.692 $Y=1.54 $X2=0.24
+ $Y2=0
cc_105 N_A_83_87#_c_75_n N_VGND_c_276_n 0.00120268f $X=0.67 $Y=1.63 $X2=0.24
+ $Y2=0
cc_106 N_A_83_87#_M1000_g N_VGND_c_280_n 0.00931089f $X=0.665 $Y=0.94 $X2=2.16
+ $Y2=0
cc_107 N_A_83_87#_c_71_n N_VGND_c_280_n 0.0325736f $X=1.66 $Y=0.66 $X2=2.16
+ $Y2=0
cc_108 N_A_83_87#_c_71_n N_A_460_107#_c_306_n 0.0187895f $X=1.66 $Y=0.66 $X2=0
+ $Y2=0
cc_109 N_A_83_87#_c_71_n N_A_460_107#_c_312_n 0.00614935f $X=1.66 $Y=0.66 $X2=0
+ $Y2=0
cc_110 N_A_83_87#_c_73_n N_A_460_107#_c_312_n 0.00613045f $X=2.205 $Y=1.54 $X2=0
+ $Y2=0
cc_111 N_B1_M1006_g N_A2_M1001_g 0.033882f $X=1.9 $Y=2.965 $X2=0 $Y2=0
cc_112 N_B1_M1005_g N_A2_M1003_g 0.0193985f $X=2.05 $Y=0.91 $X2=0 $Y2=0
cc_113 N_B1_c_129_n A2 5.36918e-19 $X=1.835 $Y=1.89 $X2=0 $Y2=0
cc_114 N_B1_c_129_n N_A2_c_165_n 0.0439826f $X=1.835 $Y=1.89 $X2=0 $Y2=0
cc_115 N_B1_c_130_n X 0.00509171f $X=1.835 $Y=1.89 $X2=0 $Y2=0
cc_116 N_B1_M1006_g N_VPWR_c_243_n 0.0959826f $X=1.9 $Y=2.965 $X2=0.24 $Y2=0
cc_117 N_B1_c_130_n N_VPWR_c_243_n 0.0680207f $X=1.835 $Y=1.89 $X2=0.24 $Y2=0
cc_118 N_B1_M1006_g N_VPWR_c_249_n 0.00818055f $X=1.9 $Y=2.965 $X2=0 $Y2=0
cc_119 N_B1_M1005_g N_VGND_c_276_n 0.00329258f $X=2.05 $Y=0.91 $X2=0.24 $Y2=0
cc_120 N_B1_M1005_g N_VGND_c_278_n 8.39127e-19 $X=2.05 $Y=0.91 $X2=4.08 $Y2=0
cc_121 N_B1_M1005_g N_VGND_c_280_n 0.0301625f $X=2.05 $Y=0.91 $X2=2.16 $Y2=0
cc_122 N_B1_M1005_g N_A_460_107#_c_306_n 0.0169926f $X=2.05 $Y=0.91 $X2=0 $Y2=0
cc_123 N_B1_M1005_g N_A_460_107#_c_312_n 0.00496761f $X=2.05 $Y=0.91 $X2=0 $Y2=0
cc_124 A2 N_A1_M1007_g 6.23726e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A2_M1003_g N_A1_M1004_g 0.030506f $X=2.83 $Y=0.91 $X2=0 $Y2=0
cc_126 A2 A1 0.0179584f $X=2.555 $Y=1.58 $X2=0.24 $Y2=0
cc_127 N_A2_c_165_n A1 0.0133003f $X=2.695 $Y=1.715 $X2=0.24 $Y2=0
cc_128 N_A2_M1001_g N_A1_c_201_n 0.0915444f $X=2.76 $Y=2.965 $X2=4.08 $Y2=0
cc_129 A2 N_A1_c_201_n 0.00171818f $X=2.555 $Y=1.58 $X2=4.08 $Y2=0
cc_130 N_A2_c_165_n N_A1_c_201_n 0.03502f $X=2.695 $Y=1.715 $X2=4.08 $Y2=0
cc_131 N_A2_M1001_g N_VPWR_c_246_n 0.0538731f $X=2.76 $Y=2.965 $X2=0 $Y2=0
cc_132 A2 N_VPWR_c_246_n 0.080245f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A2_c_165_n N_VPWR_c_246_n 0.00187389f $X=2.695 $Y=1.715 $X2=0 $Y2=0
cc_134 N_A2_M1001_g N_VPWR_c_249_n 0.0228802f $X=2.76 $Y=2.965 $X2=0 $Y2=0
cc_135 A2 N_VPWR_c_249_n 0.0110476f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A2_M1003_g N_VGND_c_278_n 0.0320804f $X=2.83 $Y=0.91 $X2=4.08 $Y2=0
cc_137 N_A2_M1003_g N_VGND_c_280_n 0.005327f $X=2.83 $Y=0.91 $X2=2.16 $Y2=0
cc_138 N_A2_M1003_g N_A_460_107#_c_306_n 0.0167032f $X=2.83 $Y=0.91 $X2=0 $Y2=0
cc_139 N_A2_M1003_g N_A_460_107#_c_308_n 0.0316632f $X=2.83 $Y=0.91 $X2=0.24
+ $Y2=0
cc_140 A2 N_A_460_107#_c_308_n 0.00924444f $X=2.555 $Y=1.58 $X2=0.24 $Y2=0
cc_141 N_A2_M1003_g N_A_460_107#_c_312_n 8.34821e-19 $X=2.83 $Y=0.91 $X2=0 $Y2=0
cc_142 A2 N_A_460_107#_c_312_n 0.00209616f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_143 N_A2_c_165_n N_A_460_107#_c_312_n 0.00207433f $X=2.695 $Y=1.715 $X2=0
+ $Y2=0
cc_144 N_A1_M1007_g N_VPWR_c_246_n 0.109371f $X=3.54 $Y=2.965 $X2=0 $Y2=0
cc_145 A1 N_VPWR_c_246_n 0.0598175f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_146 N_A1_c_201_n N_VPWR_c_246_n 0.00297548f $X=3.475 $Y=1.67 $X2=0 $Y2=0
cc_147 N_A1_M1007_g N_VPWR_c_249_n 0.00241703f $X=3.54 $Y=2.965 $X2=0 $Y2=0
cc_148 N_A1_M1004_g N_VGND_c_278_n 0.0323077f $X=3.63 $Y=0.91 $X2=4.08 $Y2=0
cc_149 N_A1_M1004_g N_VGND_c_280_n 0.00597233f $X=3.63 $Y=0.91 $X2=2.16 $Y2=0
cc_150 N_A1_M1004_g N_A_460_107#_c_308_n 0.0291399f $X=3.63 $Y=0.91 $X2=0.24
+ $Y2=0
cc_151 A1 N_A_460_107#_c_308_n 0.0737704f $X=3.995 $Y=1.58 $X2=0.24 $Y2=0
cc_152 N_A1_c_201_n N_A_460_107#_c_308_n 0.00234813f $X=3.475 $Y=1.67 $X2=0.24
+ $Y2=0
cc_153 N_A1_M1004_g N_A_460_107#_c_309_n 0.0179396f $X=3.63 $Y=0.91 $X2=0 $Y2=0
cc_154 N_X_c_227_n N_VPWR_c_243_n 0.0614045f $X=0.51 $Y=2.34 $X2=0.24 $Y2=0
cc_155 N_X_M1002_s N_VPWR_c_249_n 0.00221032f $X=0.365 $Y=2.215 $X2=0 $Y2=0
cc_156 N_X_c_227_n N_VPWR_c_249_n 0.0569588f $X=0.51 $Y=2.34 $X2=0 $Y2=0
cc_157 N_X_c_224_n N_VGND_c_276_n 0.0330164f $X=0.275 $Y=0.71 $X2=0.24 $Y2=0
cc_158 N_X_M1000_s N_VGND_c_280_n 0.00137624f $X=0.15 $Y=0.565 $X2=2.16 $Y2=0
cc_159 N_X_c_224_n N_VGND_c_280_n 0.0251405f $X=0.275 $Y=0.71 $X2=2.16 $Y2=0
cc_160 N_VGND_c_278_n N_A_460_107#_c_306_n 0.0307506f $X=2.87 $Y=0.48 $X2=0
+ $Y2=0
cc_161 N_VGND_c_280_n N_A_460_107#_c_306_n 0.0324443f $X=3.59 $Y=0.48 $X2=0
+ $Y2=0
cc_162 N_VGND_M1003_d N_A_460_107#_c_308_n 0.00414316f $X=3.08 $Y=0.535 $X2=0.24
+ $Y2=0
cc_163 N_VGND_c_278_n N_A_460_107#_c_308_n 0.0540633f $X=2.87 $Y=0.48 $X2=0.24
+ $Y2=0
cc_164 N_VGND_c_280_n N_A_460_107#_c_308_n 0.0141109f $X=3.59 $Y=0.48 $X2=0.24
+ $Y2=0
cc_165 N_VGND_c_278_n N_A_460_107#_c_309_n 0.0307506f $X=2.87 $Y=0.48 $X2=0
+ $Y2=0
cc_166 N_VGND_c_280_n N_A_460_107#_c_309_n 0.0332851f $X=3.59 $Y=0.48 $X2=0
+ $Y2=0
