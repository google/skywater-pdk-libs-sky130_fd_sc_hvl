* File: sky130_fd_sc_hvl__dfxtp_1.spice
* Created: Fri Aug 28 09:34:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__dfxtp_1.pex.spice"
.subckt sky130_fd_sc_hvl__dfxtp_1  VNB VPB CLK D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1022 N_VGND_M1022_d N_CLK_M1022_g N_A_30_127#_M1022_s N_VNB_M1022_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1004 N_A_339_559#_M1004_d N_A_30_127#_M1004_g N_VGND_M1022_d N_VNB_M1022_b NHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1016 N_A_605_563#_M1016_d N_D_M1016_g N_VGND_M1016_s N_VNB_M1022_b NHV L=0.5
+ W=0.42 AD=0.084 AS=0.1197 PD=0.82 PS=1.41 NRD=32.5698 NRS=0 M=1 R=0.84
+ SA=250000 SB=250007 A=0.21 P=1.84 MULT=1
MM1013 N_A_780_574#_M1013_d N_A_30_127#_M1013_g N_A_605_563#_M1016_d
+ N_VNB_M1022_b NHV L=0.5 W=0.42 AD=0.09975 AS=0.084 PD=0.895 PS=0.82
+ NRD=37.9962 NRS=0 M=1 R=0.84 SA=250001 SB=250006 A=0.21 P=1.84 MULT=1
MM1005 A_1015_113# N_A_339_559#_M1005_g N_A_780_574#_M1013_d N_VNB_M1022_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.09975 PD=0.63 PS=0.895 NRD=13.566 NRS=14.9226 M=1
+ R=0.84 SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1007 N_VGND_M1007_d N_A_1024_371#_M1007_g A_1015_113# N_VNB_M1022_b NHV L=0.5
+ W=0.42 AD=0.114854 AS=0.0441 PD=0.879487 PS=0.63 NRD=31.2132 NRS=13.566 M=1
+ R=0.84 SA=250003 SB=250004 A=0.21 P=1.84 MULT=1
MM1021 N_A_1024_371#_M1021_d N_A_780_574#_M1021_g N_VGND_M1007_d N_VNB_M1022_b
+ NHV L=0.5 W=0.75 AD=0.166635 AS=0.205096 PD=1.46795 PS=1.57051 NRD=0
+ NRS=12.1524 M=1 R=1.5 SA=250002 SB=250002 A=0.375 P=2.5 MULT=1
MM1010 N_A_1455_543#_M1010_d N_A_339_559#_M1010_g N_A_1024_371#_M1021_d
+ N_VNB_M1022_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.0933154 PD=0.7 PS=0.822051 NRD=0
+ NRS=31.2132 M=1 R=0.84 SA=250004 SB=250003 A=0.21 P=1.84 MULT=1
MM1002 A_1687_113# N_A_30_127#_M1002_g N_A_1455_543#_M1010_d N_VNB_M1022_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250005 SB=250002 A=0.21 P=1.84 MULT=1
MM1008 N_VGND_M1008_d N_A_1729_87#_M1008_g A_1687_113# N_VNB_M1022_b NHV L=0.5
+ W=0.42 AD=0.115823 AS=0.0441 PD=0.940513 PS=0.63 NRD=75.9924 NRS=13.566 M=1
+ R=0.84 SA=250006 SB=250001 A=0.21 P=1.84 MULT=1
MM1019 N_A_1729_87#_M1019_d N_A_1455_543#_M1019_g N_VGND_M1008_d N_VNB_M1022_b
+ NHV L=0.5 W=0.75 AD=0.21375 AS=0.206827 PD=2.07 PS=1.67949 NRD=0 NRS=0 M=1
+ R=1.5 SA=250004 SB=250000 A=0.375 P=2.5 MULT=1
MM1023 N_Q_M1023_d N_A_1729_87#_M1023_g N_VGND_M1023_s N_VNB_M1022_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.21375 PD=2.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1011 N_VPWR_M1011_d N_CLK_M1011_g N_A_30_127#_M1011_s N_VPB_M1011_b PHV L=0.5
+ W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1001 N_A_339_559#_M1001_d N_A_30_127#_M1001_g N_VPWR_M1011_d N_VPB_M1011_b PHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1017 N_A_605_563#_M1017_d N_D_M1017_g N_VPWR_M1017_s N_VPB_M1011_b PHV L=0.5
+ W=0.42 AD=0.0826 AS=0.1113 PD=0.85 PS=1.37 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250005 A=0.21 P=1.84 MULT=1
MM1012 N_A_780_574#_M1012_d N_A_339_559#_M1012_g N_A_605_563#_M1017_d
+ N_VPB_M1011_b PHV L=0.5 W=0.42 AD=0.129575 AS=0.0826 PD=1.085 PS=0.85
+ NRD=84.1164 NRS=43.1851 M=1 R=0.84 SA=250001 SB=250004 A=0.21 P=1.84 MULT=1
MM1000 A_982_543# N_A_30_127#_M1000_g N_A_780_574#_M1012_d N_VPB_M1011_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.129575 PD=0.63 PS=1.085 NRD=22.729 NRS=22.729 M=1
+ R=0.84 SA=250001 SB=250005 A=0.21 P=1.84 MULT=1
MM1006 N_VPWR_M1006_d N_A_1024_371#_M1006_g A_982_543# N_VPB_M1011_b PHV L=0.5
+ W=0.42 AD=0.0920451 AS=0.0441 PD=0.81338 PS=0.63 NRD=74.6428 NRS=22.729 M=1
+ R=0.84 SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1003 N_A_1024_371#_M1003_d N_A_780_574#_M1003_g N_VPWR_M1006_d N_VPB_M1011_b
+ PHV L=0.5 W=1 AD=0.14 AS=0.219155 PD=1.28 PS=1.93662 NRD=0 NRS=0 M=1 R=2
+ SA=250001 SB=250002 A=0.5 P=3 MULT=1
MM1020 N_A_1455_543#_M1020_d N_A_30_127#_M1020_g N_A_1024_371#_M1003_d
+ N_VPB_M1011_b PHV L=0.5 W=1 AD=0.574789 AS=0.14 PD=2.64789 PS=1.28 NRD=96.4359
+ NRS=0 M=1 R=2 SA=250002 SB=250002 A=0.5 P=3 MULT=1
MM1014 A_1731_543# N_A_339_559#_M1014_g N_A_1455_543#_M1020_d N_VPB_M1011_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.241411 PD=0.63 PS=1.11211 NRD=22.729 NRS=43.1851
+ M=1 R=0.84 SA=250005 SB=250002 A=0.21 P=1.84 MULT=1
MM1015 N_VPWR_M1015_d N_A_1729_87#_M1015_g A_1731_543# N_VPB_M1011_b PHV L=0.5
+ W=0.42 AD=0.0920451 AS=0.0441 PD=0.81338 PS=0.63 NRD=43.1851 NRS=22.729 M=1
+ R=0.84 SA=250006 SB=250001 A=0.21 P=1.84 MULT=1
MM1018 N_A_1729_87#_M1018_d N_A_1455_543#_M1018_g N_VPWR_M1015_d N_VPB_M1011_b
+ PHV L=0.5 W=1 AD=0.265 AS=0.219155 PD=2.53 PS=1.93662 NRD=0 NRS=0 M=1 R=2
+ SA=250003 SB=250000 A=0.5 P=3 MULT=1
MM1009 N_Q_M1009_d N_A_1729_87#_M1009_g N_VPWR_M1009_s N_VPB_M1011_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.3975 PD=3.53 PS=3.53 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
DX24_noxref N_VNB_M1022_b N_VPB_M1011_b NWDIODE A=32.916 P=30.52
*
.include "sky130_fd_sc_hvl__dfxtp_1.pxi.spice"
*
.ends
*
*
