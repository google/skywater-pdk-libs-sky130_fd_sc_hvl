# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
SITE unithvdbl
  SYMMETRY y ;
  CLASS CORE ;
  SIZE  8.640000 BY  8.140000 ;
END unithvdbl
MACRO sky130_fd_sc_hvl__lsbufhv2hv_hl_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__lsbufhv2hv_hl_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  8.140000 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355000 1.775000 4.685000 2.900000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.995000 0.495000 3.395000 4.065000 ;
    END
  END X
  PIN LOWHVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 8.570000 3.305000 ;
    END
  END LOWHVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 8.640000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 8.640000 8.255000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 8.640000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 8.640000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.985000 0.800000 4.155000 ;
      RECT 0.000000  8.055000 8.640000 8.225000 ;
      RECT 3.130000  4.265000 5.095000 4.835000 ;
      RECT 3.565000  0.365000 4.515000 1.265000 ;
      RECT 3.565000  1.435000 5.115000 1.605000 ;
      RECT 3.565000  1.605000 3.895000 2.065000 ;
      RECT 3.565000  2.485000 4.185000 4.265000 ;
      RECT 4.865000  0.495000 5.115000 1.435000 ;
      RECT 4.865000  1.605000 5.115000 3.315000 ;
      RECT 7.425000  3.985000 8.640000 4.155000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.155000  8.055000 0.325000 8.225000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  8.055000 0.805000 8.225000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  8.055000 1.285000 8.225000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  8.055000 1.765000 8.225000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  8.055000 2.245000 8.225000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  8.055000 2.725000 8.225000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  8.055000 3.205000 8.225000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  8.055000 3.685000 8.225000 ;
      RECT 3.595000  0.395000 3.765000 0.565000 ;
      RECT 3.630000  3.075000 3.800000 3.245000 ;
      RECT 3.955000  0.395000 4.125000 0.565000 ;
      RECT 3.990000  3.075000 4.160000 3.245000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  8.055000 4.165000 8.225000 ;
      RECT 4.315000  0.395000 4.485000 0.565000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  8.055000 4.645000 8.225000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  8.055000 5.125000 8.225000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  8.055000 5.605000 8.225000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  8.055000 6.085000 8.225000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  8.055000 6.565000 8.225000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  8.055000 7.045000 8.225000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  8.055000 7.525000 8.225000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 7.835000  8.055000 8.005000 8.225000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.985000 8.485000 4.155000 ;
      RECT 8.315000  8.055000 8.485000 8.225000 ;
    LAYER met1 ;
      RECT 0.000000 -0.115000 8.640000 0.115000 ;
      RECT 0.000000  0.255000 8.640000 0.625000 ;
      RECT 0.000000  3.445000 8.640000 3.815000 ;
  END
END sky130_fd_sc_hvl__lsbufhv2hv_hl_1
END LIBRARY
