* File: sky130_fd_sc_hvl__and3_1.spice
* Created: Wed Sep  2 09:03:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__and3_1.pex.spice"
.subckt sky130_fd_sc_hvl__and3_1  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 A_201_173# N_A_M1002_g N_A_30_517#_M1002_s N_VNB_M1002_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.1302 PD=0.63 PS=1.46 NRD=13.566 NRS=6.783 M=1 R=0.84 SA=250000
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1003 A_343_173# N_B_M1003_g A_201_173# N_VNB_M1002_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=13.566 NRS=13.566 M=1 R=0.84 SA=250001
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1004 N_VGND_M1004_d N_C_M1004_g A_343_173# N_VNB_M1002_b NHV L=0.5 W=0.42
+ AD=0.109146 AS=0.0441 PD=0.897436 PS=0.63 NRD=59.7132 NRS=13.566 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1001 N_X_M1001_d N_A_30_517#_M1001_g N_VGND_M1004_d N_VNB_M1002_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.194904 PD=2.03 PS=1.60256 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_30_517#_M1007_s N_VPB_M1007_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1000 N_A_30_517#_M1000_d N_B_M1000_g N_VPWR_M1007_d N_VPB_M1007_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250001
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1006 N_VPWR_M1006_d N_C_M1006_g N_A_30_517#_M1000_d N_VPB_M1007_b PHV L=0.5
+ W=0.42 AD=0.103622 AS=0.0588 PD=0.829062 PS=0.7 NRD=52.2958 NRS=0 M=1 R=0.84
+ SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1005 N_X_M1005_d N_A_30_517#_M1005_g N_VPWR_M1006_d N_VPB_M1007_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.370078 PD=3.57 PS=2.96094 NRD=0 NRS=0 M=1 R=3 SA=250001
+ SB=250000 A=0.75 P=4 MULT=1
DX8_noxref N_VNB_M1002_b N_VPB_M1007_b NWDIODE A=11.7 P=14.2
*
.include "sky130_fd_sc_hvl__and3_1.pxi.spice"
*
.ends
*
*
