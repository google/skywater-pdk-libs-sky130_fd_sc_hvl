* File: sky130_fd_sc_hvl__dlxtp_1.spice
* Created: Wed Sep  2 09:06:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__dlxtp_1.pex.spice"
.subckt sky130_fd_sc_hvl__dlxtp_1  VNB VPB GATE D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_GATE_M1010_g N_A_30_443#_M1010_s N_VNB_M1010_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1000 N_A_384_107#_M1000_d N_A_30_443#_M1000_g N_VGND_M1010_d N_VNB_M1010_b NHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1004 N_A_650_107#_M1004_d N_D_M1004_g N_VGND_M1004_s N_VNB_M1010_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1015 N_A_806_107#_M1015_d N_A_384_107#_M1015_g N_A_650_107#_M1004_d
+ N_VNB_M1010_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0
+ M=1 R=0.84 SA=250001 SB=250002 A=0.21 P=1.84 MULT=1
MM1007 A_962_107# N_A_30_443#_M1007_g N_A_806_107#_M1015_d N_VNB_M1010_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1012 N_VGND_M1012_d N_A_1004_81#_M1012_g A_962_107# N_VNB_M1010_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1003 N_VGND_M1003_d N_A_806_107#_M1003_g N_A_1004_81#_M1003_s N_VNB_M1010_b
+ NHV L=0.5 W=0.42 AD=0.0933154 AS=0.1113 PD=0.822051 PS=1.37 NRD=31.2132 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1009 N_Q_M1009_d N_A_806_107#_M1009_g N_VGND_M1003_d N_VNB_M1010_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.166635 PD=2.03 PS=1.46795 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_GATE_M1005_g N_A_30_443#_M1005_s N_VPB_M1005_b PHV L=0.5
+ W=0.75 AD=0.21375 AS=0.19875 PD=1.32 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1011 N_A_384_107#_M1011_d N_A_30_443#_M1011_g N_VPWR_M1005_d N_VPB_M1005_b PHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.21375 PD=2.03 PS=1.32 NRD=0 NRS=73.8406 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1013 N_A_650_107#_M1013_d N_D_M1013_g N_VPWR_M1013_s N_VPB_M1005_b PHV L=0.5
+ W=0.75 AD=0.133125 AS=0.2025 PD=1.105 PS=2.04 NRD=19.0809 NRS=1.2606 M=1 R=1.5
+ SA=250000 SB=250002 A=0.375 P=2.5 MULT=1
MM1006 N_A_806_107#_M1006_d N_A_30_443#_M1006_g N_A_650_107#_M1013_d
+ N_VPB_M1005_b PHV L=0.5 W=0.75 AD=0.166635 AS=0.133125 PD=1.46795 PS=1.105
+ NRD=0 NRS=0 M=1 R=1.5 SA=250001 SB=250001 A=0.375 P=2.5 MULT=1
MM1014 A_1014_587# N_A_384_107#_M1014_g N_A_806_107#_M1006_d N_VPB_M1005_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0933154 PD=0.63 PS=0.822051 NRD=22.729 NRS=52.2958
+ M=1 R=0.84 SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1001 N_VPWR_M1001_d N_A_1004_81#_M1001_g A_1014_587# N_VPB_M1005_b PHV L=0.5
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1008 N_VPWR_M1008_d N_A_806_107#_M1008_g N_A_1004_81#_M1008_s N_VPB_M1005_b
+ PHV L=0.5 W=0.42 AD=0.103622 AS=0.1197 PD=0.829062 PS=1.41 NRD=54.5687 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1002 N_Q_M1002_d N_A_806_107#_M1002_g N_VPWR_M1008_d N_VPB_M1005_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.370078 PD=3.57 PS=2.96094 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
DX16_noxref N_VNB_M1010_b N_VPB_M1005_b NWDIODE A=22.932 P=22.84
*
.include "sky130_fd_sc_hvl__dlxtp_1.pxi.spice"
*
.ends
*
*
