* File: sky130_fd_sc_hvl__lsbuflv2hv_1.pxi.spice
* Created: Wed Sep  2 09:07:42 2020
* 
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%VNB N_VNB_M1014_b VNB VNB N_VNB_c_25_p
+ N_VNB_c_15_p VNB VNB PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%VNB
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%VPB N_VPB_X20_noxref_D1 N_VPB_M1018_b VPB
+ N_VPB_c_91_n N_VPB_c_101_p N_VPB_c_92_n VPB
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%VPB
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%LVPWR N_LVPWR_M1004_d N_LVPWR_M1004_b
+ N_LVPWR_c_167_p LVPWR N_LVPWR_c_164_n LVPWR
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%LVPWR
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A N_A_c_215_n N_A_c_216_n N_A_M1014_g
+ N_A_M1004_g N_A_c_217_n A A N_A_c_219_n PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_404_1133# N_A_404_1133#_M1014_s
+ N_A_404_1133#_M1004_s N_A_404_1133#_c_247_n N_A_404_1133#_M1002_g
+ N_A_404_1133#_c_248_n N_A_404_1133#_M1003_g N_A_404_1133#_c_249_n
+ N_A_404_1133#_M1008_g N_A_404_1133#_c_250_n N_A_404_1133#_M1015_g
+ N_A_404_1133#_M1017_g N_A_404_1133#_c_251_n N_A_404_1133#_M1010_g
+ N_A_404_1133#_c_252_n N_A_404_1133#_M1011_g N_A_404_1133#_c_254_n
+ N_A_404_1133#_c_255_n N_A_404_1133#_c_256_n N_A_404_1133#_c_257_n
+ N_A_404_1133#_c_272_n N_A_404_1133#_c_258_n N_A_404_1133#_c_259_n
+ N_A_404_1133#_c_276_n N_A_404_1133#_c_292_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_404_1133#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_1197_107# N_A_1197_107#_M1000_d
+ N_A_1197_107#_M1009_d N_A_1197_107#_M1019_d N_A_1197_107#_M1018_s
+ N_A_1197_107#_c_372_p N_A_1197_107#_c_365_n N_A_1197_107#_c_350_n
+ N_A_1197_107#_c_354_n N_A_1197_107#_c_355_n N_A_1197_107#_c_356_n
+ N_A_1197_107#_c_374_p N_A_1197_107#_c_351_n N_A_1197_107#_c_369_n
+ N_A_1197_107#_c_352_n N_A_1197_107#_c_360_n N_A_1197_107#_c_362_n
+ N_A_1197_107#_M1006_g PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_1197_107#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_772_151# N_A_772_151#_M1015_d
+ N_A_772_151#_M1017_d N_A_772_151#_c_426_n N_A_772_151#_M1000_g
+ N_A_772_151#_c_427_n N_A_772_151#_M1007_g N_A_772_151#_c_428_n
+ N_A_772_151#_M1009_g N_A_772_151#_c_429_n N_A_772_151#_M1012_g
+ N_A_772_151#_c_430_n N_A_772_151#_M1019_g N_A_772_151#_c_432_n
+ N_A_772_151#_c_433_n N_A_772_151#_c_434_n N_A_772_151#_c_443_n
+ N_A_772_151#_c_435_n N_A_772_151#_c_444_n N_A_772_151#_c_436_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_772_151#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_504_1221# N_A_504_1221#_M1002_s
+ N_A_504_1221#_M1008_s N_A_504_1221#_M1011_s N_A_504_1221#_M1006_s
+ N_A_504_1221#_c_504_n N_A_504_1221#_c_517_n N_A_504_1221#_M1013_g
+ N_A_504_1221#_c_505_n N_A_504_1221#_M1016_g N_A_504_1221#_M1018_g
+ N_A_504_1221#_c_521_n N_A_504_1221#_c_537_n N_A_504_1221#_c_539_n
+ N_A_504_1221#_c_507_n N_A_504_1221#_c_542_n N_A_504_1221#_c_544_n
+ N_A_504_1221#_c_508_n N_A_504_1221#_c_510_n N_A_504_1221#_c_526_n
+ N_A_504_1221#_c_511_n N_A_504_1221#_c_528_n N_A_504_1221#_c_572_p
+ N_A_504_1221#_c_529_n N_A_504_1221#_c_512_n N_A_504_1221#_c_513_n
+ N_A_504_1221#_c_514_n N_A_504_1221#_c_532_n N_A_504_1221#_c_515_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_504_1221#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_1711_885# N_A_1711_885#_M1016_s
+ N_A_1711_885#_M1013_s N_A_1711_885#_M1001_g N_A_1711_885#_M1005_g
+ N_A_1711_885#_c_616_n N_A_1711_885#_c_609_n N_A_1711_885#_c_611_n
+ N_A_1711_885#_c_612_n N_A_1711_885#_c_634_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%A_1711_885#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%VPWR N_VPWR_M1018_d N_VPWR_M1006_d
+ N_VPWR_M1013_d VPWR VPWR N_VPWR_c_657_n N_VPWR_c_660_n N_VPWR_c_655_n
+ N_VPWR_c_668_n N_VPWR_c_656_n VPWR VPWR PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%VPWR
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%X N_X_M1005_d N_X_M1001_d X X X X X
+ N_X_c_725_n X X PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%X
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%VGND N_VGND_M1002_d N_VGND_M1003_d
+ N_VGND_M1014_d N_VGND_M1010_d N_VGND_M1000_s N_VGND_M1007_s N_VGND_M1012_s
+ N_VGND_M1016_d N_VGND_c_738_n N_VGND_c_740_n N_VGND_c_742_n N_VGND_c_743_n
+ N_VGND_c_745_n N_VGND_c_747_n N_VGND_c_749_n N_VGND_c_751_n N_VGND_c_753_n
+ VGND VGND N_VGND_c_755_n N_VGND_c_756_n N_VGND_c_787_n N_VGND_c_758_n
+ N_VGND_c_793_n N_VGND_c_760_n N_VGND_c_806_n N_VGND_c_809_n N_VGND_c_761_n
+ N_VGND_c_763_n N_VGND_c_765_n N_VGND_c_767_n VGND VGND
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_1%VGND
cc_1 N_VNB_M1014_b N_VPB_c_91_n 0.0021751f $X=-0.33 $Y=-0.265 $X2=0.24 $Y2=4.07
cc_2 N_VNB_M1014_b N_VPB_c_92_n 0.079871f $X=-0.33 $Y=-0.265 $X2=10.32 $Y2=4.07
cc_3 N_VNB_M1014_b LVPWR 0.156699f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_4 N_VNB_M1014_b N_A_c_215_n 0.0315583f $X=-0.33 $Y=-0.265 $X2=0 $Y2=3.985
cc_5 N_VNB_M1014_b N_A_c_216_n 0.0215558f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_M1014_b N_A_c_217_n 0.00851298f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_7 N_VNB_M1014_b A 0.0248803f $X=-0.33 $Y=-0.265 $X2=0 $Y2=3.955
cc_8 N_VNB_M1014_b N_A_c_219_n 0.0812462f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_M1014_b N_A_404_1133#_c_247_n 0.0411781f $X=-0.33 $Y=-0.265 $X2=-0.33
+ $Y2=1.885
cc_10 N_VNB_M1014_b N_A_404_1133#_c_248_n 0.0358616f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1014_b N_A_404_1133#_c_249_n 0.0358616f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1014_b N_A_404_1133#_c_250_n 0.0223696f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1014_b N_A_404_1133#_c_251_n 0.0358616f $X=-0.33 $Y=-0.265 $X2=7.92
+ $Y2=4.07
cc_14 N_VNB_M1014_b N_A_404_1133#_c_252_n 0.376504f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_15 N_VNB_c_15_p N_A_404_1133#_c_252_n 0.00160584f $X=10.32 $Y=8.14 $X2=10.32
+ $Y2=4.07
cc_16 N_VNB_M1014_b N_A_404_1133#_c_254_n 0.0125974f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_17 N_VNB_M1014_b N_A_404_1133#_c_255_n 0.00411489f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1014_b N_A_404_1133#_c_256_n 0.164089f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_19 N_VNB_M1014_b N_A_404_1133#_c_257_n 0.035967f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_20 N_VNB_M1014_b N_A_404_1133#_c_258_n 0.00652689f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_21 N_VNB_M1014_b N_A_404_1133#_c_259_n 0.0344484f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_22 N_VNB_M1014_b N_A_1197_107#_c_350_n 0.00599753f $X=-0.33 $Y=-0.265
+ $X2=7.92 $Y2=4.07
cc_23 N_VNB_M1014_b N_A_1197_107#_c_351_n 0.0145123f $X=-0.33 $Y=-0.265
+ $X2=10.32 $Y2=4.07
cc_24 N_VNB_M1014_b N_A_1197_107#_c_352_n 0.0715552f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_25 N_VNB_c_25_p N_A_1197_107#_c_352_n 7.98897e-19 $X=10.32 $Y=0 $X2=0 $Y2=0
cc_26 N_VNB_M1014_b N_A_772_151#_c_426_n 0.0398058f $X=-0.33 $Y=-0.265 $X2=-0.33
+ $Y2=1.885
cc_27 N_VNB_M1014_b N_A_772_151#_c_427_n 0.0358616f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_28 N_VNB_M1014_b N_A_772_151#_c_428_n 0.0358616f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_29 N_VNB_M1014_b N_A_772_151#_c_429_n 0.0358616f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_30 N_VNB_M1014_b N_A_772_151#_c_430_n 0.222739f $X=-0.33 $Y=-0.265 $X2=7.92
+ $Y2=4.07
cc_31 N_VNB_c_25_p N_A_772_151#_c_430_n 0.00160584f $X=10.32 $Y=0 $X2=7.92
+ $Y2=4.07
cc_32 N_VNB_M1014_b N_A_772_151#_c_432_n 0.0244016f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_33 N_VNB_M1014_b N_A_772_151#_c_433_n 0.0185531f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_34 N_VNB_M1014_b N_A_772_151#_c_434_n 0.014445f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_35 N_VNB_M1014_b N_A_772_151#_c_435_n 0.0384012f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_36 N_VNB_M1014_b N_A_772_151#_c_436_n 0.084631f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_37 N_VNB_M1014_b N_A_504_1221#_c_504_n 0.0621692f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_38 N_VNB_M1014_b N_A_504_1221#_c_505_n 0.0873403f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_39 N_VNB_c_15_p N_A_504_1221#_c_505_n 0.00181995f $X=10.32 $Y=8.14 $X2=0
+ $Y2=0
cc_40 N_VNB_M1014_b N_A_504_1221#_c_507_n 0.0134401f $X=-0.33 $Y=-0.265
+ $X2=10.32 $Y2=4.07
cc_41 N_VNB_M1014_b N_A_504_1221#_c_508_n 0.072465f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_42 N_VNB_c_15_p N_A_504_1221#_c_508_n 7.98897e-19 $X=10.32 $Y=8.14 $X2=0
+ $Y2=0
cc_43 N_VNB_M1014_b N_A_504_1221#_c_510_n 0.071364f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_44 N_VNB_M1014_b N_A_504_1221#_c_511_n 0.0424618f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_45 N_VNB_M1014_b N_A_504_1221#_c_512_n 0.0133586f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_M1014_b N_A_504_1221#_c_513_n 0.0134401f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_47 N_VNB_M1014_b N_A_504_1221#_c_514_n 0.0113458f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_M1014_b N_A_504_1221#_c_515_n 0.036449f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_49 N_VNB_M1014_b N_A_1711_885#_M1005_g 0.0682348f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_c_15_p N_A_1711_885#_M1005_g 0.00161049f $X=10.32 $Y=8.14 $X2=0
+ $Y2=0
cc_51 N_VNB_M1014_b N_A_1711_885#_c_609_n 0.0496534f $X=-0.33 $Y=-0.265 $X2=7.92
+ $Y2=4.07
cc_52 N_VNB_c_15_p N_A_1711_885#_c_609_n 7.98897e-19 $X=10.32 $Y=8.14 $X2=7.92
+ $Y2=4.07
cc_53 N_VNB_M1014_b N_A_1711_885#_c_611_n 0.00203039f $X=-0.33 $Y=-0.265
+ $X2=10.32 $Y2=4.07
cc_54 N_VNB_M1014_b N_A_1711_885#_c_612_n 0.0377119f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_55 N_VNB_M1014_b N_VPWR_c_655_n 0.0939361f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_56 N_VNB_M1014_b N_VPWR_c_656_n 0.271949f $X=-0.33 $Y=-0.265 $X2=4.8
+ $Y2=4.068
cc_57 N_VNB_M1014_b X 0.0443485f $X=-0.33 $Y=-0.265 $X2=0 $Y2=3.955
cc_58 N_VNB_c_15_p X 7.98897e-19 $X=10.32 $Y=8.14 $X2=0 $Y2=3.955
cc_59 N_VNB_M1014_b X 0.0234434f $X=-0.33 $Y=-0.265 $X2=4.8 $Y2=4.07
cc_60 N_VNB_M1014_b N_VGND_c_738_n 0.0718145f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_61 N_VNB_c_15_p N_VGND_c_738_n 0.00332742f $X=10.32 $Y=8.14 $X2=10.32
+ $Y2=4.07
cc_62 N_VNB_M1014_b N_VGND_c_740_n 0.0481389f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_63 N_VNB_c_15_p N_VGND_c_740_n 0.00198821f $X=10.32 $Y=8.14 $X2=10.32
+ $Y2=4.07
cc_64 N_VNB_M1014_b N_VGND_c_742_n 0.00570671f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_65 N_VNB_M1014_b N_VGND_c_743_n 0.118091f $X=-0.33 $Y=-0.265 $X2=4.8 $Y2=4.07
cc_66 N_VNB_c_15_p N_VGND_c_743_n 0.00531562f $X=10.32 $Y=8.14 $X2=4.8 $Y2=4.07
cc_67 N_VNB_M1014_b N_VGND_c_745_n 0.0718145f $X=-0.33 $Y=-0.265 $X2=5.28
+ $Y2=4.07
cc_68 N_VNB_c_25_p N_VGND_c_745_n 0.00332742f $X=10.32 $Y=0 $X2=5.28 $Y2=4.07
cc_69 N_VNB_M1014_b N_VGND_c_747_n 0.0481389f $X=-0.33 $Y=-0.265 $X2=7.92
+ $Y2=4.07
cc_70 N_VNB_c_25_p N_VGND_c_747_n 0.00198821f $X=10.32 $Y=0 $X2=7.92 $Y2=4.07
cc_71 N_VNB_M1014_b N_VGND_c_749_n 0.118091f $X=-0.33 $Y=-0.265 $X2=10.32
+ $Y2=4.07
cc_72 N_VNB_c_25_p N_VGND_c_749_n 0.00531562f $X=10.32 $Y=0 $X2=10.32 $Y2=4.07
cc_73 N_VNB_M1014_b N_VGND_c_751_n 0.0443345f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_74 N_VNB_c_15_p N_VGND_c_751_n 0.00198821f $X=10.32 $Y=8.14 $X2=0 $Y2=0
cc_75 N_VNB_M1014_b N_VGND_c_753_n 0.0443345f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_76 N_VNB_c_25_p N_VGND_c_753_n 0.00198821f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_77 N_VNB_M1014_b N_VGND_c_755_n 0.088056f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_78 N_VNB_M1014_b N_VGND_c_756_n 0.0262752f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_79 N_VNB_c_25_p N_VGND_c_756_n 0.00102546f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_80 N_VNB_M1014_b N_VGND_c_758_n 0.0262752f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_81 N_VNB_c_25_p N_VGND_c_758_n 0.00102546f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_82 N_VNB_M1014_b N_VGND_c_760_n 0.0461766f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_83 N_VNB_M1014_b N_VGND_c_761_n 0.369793f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_84 N_VNB_c_25_p N_VGND_c_761_n 1.11823f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_85 N_VNB_M1014_b N_VGND_c_763_n 0.0294115f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_86 N_VNB_c_15_p N_VGND_c_763_n 0.00159492f $X=10.32 $Y=8.14 $X2=0 $Y2=0
cc_87 N_VNB_M1014_b N_VGND_c_765_n 0.328524f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_88 N_VNB_c_15_p N_VGND_c_765_n 1.11834f $X=10.32 $Y=8.14 $X2=0 $Y2=0
cc_89 N_VNB_M1014_b N_VGND_c_767_n 0.0167066f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_90 N_VNB_c_25_p N_VGND_c_767_n 8.02293e-19 $X=10.32 $Y=0 $X2=0 $Y2=0
cc_91 N_VPB_c_92_n N_LVPWR_M1004_b 0.00792118f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_92 N_VPB_X20_noxref_D1 LVPWR 0.050189f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_93 N_VPB_M1018_b LVPWR 0.0937645f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_94 N_VPB_c_92_n N_LVPWR_c_164_n 0.0433246f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_95 N_VPB_c_92_n N_A_404_1133#_c_255_n 0.0252548f $X=10.32 $Y=4.07 $X2=4.8
+ $Y2=0.058
cc_96 N_VPB_c_92_n N_A_1197_107#_c_354_n 0.00396985f $X=10.32 $Y=4.07 $X2=0
+ $Y2=0
cc_97 N_VPB_M1018_b N_A_1197_107#_c_355_n 0.0156528f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_98 N_VPB_M1018_b N_A_1197_107#_c_356_n 0.020028f $X=6.335 $Y=2.465 $X2=0.24
+ $Y2=8.14
cc_99 N_VPB_c_101_p N_A_1197_107#_c_356_n 0.00784462f $X=10.32 $Y=4.07 $X2=0.24
+ $Y2=8.14
cc_100 N_VPB_c_92_n N_A_1197_107#_c_356_n 0.0270266f $X=10.32 $Y=4.07 $X2=0.24
+ $Y2=8.14
cc_101 N_VPB_M1018_b N_A_1197_107#_c_351_n 0.00689188f $X=6.335 $Y=2.465
+ $X2=10.32 $Y2=8.14
cc_102 N_VPB_M1018_b N_A_1197_107#_c_360_n 0.135402f $X=6.335 $Y=2.465 $X2=4.8
+ $Y2=8.14
cc_103 N_VPB_c_101_p N_A_1197_107#_c_360_n 0.0038941f $X=10.32 $Y=4.07 $X2=4.8
+ $Y2=8.14
cc_104 N_VPB_M1018_b N_A_1197_107#_c_362_n 0.00993716f $X=6.335 $Y=2.465
+ $X2=5.28 $Y2=8.14
cc_105 N_VPB_c_101_p N_A_1197_107#_c_362_n 0.00533646f $X=10.32 $Y=4.07 $X2=5.28
+ $Y2=8.14
cc_106 N_VPB_c_92_n N_A_1197_107#_c_362_n 0.00243411f $X=10.32 $Y=4.07 $X2=5.28
+ $Y2=8.14
cc_107 N_VPB_M1018_b N_A_772_151#_c_430_n 0.078156f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_108 N_VPB_M1018_b N_A_504_1221#_c_504_n 0.0309838f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_109 N_VPB_M1018_b N_A_504_1221#_c_517_n 0.0267665f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_VPB_c_101_p N_A_504_1221#_c_517_n 0.0181139f $X=10.32 $Y=4.07 $X2=0
+ $Y2=0
cc_111 N_VPB_c_92_n N_A_504_1221#_c_517_n 0.00970178f $X=10.32 $Y=4.07 $X2=0
+ $Y2=0
cc_112 N_VPB_M1018_b N_A_504_1221#_c_505_n 0.0336745f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_VPB_M1018_b N_A_504_1221#_c_521_n 0.0981784f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_114 N_VPB_c_101_p N_A_504_1221#_c_521_n 0.00523258f $X=10.32 $Y=4.07 $X2=0
+ $Y2=0
cc_115 N_VPB_c_92_n N_A_504_1221#_c_521_n 0.00914126f $X=10.32 $Y=4.07 $X2=0
+ $Y2=0
cc_116 N_VPB_M1018_b N_A_504_1221#_c_510_n 0.0559093f $X=6.335 $Y=2.465
+ $X2=10.32 $Y2=8.14
cc_117 N_VPB_c_92_n N_A_504_1221#_c_510_n 0.0308152f $X=10.32 $Y=4.07 $X2=10.32
+ $Y2=8.14
cc_118 N_VPB_M1018_b N_A_504_1221#_c_526_n 0.0828797f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_119 N_VPB_M1018_b N_A_504_1221#_c_511_n 0.0094031f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_VPB_M1018_b N_A_504_1221#_c_528_n 0.00377304f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_121 N_VPB_M1018_b N_A_504_1221#_c_529_n 0.138015f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_122 N_VPB_M1018_b N_A_504_1221#_c_514_n 0.0148513f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_123 N_VPB_c_92_n N_A_504_1221#_c_514_n 0.00180482f $X=10.32 $Y=4.07 $X2=0
+ $Y2=0
cc_124 N_VPB_M1018_b N_A_504_1221#_c_532_n 0.00504693f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_VPB_M1018_b N_A_504_1221#_c_515_n 0.00270883f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_126 N_VPB_M1018_b N_A_1711_885#_M1001_g 0.0571881f $X=6.335 $Y=2.465
+ $X2=-0.33 $Y2=-0.265
cc_127 N_VPB_c_101_p N_A_1711_885#_M1001_g 0.0175857f $X=10.32 $Y=4.07 $X2=-0.33
+ $Y2=-0.265
cc_128 N_VPB_c_92_n N_A_1711_885#_M1001_g 0.00970178f $X=10.32 $Y=4.07 $X2=-0.33
+ $Y2=-0.265
cc_129 N_VPB_M1018_b N_A_1711_885#_c_616_n 0.0232401f $X=6.335 $Y=2.465 $X2=0.24
+ $Y2=0
cc_130 N_VPB_c_101_p N_A_1711_885#_c_616_n 0.0158392f $X=10.32 $Y=4.07 $X2=0.24
+ $Y2=0
cc_131 N_VPB_c_92_n N_A_1711_885#_c_616_n 0.00101808f $X=10.32 $Y=4.07 $X2=0.24
+ $Y2=0
cc_132 N_VPB_M1018_b N_A_1711_885#_c_611_n 0.00203039f $X=6.335 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_VPB_M1018_b N_A_1711_885#_c_612_n 0.00832153f $X=6.335 $Y=2.465
+ $X2=0.24 $Y2=8.14
cc_134 N_VPB_M1018_b N_VPWR_c_657_n 0.00823544f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_135 N_VPB_c_101_p N_VPWR_c_657_n 0.0274404f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_136 N_VPB_c_92_n N_VPWR_c_657_n 0.00213221f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_137 N_VPB_M1018_b N_VPWR_c_660_n 0.0406421f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_138 N_VPB_c_101_p N_VPWR_c_660_n 0.0254284f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_139 N_VPB_c_92_n N_VPWR_c_660_n 0.00166879f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_140 N_VPB_X20_noxref_D1 N_VPWR_c_655_n 0.0336658f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_141 N_VPB_M1018_b N_VPWR_c_655_n 0.0709744f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_142 N_VPB_c_91_n N_VPWR_c_655_n 0.00613319f $X=0.24 $Y=4.07 $X2=0 $Y2=0
cc_143 N_VPB_c_101_p N_VPWR_c_655_n 0.018878f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_144 N_VPB_c_92_n N_VPWR_c_655_n 1.11192f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_145 N_VPB_M1018_b N_VPWR_c_668_n 0.00453345f $X=6.335 $Y=2.465 $X2=0.24
+ $Y2=8.14
cc_146 N_VPB_c_101_p N_VPWR_c_668_n 0.0275229f $X=10.32 $Y=4.07 $X2=0.24
+ $Y2=8.14
cc_147 N_VPB_c_92_n N_VPWR_c_668_n 0.00222323f $X=10.32 $Y=4.07 $X2=0.24
+ $Y2=8.14
cc_148 N_VPB_X20_noxref_D1 N_VPWR_c_656_n 0.0565882f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_149 N_VPB_M1018_b N_VPWR_c_656_n 0.0412639f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_150 N_VPB_c_91_n N_VPWR_c_656_n 0.00613319f $X=0.24 $Y=4.07 $X2=0 $Y2=0
cc_151 N_VPB_c_101_p N_VPWR_c_656_n 0.013686f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_152 N_VPB_c_92_n N_VPWR_c_656_n 1.11364f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_153 N_VPB_M1018_b X 0.0077824f $X=6.335 $Y=2.465 $X2=-0.33 $Y2=-0.265
cc_154 N_VPB_M1018_b N_X_c_725_n 0.0518911f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_155 N_VPB_c_101_p N_X_c_725_n 0.0158392f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_156 N_VPB_c_92_n N_X_c_725_n 0.00101808f $X=10.32 $Y=4.07 $X2=0 $Y2=0
cc_157 N_VPB_M1018_b X 0.00990693f $X=6.335 $Y=2.465 $X2=0 $Y2=0
cc_158 N_LVPWR_M1004_b N_A_c_215_n 0.0176162f $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_159 N_LVPWR_M1004_b N_A_M1004_g 0.0225938f $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_160 N_LVPWR_c_167_p N_A_M1004_g 0.00135859f $X=3.57 $Y=2.33 $X2=0 $Y2=0
cc_161 LVPWR N_A_M1004_g 0.0109749f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_162 N_LVPWR_c_164_n N_A_M1004_g 0.00417272f $X=3.93 $Y=3.19 $X2=0 $Y2=0
cc_163 N_LVPWR_M1004_b N_A_c_217_n 6.60476e-19 $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_164 N_LVPWR_M1004_b N_A_c_219_n 0.00547003f $X=2.8 $Y=2.015 $X2=0.24 $Y2=0
cc_165 LVPWR N_A_404_1133#_M1004_s 5.28909e-19 $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_166 N_LVPWR_M1004_b N_A_404_1133#_M1017_g 0.0221724f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_167 N_LVPWR_c_167_p N_A_404_1133#_M1017_g 0.00208937f $X=3.57 $Y=2.33 $X2=0
+ $Y2=0
cc_168 LVPWR N_A_404_1133#_M1017_g 0.00767826f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_169 N_LVPWR_c_164_n N_A_404_1133#_M1017_g 0.0112605f $X=3.93 $Y=3.19 $X2=0
+ $Y2=0
cc_170 N_LVPWR_M1004_b N_A_404_1133#_c_254_n 0.00262762f $X=2.8 $Y=2.015
+ $X2=0.24 $Y2=0
cc_171 N_LVPWR_c_167_p N_A_404_1133#_c_254_n 0.00156473f $X=3.57 $Y=2.33
+ $X2=0.24 $Y2=0
cc_172 N_LVPWR_M1004_b N_A_404_1133#_c_255_n 0.0500919f $X=2.8 $Y=2.015 $X2=4.8
+ $Y2=0.058
cc_173 N_LVPWR_c_167_p N_A_404_1133#_c_255_n 8.98083e-19 $X=3.57 $Y=2.33 $X2=4.8
+ $Y2=0.058
cc_174 LVPWR N_A_404_1133#_c_255_n 0.0236806f $X=0.07 $Y=3.02 $X2=4.8 $Y2=0.058
cc_175 N_LVPWR_c_164_n N_A_404_1133#_c_255_n 0.0814701f $X=3.93 $Y=3.19 $X2=4.8
+ $Y2=0.058
cc_176 N_LVPWR_M1004_b N_A_404_1133#_c_272_n 0.0232362f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_177 N_LVPWR_c_167_p N_A_404_1133#_c_272_n 0.00429663f $X=3.57 $Y=2.33 $X2=0
+ $Y2=0
cc_178 N_LVPWR_c_167_p N_A_404_1133#_c_258_n 0.0229916f $X=3.57 $Y=2.33 $X2=0
+ $Y2=0
cc_179 N_LVPWR_M1004_b N_A_404_1133#_c_259_n 0.0124783f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_180 N_LVPWR_M1004_b N_A_404_1133#_c_276_n 0.016229f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_181 LVPWR N_A_404_1133#_c_276_n 0.0263553f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_182 LVPWR N_A_1197_107#_c_365_n 0.0149945f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_183 LVPWR N_A_1197_107#_c_350_n 0.0103948f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_184 LVPWR N_A_1197_107#_c_355_n 0.0277879f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_185 LVPWR N_A_1197_107#_c_351_n 0.0313648f $X=0.07 $Y=3.02 $X2=10.32 $Y2=8.14
cc_186 LVPWR N_A_1197_107#_c_369_n 0.0155178f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_187 LVPWR N_A_1197_107#_c_360_n 0.0180443f $X=0.07 $Y=3.02 $X2=4.8 $Y2=8.14
cc_188 LVPWR N_A_1197_107#_c_362_n 0.00998653f $X=0.07 $Y=3.02 $X2=5.28 $Y2=8.14
cc_189 LVPWR N_A_772_151#_M1017_d 0.00288751f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_190 LVPWR N_A_772_151#_c_430_n 0.0145666f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_191 N_LVPWR_M1004_b N_A_772_151#_c_434_n 0.00801775f $X=2.8 $Y=2.015 $X2=0
+ $Y2=0
cc_192 N_LVPWR_c_167_p N_A_772_151#_c_434_n 0.00252726f $X=3.57 $Y=2.33 $X2=0
+ $Y2=0
cc_193 LVPWR N_A_772_151#_c_434_n 0.0235018f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_194 LVPWR N_A_772_151#_c_443_n 0.0320105f $X=0.07 $Y=3.02 $X2=10.32 $Y2=8.14
cc_195 N_LVPWR_M1004_b N_A_772_151#_c_444_n 0.016687f $X=2.8 $Y=2.015 $X2=10.32
+ $Y2=0
cc_196 LVPWR N_A_772_151#_c_444_n 0.0115771f $X=0.07 $Y=3.02 $X2=10.32 $Y2=0
cc_197 N_LVPWR_c_164_n N_A_772_151#_c_444_n 0.0160139f $X=3.93 $Y=3.19 $X2=10.32
+ $Y2=0
cc_198 LVPWR N_A_772_151#_c_436_n 0.0360894f $X=0.07 $Y=3.02 $X2=0.24 $Y2=8.14
cc_199 LVPWR N_A_504_1221#_M1006_s 4.36537e-19 $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_200 LVPWR N_A_504_1221#_c_528_n 0.0151454f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_201 LVPWR N_A_504_1221#_c_514_n 0.0407311f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_202 LVPWR N_VPWR_c_660_n 0.0536317f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_203 N_LVPWR_M1004_b N_VPWR_c_655_n 0.00793792f $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_204 LVPWR N_VPWR_c_655_n 1.09632f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_205 N_LVPWR_c_164_n N_VPWR_c_655_n 0.0680381f $X=3.93 $Y=3.19 $X2=0 $Y2=0
cc_206 N_LVPWR_M1004_b N_VPWR_c_656_n 0.00618401f $X=2.8 $Y=2.015 $X2=0 $Y2=0
cc_207 N_LVPWR_c_164_n N_VPWR_c_656_n 0.0268368f $X=3.93 $Y=3.19 $X2=0 $Y2=0
cc_208 N_A_c_216_n N_A_404_1133#_c_250_n 0.014409f $X=3.355 $Y=1.705 $X2=0.24
+ $Y2=0
cc_209 N_A_M1004_g N_A_404_1133#_M1017_g 0.019196f $X=3.355 $Y=2.615 $X2=0 $Y2=0
cc_210 N_A_c_217_n N_A_404_1133#_c_254_n 0.0226068f $X=3.355 $Y=1.87 $X2=0.24
+ $Y2=0
cc_211 N_A_M1004_g N_A_404_1133#_c_255_n 0.00201071f $X=3.355 $Y=2.615 $X2=4.8
+ $Y2=0.058
cc_212 N_A_c_215_n N_A_404_1133#_c_257_n 0.00930167f $X=3.28 $Y=1.87 $X2=5.28
+ $Y2=8.14
cc_213 N_A_c_216_n N_A_404_1133#_c_257_n 0.00615095f $X=3.355 $Y=1.705 $X2=5.28
+ $Y2=8.14
cc_214 A N_A_404_1133#_c_257_n 0.0165667f $X=2.555 $Y=1.58 $X2=5.28 $Y2=8.14
cc_215 N_A_c_219_n N_A_404_1133#_c_257_n 0.00155799f $X=2.66 $Y=1.695 $X2=5.28
+ $Y2=8.14
cc_216 N_A_c_215_n N_A_404_1133#_c_272_n 0.00930167f $X=3.28 $Y=1.87 $X2=0 $Y2=0
cc_217 N_A_M1004_g N_A_404_1133#_c_272_n 0.00805052f $X=3.355 $Y=2.615 $X2=0
+ $Y2=0
cc_218 A N_A_404_1133#_c_272_n 0.015787f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_219 N_A_c_219_n N_A_404_1133#_c_272_n 0.00146896f $X=2.66 $Y=1.695 $X2=0
+ $Y2=0
cc_220 N_A_c_215_n N_A_404_1133#_c_258_n 0.00131023f $X=3.28 $Y=1.87 $X2=0 $Y2=0
cc_221 N_A_c_217_n N_A_404_1133#_c_258_n 0.0196537f $X=3.355 $Y=1.87 $X2=0 $Y2=0
cc_222 N_A_c_215_n N_A_404_1133#_c_292_n 0.0104509f $X=3.28 $Y=1.87 $X2=0 $Y2=0
cc_223 A N_A_404_1133#_c_292_n 0.0198664f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_224 N_A_M1004_g N_VPWR_c_655_n 3.17298e-19 $X=3.355 $Y=2.615 $X2=0 $Y2=0
cc_225 N_A_c_216_n N_VGND_c_742_n 0.00386936f $X=3.355 $Y=1.705 $X2=0.24
+ $Y2=8.14
cc_226 N_A_c_216_n N_VGND_c_756_n 0.00555051f $X=3.355 $Y=1.705 $X2=0 $Y2=0
cc_227 N_A_c_216_n N_VGND_c_761_n 0.00523016f $X=3.355 $Y=1.705 $X2=0 $Y2=0
cc_228 N_A_404_1133#_c_250_n N_A_772_151#_c_432_n 0.00286882f $X=3.785 $Y=1.705
+ $X2=0 $Y2=0
cc_229 N_A_404_1133#_c_250_n N_A_772_151#_c_433_n 0.00280304f $X=3.785 $Y=1.705
+ $X2=0.24 $Y2=8.14
cc_230 N_A_404_1133#_M1017_g N_A_772_151#_c_433_n 0.00253691f $X=3.785 $Y=2.615
+ $X2=0.24 $Y2=8.14
cc_231 N_A_404_1133#_c_258_n N_A_772_151#_c_433_n 0.020811f $X=4.145 $Y=1.87
+ $X2=0.24 $Y2=8.14
cc_232 N_A_404_1133#_c_259_n N_A_772_151#_c_433_n 0.00542196f $X=4.145 $Y=1.87
+ $X2=0.24 $Y2=8.14
cc_233 N_A_404_1133#_M1017_g N_A_772_151#_c_434_n 0.00123902f $X=3.785 $Y=2.615
+ $X2=0 $Y2=0
cc_234 N_A_404_1133#_c_258_n N_A_772_151#_c_434_n 0.0353505f $X=4.145 $Y=1.87
+ $X2=0 $Y2=0
cc_235 N_A_404_1133#_c_259_n N_A_772_151#_c_434_n 0.0105631f $X=4.145 $Y=1.87
+ $X2=0 $Y2=0
cc_236 N_A_404_1133#_c_258_n N_A_772_151#_c_435_n 0.0316368f $X=4.145 $Y=1.87
+ $X2=0 $Y2=0
cc_237 N_A_404_1133#_c_259_n N_A_772_151#_c_435_n 0.0102771f $X=4.145 $Y=1.87
+ $X2=0 $Y2=0
cc_238 N_A_404_1133#_c_247_n N_A_504_1221#_c_537_n 0.0381272f $X=2.27 $Y=5.995
+ $X2=0 $Y2=0
cc_239 N_A_404_1133#_c_248_n N_A_504_1221#_c_537_n 0.0401197f $X=3.05 $Y=5.995
+ $X2=0 $Y2=0
cc_240 N_A_404_1133#_c_252_n N_A_504_1221#_c_539_n 0.117263f $X=5.39 $Y=5.995
+ $X2=10.32 $Y2=8.14
cc_241 N_A_404_1133#_c_255_n N_A_504_1221#_c_539_n 0.0229895f $X=3.03 $Y=4.65
+ $X2=10.32 $Y2=8.14
cc_242 N_A_404_1133#_c_252_n N_A_504_1221#_c_507_n 0.0335781f $X=5.39 $Y=5.995
+ $X2=10.32 $Y2=8.14
cc_243 N_A_404_1133#_c_249_n N_A_504_1221#_c_542_n 0.0401197f $X=3.83 $Y=5.995
+ $X2=0 $Y2=0
cc_244 N_A_404_1133#_c_251_n N_A_504_1221#_c_542_n 0.0401197f $X=4.61 $Y=5.995
+ $X2=0 $Y2=0
cc_245 N_A_404_1133#_c_252_n N_A_504_1221#_c_544_n 0.124218f $X=5.39 $Y=5.995
+ $X2=4.8 $Y2=0.058
cc_246 N_A_404_1133#_c_252_n N_A_504_1221#_c_508_n 0.0429997f $X=5.39 $Y=5.995
+ $X2=0.24 $Y2=8.14
cc_247 N_A_404_1133#_c_252_n N_A_504_1221#_c_511_n 0.0100783f $X=5.39 $Y=5.995
+ $X2=0 $Y2=0
cc_248 N_A_404_1133#_c_252_n N_A_504_1221#_c_513_n 0.0175374f $X=5.39 $Y=5.995
+ $X2=0 $Y2=0
cc_249 N_A_404_1133#_c_255_n N_VPWR_c_655_n 0.0361756f $X=3.03 $Y=4.65 $X2=0
+ $Y2=0
cc_250 N_A_404_1133#_c_276_n N_VPWR_c_655_n 3.87848e-19 $X=3.075 $Y=3.055 $X2=0
+ $Y2=0
cc_251 N_A_404_1133#_c_255_n N_VPWR_c_656_n 0.0547753f $X=3.03 $Y=4.65 $X2=0
+ $Y2=0
cc_252 N_A_404_1133#_c_256_n N_VPWR_c_656_n 0.00922839f $X=3.03 $Y=4.65 $X2=0
+ $Y2=0
cc_253 N_A_404_1133#_c_247_n N_VGND_c_738_n 0.0146836f $X=2.27 $Y=5.995 $X2=0
+ $Y2=0
cc_254 N_A_404_1133#_c_248_n N_VGND_c_738_n 0.0146836f $X=3.05 $Y=5.995 $X2=0
+ $Y2=0
cc_255 N_A_404_1133#_c_247_n N_VGND_c_740_n 0.0034209f $X=2.27 $Y=5.995 $X2=0
+ $Y2=0
cc_256 N_A_404_1133#_c_250_n N_VGND_c_742_n 0.00386936f $X=3.785 $Y=1.705
+ $X2=0.24 $Y2=8.14
cc_257 N_A_404_1133#_c_254_n N_VGND_c_742_n 0.00139629f $X=3.75 $Y=1.87 $X2=0.24
+ $Y2=8.14
cc_258 N_A_404_1133#_c_257_n N_VGND_c_742_n 0.001542f $X=3.14 $Y=0.9 $X2=0.24
+ $Y2=8.14
cc_259 N_A_404_1133#_c_258_n N_VGND_c_742_n 0.0179406f $X=4.145 $Y=1.87 $X2=0.24
+ $Y2=8.14
cc_260 N_A_404_1133#_c_249_n N_VGND_c_743_n 0.0146836f $X=3.83 $Y=5.995 $X2=0
+ $Y2=0
cc_261 N_A_404_1133#_c_251_n N_VGND_c_743_n 0.0179057f $X=4.61 $Y=5.995 $X2=0
+ $Y2=0
cc_262 N_A_404_1133#_c_252_n N_VGND_c_743_n 0.00366145f $X=5.39 $Y=5.995 $X2=0
+ $Y2=0
cc_263 N_A_404_1133#_c_248_n N_VGND_c_751_n 0.00322203f $X=3.05 $Y=5.995
+ $X2=0.24 $Y2=0
cc_264 N_A_404_1133#_c_249_n N_VGND_c_751_n 0.00322203f $X=3.83 $Y=5.995
+ $X2=0.24 $Y2=0
cc_265 N_A_404_1133#_c_247_n N_VGND_c_755_n 0.0665921f $X=2.27 $Y=5.995 $X2=5.28
+ $Y2=8.14
cc_266 N_A_404_1133#_c_248_n N_VGND_c_755_n 0.00132352f $X=3.05 $Y=5.995
+ $X2=5.28 $Y2=8.14
cc_267 N_A_404_1133#_c_257_n N_VGND_c_756_n 0.0123012f $X=3.14 $Y=0.9 $X2=0
+ $Y2=0
cc_268 N_A_404_1133#_c_247_n N_VGND_c_787_n 0.00129485f $X=2.27 $Y=5.995 $X2=0
+ $Y2=0
cc_269 N_A_404_1133#_c_248_n N_VGND_c_787_n 0.0567946f $X=3.05 $Y=5.995 $X2=0
+ $Y2=0
cc_270 N_A_404_1133#_c_249_n N_VGND_c_787_n 0.0567946f $X=3.83 $Y=5.995 $X2=0
+ $Y2=0
cc_271 N_A_404_1133#_c_251_n N_VGND_c_787_n 0.00129485f $X=4.61 $Y=5.995 $X2=0
+ $Y2=0
cc_272 N_A_404_1133#_c_252_n N_VGND_c_787_n 0.00232957f $X=5.39 $Y=5.995 $X2=0
+ $Y2=0
cc_273 N_A_404_1133#_c_250_n N_VGND_c_758_n 0.00555051f $X=3.785 $Y=1.705 $X2=0
+ $Y2=0
cc_274 N_A_404_1133#_c_249_n N_VGND_c_793_n 0.00129485f $X=3.83 $Y=5.995 $X2=0
+ $Y2=0
cc_275 N_A_404_1133#_c_251_n N_VGND_c_793_n 0.0567946f $X=4.61 $Y=5.995 $X2=0
+ $Y2=0
cc_276 N_A_404_1133#_c_252_n N_VGND_c_793_n 0.0596044f $X=5.39 $Y=5.995 $X2=0
+ $Y2=0
cc_277 N_A_404_1133#_c_250_n N_VGND_c_761_n 0.00523016f $X=3.785 $Y=1.705 $X2=0
+ $Y2=0
cc_278 N_A_404_1133#_c_257_n N_VGND_c_761_n 0.0105954f $X=3.14 $Y=0.9 $X2=0
+ $Y2=0
cc_279 N_A_404_1133#_c_247_n N_VGND_c_765_n 0.0157032f $X=2.27 $Y=5.995 $X2=0
+ $Y2=0
cc_280 N_A_404_1133#_c_248_n N_VGND_c_765_n 0.0157032f $X=3.05 $Y=5.995 $X2=0
+ $Y2=0
cc_281 N_A_404_1133#_c_249_n N_VGND_c_765_n 0.0157032f $X=3.83 $Y=5.995 $X2=0
+ $Y2=0
cc_282 N_A_404_1133#_c_251_n N_VGND_c_765_n 0.0157032f $X=4.61 $Y=5.995 $X2=0
+ $Y2=0
cc_283 N_A_404_1133#_c_252_n N_VGND_c_765_n 0.0212017f $X=5.39 $Y=5.995 $X2=0
+ $Y2=0
cc_284 N_A_1197_107#_c_372_p N_A_772_151#_c_426_n 0.0401197f $X=6.125 $Y=0.68
+ $X2=0 $Y2=0
cc_285 N_A_1197_107#_c_372_p N_A_772_151#_c_427_n 0.0401197f $X=6.125 $Y=0.68
+ $X2=0 $Y2=0
cc_286 N_A_1197_107#_c_374_p N_A_772_151#_c_428_n 0.0401197f $X=7.685 $Y=0.68
+ $X2=0 $Y2=0
cc_287 N_A_1197_107#_c_374_p N_A_772_151#_c_429_n 0.0401197f $X=7.685 $Y=0.68
+ $X2=0.24 $Y2=0
cc_288 N_A_1197_107#_c_365_n N_A_772_151#_c_430_n 0.0595693f $X=7.165 $Y=2.31
+ $X2=0 $Y2=0
cc_289 N_A_1197_107#_c_350_n N_A_772_151#_c_430_n 0.0200524f $X=6.29 $Y=2.31
+ $X2=0 $Y2=0
cc_290 N_A_1197_107#_c_355_n N_A_772_151#_c_430_n 0.00172854f $X=7.33 $Y=3.395
+ $X2=0 $Y2=0
cc_291 N_A_1197_107#_c_374_p N_A_772_151#_c_430_n 0.00443612f $X=7.685 $Y=0.68
+ $X2=0 $Y2=0
cc_292 N_A_1197_107#_c_351_n N_A_772_151#_c_430_n 0.0994932f $X=9.08 $Y=2.31
+ $X2=0 $Y2=0
cc_293 N_A_1197_107#_c_369_n N_A_772_151#_c_430_n 0.0425514f $X=7.85 $Y=2.31
+ $X2=0 $Y2=0
cc_294 N_A_1197_107#_c_352_n N_A_772_151#_c_430_n 0.0429997f $X=9.245 $Y=0.68
+ $X2=0 $Y2=0
cc_295 N_A_1197_107#_c_360_n N_A_772_151#_c_430_n 0.0712039f $X=7.33 $Y=3.56
+ $X2=0 $Y2=0
cc_296 N_A_1197_107#_c_350_n N_A_772_151#_c_443_n 0.0277655f $X=6.29 $Y=2.31
+ $X2=10.32 $Y2=8.14
cc_297 N_A_1197_107#_c_354_n N_A_504_1221#_c_521_n 0.0456276f $X=7.165 $Y=4.635
+ $X2=0 $Y2=0
cc_298 N_A_1197_107#_c_356_n N_A_504_1221#_c_521_n 0.017714f $X=7.33 $Y=4.47
+ $X2=0 $Y2=0
cc_299 N_A_1197_107#_c_360_n N_A_504_1221#_c_521_n 0.0107531f $X=7.33 $Y=3.56
+ $X2=0 $Y2=0
cc_300 N_A_1197_107#_c_362_n N_A_504_1221#_c_521_n 0.00384278f $X=7.67 $Y=3.56
+ $X2=0 $Y2=0
cc_301 N_A_1197_107#_c_354_n N_A_504_1221#_c_510_n 0.0250923f $X=7.165 $Y=4.635
+ $X2=10.32 $Y2=8.14
cc_302 N_A_1197_107#_c_356_n N_A_504_1221#_c_510_n 0.0144968f $X=7.33 $Y=4.47
+ $X2=10.32 $Y2=8.14
cc_303 N_A_1197_107#_c_360_n N_A_504_1221#_c_510_n 9.41636e-19 $X=7.33 $Y=3.56
+ $X2=10.32 $Y2=8.14
cc_304 N_A_1197_107#_c_362_n N_A_504_1221#_c_510_n 0.00442739f $X=7.67 $Y=3.56
+ $X2=10.32 $Y2=8.14
cc_305 N_A_1197_107#_c_365_n N_A_504_1221#_c_528_n 0.0146618f $X=7.165 $Y=2.31
+ $X2=0 $Y2=0
cc_306 N_A_1197_107#_c_355_n N_A_504_1221#_c_528_n 0.0150559f $X=7.33 $Y=3.395
+ $X2=0 $Y2=0
cc_307 N_A_1197_107#_c_360_n N_A_504_1221#_c_528_n 7.80231e-19 $X=7.33 $Y=3.56
+ $X2=0 $Y2=0
cc_308 N_A_1197_107#_c_365_n N_A_504_1221#_c_514_n 0.00518824f $X=7.165 $Y=2.31
+ $X2=0 $Y2=0
cc_309 N_A_1197_107#_c_350_n N_A_504_1221#_c_514_n 0.00152927f $X=6.29 $Y=2.31
+ $X2=0 $Y2=0
cc_310 N_A_1197_107#_c_355_n N_A_504_1221#_c_514_n 0.01755f $X=7.33 $Y=3.395
+ $X2=0 $Y2=0
cc_311 N_A_1197_107#_c_360_n N_A_504_1221#_c_514_n 0.00675584f $X=7.33 $Y=3.56
+ $X2=0 $Y2=0
cc_312 N_A_1197_107#_c_362_n N_A_504_1221#_c_514_n 0.00570418f $X=7.67 $Y=3.56
+ $X2=0 $Y2=0
cc_313 N_A_1197_107#_c_354_n N_VPWR_c_657_n 0.0154109f $X=7.165 $Y=4.635 $X2=0
+ $Y2=0
cc_314 N_A_1197_107#_c_356_n N_VPWR_c_657_n 0.002585f $X=7.33 $Y=4.47 $X2=0
+ $Y2=0
cc_315 N_A_1197_107#_c_355_n N_VPWR_c_660_n 0.0144973f $X=7.33 $Y=3.395 $X2=0
+ $Y2=0
cc_316 N_A_1197_107#_c_351_n N_VPWR_c_660_n 0.0279184f $X=9.08 $Y=2.31 $X2=0
+ $Y2=0
cc_317 N_A_1197_107#_c_360_n N_VPWR_c_660_n 0.0230299f $X=7.33 $Y=3.56 $X2=0
+ $Y2=0
cc_318 N_A_1197_107#_c_362_n N_VPWR_c_660_n 0.0224772f $X=7.67 $Y=3.56 $X2=0
+ $Y2=0
cc_319 N_A_1197_107#_c_355_n N_VPWR_c_655_n 3.90571e-19 $X=7.33 $Y=3.395 $X2=0
+ $Y2=0
cc_320 N_A_1197_107#_c_356_n N_VPWR_c_655_n 0.00532287f $X=7.33 $Y=4.47 $X2=0
+ $Y2=0
cc_321 N_A_1197_107#_c_360_n N_VPWR_c_655_n 0.0153452f $X=7.33 $Y=3.56 $X2=0
+ $Y2=0
cc_322 N_A_1197_107#_c_362_n N_VPWR_c_655_n 0.0496017f $X=7.67 $Y=3.56 $X2=0
+ $Y2=0
cc_323 N_A_1197_107#_M1018_s N_VPWR_c_656_n 8.34083e-19 $X=6.665 $Y=4.425 $X2=0
+ $Y2=0
cc_324 N_A_1197_107#_c_354_n N_VPWR_c_656_n 0.074493f $X=7.165 $Y=4.635 $X2=0
+ $Y2=0
cc_325 N_A_1197_107#_c_356_n N_VPWR_c_656_n 0.0159329f $X=7.33 $Y=4.47 $X2=0
+ $Y2=0
cc_326 N_A_1197_107#_c_372_p N_VGND_c_745_n 0.0211458f $X=6.125 $Y=0.68 $X2=0
+ $Y2=0
cc_327 N_A_1197_107#_c_374_p N_VGND_c_749_n 0.0211458f $X=7.685 $Y=0.68
+ $X2=10.32 $Y2=8.14
cc_328 N_A_1197_107#_c_372_p N_VGND_c_760_n 0.0648349f $X=6.125 $Y=0.68 $X2=0
+ $Y2=0
cc_329 N_A_1197_107#_c_372_p N_VGND_c_806_n 0.0648349f $X=6.125 $Y=0.68 $X2=0
+ $Y2=0
cc_330 N_A_1197_107#_c_365_n N_VGND_c_806_n 0.0424704f $X=7.165 $Y=2.31 $X2=0
+ $Y2=0
cc_331 N_A_1197_107#_c_374_p N_VGND_c_806_n 0.0648349f $X=7.685 $Y=0.68 $X2=0
+ $Y2=0
cc_332 N_A_1197_107#_c_374_p N_VGND_c_809_n 0.0648349f $X=7.685 $Y=0.68 $X2=0
+ $Y2=0
cc_333 N_A_1197_107#_c_351_n N_VGND_c_809_n 0.0425081f $X=9.08 $Y=2.31 $X2=0
+ $Y2=0
cc_334 N_A_1197_107#_c_352_n N_VGND_c_809_n 0.0673371f $X=9.245 $Y=0.68 $X2=0
+ $Y2=0
cc_335 N_A_1197_107#_c_372_p N_VGND_c_761_n 0.0240827f $X=6.125 $Y=0.68 $X2=0
+ $Y2=0
cc_336 N_A_1197_107#_c_374_p N_VGND_c_761_n 0.0240827f $X=7.685 $Y=0.68 $X2=0
+ $Y2=0
cc_337 N_A_1197_107#_c_352_n N_VGND_c_761_n 0.0337346f $X=9.245 $Y=0.68 $X2=0
+ $Y2=0
cc_338 N_A_772_151#_c_430_n N_A_504_1221#_c_528_n 0.0075528f $X=8.855 $Y=2.145
+ $X2=0 $Y2=0
cc_339 N_A_772_151#_c_430_n N_A_504_1221#_c_514_n 0.00656921f $X=8.855 $Y=2.145
+ $X2=0 $Y2=0
cc_340 N_A_772_151#_c_430_n N_VPWR_c_660_n 0.0136723f $X=8.855 $Y=2.145 $X2=0
+ $Y2=0
cc_341 N_A_772_151#_c_432_n N_VGND_c_742_n 0.00154986f $X=4 $Y=0.9 $X2=0.24
+ $Y2=8.14
cc_342 N_A_772_151#_c_426_n N_VGND_c_745_n 0.0146836f $X=5.735 $Y=2.145 $X2=0
+ $Y2=0
cc_343 N_A_772_151#_c_427_n N_VGND_c_745_n 0.0146836f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_344 N_A_772_151#_c_426_n N_VGND_c_747_n 0.0034209f $X=5.735 $Y=2.145
+ $X2=10.32 $Y2=8.14
cc_345 N_A_772_151#_c_428_n N_VGND_c_749_n 0.0146836f $X=7.295 $Y=2.145
+ $X2=10.32 $Y2=8.14
cc_346 N_A_772_151#_c_429_n N_VGND_c_749_n 0.0179057f $X=8.075 $Y=2.145
+ $X2=10.32 $Y2=8.14
cc_347 N_A_772_151#_c_430_n N_VGND_c_749_n 0.00366145f $X=8.855 $Y=2.145
+ $X2=10.32 $Y2=8.14
cc_348 N_A_772_151#_c_427_n N_VGND_c_753_n 0.00322203f $X=6.515 $Y=2.145
+ $X2=5.28 $Y2=0
cc_349 N_A_772_151#_c_428_n N_VGND_c_753_n 0.00322203f $X=7.295 $Y=2.145
+ $X2=5.28 $Y2=0
cc_350 N_A_772_151#_c_432_n N_VGND_c_758_n 0.0120367f $X=4 $Y=0.9 $X2=0 $Y2=0
cc_351 N_A_772_151#_c_426_n N_VGND_c_760_n 0.0582646f $X=5.735 $Y=2.145 $X2=0
+ $Y2=0
cc_352 N_A_772_151#_c_427_n N_VGND_c_760_n 0.00129485f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_353 N_A_772_151#_c_433_n N_VGND_c_760_n 0.027388f $X=4.645 $Y=2.145 $X2=0
+ $Y2=0
cc_354 N_A_772_151#_c_443_n N_VGND_c_760_n 0.0457912f $X=5.625 $Y=2.31 $X2=0
+ $Y2=0
cc_355 N_A_772_151#_c_435_n N_VGND_c_760_n 0.0237705f $X=4.645 $Y=1.41 $X2=0
+ $Y2=0
cc_356 N_A_772_151#_c_436_n N_VGND_c_760_n 0.00991638f $X=5.485 $Y=2.31 $X2=0
+ $Y2=0
cc_357 N_A_772_151#_c_426_n N_VGND_c_806_n 0.00129485f $X=5.735 $Y=2.145 $X2=0
+ $Y2=0
cc_358 N_A_772_151#_c_427_n N_VGND_c_806_n 0.0567946f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_359 N_A_772_151#_c_428_n N_VGND_c_806_n 0.0567946f $X=7.295 $Y=2.145 $X2=0
+ $Y2=0
cc_360 N_A_772_151#_c_429_n N_VGND_c_806_n 0.00129485f $X=8.075 $Y=2.145 $X2=0
+ $Y2=0
cc_361 N_A_772_151#_c_430_n N_VGND_c_806_n 0.00232957f $X=8.855 $Y=2.145 $X2=0
+ $Y2=0
cc_362 N_A_772_151#_c_428_n N_VGND_c_809_n 0.00129485f $X=7.295 $Y=2.145 $X2=0
+ $Y2=0
cc_363 N_A_772_151#_c_429_n N_VGND_c_809_n 0.0567946f $X=8.075 $Y=2.145 $X2=0
+ $Y2=0
cc_364 N_A_772_151#_c_430_n N_VGND_c_809_n 0.0596044f $X=8.855 $Y=2.145 $X2=0
+ $Y2=0
cc_365 N_A_772_151#_c_426_n N_VGND_c_761_n 0.0157032f $X=5.735 $Y=2.145 $X2=0
+ $Y2=0
cc_366 N_A_772_151#_c_427_n N_VGND_c_761_n 0.0157032f $X=6.515 $Y=2.145 $X2=0
+ $Y2=0
cc_367 N_A_772_151#_c_428_n N_VGND_c_761_n 0.0157032f $X=7.295 $Y=2.145 $X2=0
+ $Y2=0
cc_368 N_A_772_151#_c_429_n N_VGND_c_761_n 0.0157032f $X=8.075 $Y=2.145 $X2=0
+ $Y2=0
cc_369 N_A_772_151#_c_430_n N_VGND_c_761_n 0.0212017f $X=8.855 $Y=2.145 $X2=0
+ $Y2=0
cc_370 N_A_772_151#_c_432_n N_VGND_c_761_n 0.0112977f $X=4 $Y=0.9 $X2=0 $Y2=0
cc_371 N_A_504_1221#_c_517_n N_A_1711_885#_M1001_g 0.0140023f $X=9.07 $Y=5.805
+ $X2=-0.33 $Y2=-0.265
cc_372 N_A_504_1221#_c_505_n N_A_1711_885#_M1001_g 0.00729839f $X=9.07 $Y=6.975
+ $X2=-0.33 $Y2=-0.265
cc_373 N_A_504_1221#_c_505_n N_A_1711_885#_M1005_g 0.0214213f $X=9.07 $Y=6.975
+ $X2=0 $Y2=0
cc_374 N_A_504_1221#_c_517_n N_A_1711_885#_c_616_n 0.0323219f $X=9.07 $Y=5.805
+ $X2=0.24 $Y2=0
cc_375 N_A_504_1221#_c_505_n N_A_1711_885#_c_616_n 0.0223325f $X=9.07 $Y=6.975
+ $X2=0.24 $Y2=0
cc_376 N_A_504_1221#_c_521_n N_A_1711_885#_c_616_n 0.0198137f $X=7.825 $Y=4.635
+ $X2=0.24 $Y2=0
cc_377 N_A_504_1221#_c_572_p N_A_1711_885#_c_616_n 0.0156097f $X=7.825 $Y=5.37
+ $X2=0.24 $Y2=0
cc_378 N_A_504_1221#_c_529_n N_A_1711_885#_c_616_n 0.00597659f $X=7.825 $Y=5.37
+ $X2=0.24 $Y2=0
cc_379 N_A_504_1221#_c_512_n N_A_1711_885#_c_616_n 0.00776343f $X=7.825 $Y=6.39
+ $X2=0.24 $Y2=0
cc_380 N_A_504_1221#_c_532_n N_A_1711_885#_c_616_n 0.0118044f $X=7.825 $Y=5.83
+ $X2=0.24 $Y2=0
cc_381 N_A_504_1221#_c_505_n N_A_1711_885#_c_609_n 0.0389021f $X=9.07 $Y=6.975
+ $X2=10.32 $Y2=0
cc_382 N_A_504_1221#_c_505_n N_A_1711_885#_c_611_n 0.0533323f $X=9.07 $Y=6.975
+ $X2=0 $Y2=0
cc_383 N_A_504_1221#_c_505_n N_A_1711_885#_c_612_n 0.0216171f $X=9.07 $Y=6.975
+ $X2=0.24 $Y2=8.14
cc_384 N_A_504_1221#_c_504_n N_A_1711_885#_c_634_n 0.0311995f $X=8.82 $Y=6.39
+ $X2=0 $Y2=0
cc_385 N_A_504_1221#_c_505_n N_A_1711_885#_c_634_n 7.76856e-19 $X=9.07 $Y=6.975
+ $X2=0 $Y2=0
cc_386 N_A_504_1221#_c_512_n N_A_1711_885#_c_634_n 0.0104394f $X=7.825 $Y=6.39
+ $X2=0 $Y2=0
cc_387 N_A_504_1221#_c_517_n N_VPWR_c_657_n 5.056e-19 $X=9.07 $Y=5.805 $X2=0
+ $Y2=0
cc_388 N_A_504_1221#_c_521_n N_VPWR_c_657_n 0.0211446f $X=7.825 $Y=4.635 $X2=0
+ $Y2=0
cc_389 N_A_504_1221#_c_572_p N_VPWR_c_657_n 0.00780656f $X=7.825 $Y=5.37 $X2=0
+ $Y2=0
cc_390 N_A_504_1221#_c_510_n N_VPWR_c_655_n 0.0383422f $X=6.35 $Y=5.665 $X2=0
+ $Y2=0
cc_391 N_A_504_1221#_c_514_n N_VPWR_c_655_n 0.0280942f $X=6.83 $Y=3.3 $X2=0
+ $Y2=0
cc_392 N_A_504_1221#_c_517_n N_VPWR_c_668_n 0.0442244f $X=9.07 $Y=5.805 $X2=0.24
+ $Y2=8.14
cc_393 N_A_504_1221#_c_505_n N_VPWR_c_668_n 0.00618186f $X=9.07 $Y=6.975
+ $X2=0.24 $Y2=8.14
cc_394 N_A_504_1221#_c_517_n N_VPWR_c_656_n 0.0223603f $X=9.07 $Y=5.805 $X2=0
+ $Y2=0
cc_395 N_A_504_1221#_c_521_n N_VPWR_c_656_n 0.0143374f $X=7.825 $Y=4.635 $X2=0
+ $Y2=0
cc_396 N_A_504_1221#_c_510_n N_VPWR_c_656_n 0.0557507f $X=6.35 $Y=5.665 $X2=0
+ $Y2=0
cc_397 N_A_504_1221#_c_572_p N_VPWR_c_656_n 0.00455398f $X=7.825 $Y=5.37 $X2=0
+ $Y2=0
cc_398 N_A_504_1221#_c_537_n N_VGND_c_738_n 0.0211458f $X=2.66 $Y=6.25 $X2=0
+ $Y2=0
cc_399 N_A_504_1221#_c_542_n N_VGND_c_743_n 0.0211458f $X=4.22 $Y=6.25 $X2=0
+ $Y2=0
cc_400 N_A_504_1221#_c_537_n N_VGND_c_755_n 0.0686214f $X=2.66 $Y=6.25 $X2=5.28
+ $Y2=8.14
cc_401 N_A_504_1221#_c_537_n N_VGND_c_787_n 0.0648349f $X=2.66 $Y=6.25 $X2=0
+ $Y2=0
cc_402 N_A_504_1221#_c_539_n N_VGND_c_787_n 0.0425081f $X=4.055 $Y=5.83 $X2=0
+ $Y2=0
cc_403 N_A_504_1221#_c_542_n N_VGND_c_787_n 0.0648349f $X=4.22 $Y=6.25 $X2=0
+ $Y2=0
cc_404 N_A_504_1221#_c_542_n N_VGND_c_793_n 0.0648349f $X=4.22 $Y=6.25 $X2=0
+ $Y2=0
cc_405 N_A_504_1221#_c_544_n N_VGND_c_793_n 0.0425081f $X=5.615 $Y=5.83 $X2=0
+ $Y2=0
cc_406 N_A_504_1221#_c_508_n N_VGND_c_793_n 0.0673371f $X=5.78 $Y=6.25 $X2=0
+ $Y2=0
cc_407 N_A_504_1221#_c_505_n N_VGND_c_763_n 0.0340179f $X=9.07 $Y=6.975 $X2=0
+ $Y2=0
cc_408 N_A_504_1221#_c_505_n N_VGND_c_765_n 0.0241606f $X=9.07 $Y=6.975 $X2=0
+ $Y2=0
cc_409 N_A_504_1221#_c_537_n N_VGND_c_765_n 0.0240827f $X=2.66 $Y=6.25 $X2=0
+ $Y2=0
cc_410 N_A_504_1221#_c_542_n N_VGND_c_765_n 0.0240827f $X=4.22 $Y=6.25 $X2=0
+ $Y2=0
cc_411 N_A_504_1221#_c_508_n N_VGND_c_765_n 0.0337346f $X=5.78 $Y=6.25 $X2=0
+ $Y2=0
cc_412 N_A_1711_885#_c_616_n N_VPWR_c_657_n 0.0302319f $X=8.68 $Y=4.57 $X2=0
+ $Y2=0
cc_413 N_A_1711_885#_M1001_g N_VPWR_c_668_n 0.0563666f $X=9.895 $Y=5.175
+ $X2=0.24 $Y2=8.14
cc_414 N_A_1711_885#_c_616_n N_VPWR_c_668_n 0.0606653f $X=8.68 $Y=4.57 $X2=0.24
+ $Y2=8.14
cc_415 N_A_1711_885#_c_611_n N_VPWR_c_668_n 0.0338611f $X=9.955 $Y=6.39 $X2=0.24
+ $Y2=8.14
cc_416 N_A_1711_885#_c_612_n N_VPWR_c_668_n 0.00426906f $X=9.955 $Y=6.39
+ $X2=0.24 $Y2=8.14
cc_417 N_A_1711_885#_M1001_g N_VPWR_c_656_n 0.0193385f $X=9.895 $Y=5.175 $X2=0
+ $Y2=0
cc_418 N_A_1711_885#_c_616_n N_VPWR_c_656_n 0.0396431f $X=8.68 $Y=4.57 $X2=0
+ $Y2=0
cc_419 N_A_1711_885#_M1001_g X 0.00967557f $X=9.895 $Y=5.175 $X2=-0.33
+ $Y2=-0.265
cc_420 N_A_1711_885#_M1005_g X 0.0271496f $X=9.895 $Y=7.23 $X2=0 $Y2=0
cc_421 N_A_1711_885#_M1001_g N_X_c_725_n 0.032138f $X=9.895 $Y=5.175 $X2=0 $Y2=0
cc_422 N_A_1711_885#_M1001_g X 0.0254153f $X=9.895 $Y=5.175 $X2=0 $Y2=0
cc_423 N_A_1711_885#_c_611_n X 0.0268756f $X=9.955 $Y=6.39 $X2=0 $Y2=0
cc_424 N_A_1711_885#_M1005_g N_VGND_c_763_n 0.0387435f $X=9.895 $Y=7.23 $X2=0
+ $Y2=0
cc_425 N_A_1711_885#_c_609_n N_VGND_c_763_n 0.0317368f $X=8.68 $Y=7 $X2=0 $Y2=0
cc_426 N_A_1711_885#_c_611_n N_VGND_c_763_n 0.0338611f $X=9.955 $Y=6.39 $X2=0
+ $Y2=0
cc_427 N_A_1711_885#_c_612_n N_VGND_c_763_n 0.00426906f $X=9.955 $Y=6.39 $X2=0
+ $Y2=0
cc_428 N_A_1711_885#_M1005_g N_VGND_c_765_n 0.0208706f $X=9.895 $Y=7.23 $X2=0
+ $Y2=0
cc_429 N_A_1711_885#_c_609_n N_VGND_c_765_n 0.0338942f $X=8.68 $Y=7 $X2=0 $Y2=0
cc_430 N_VPWR_c_668_n N_X_c_725_n 0.0682113f $X=9.505 $Y=4.57 $X2=0 $Y2=0
cc_431 N_VPWR_c_656_n N_X_c_725_n 0.0434272f $X=9.685 $Y=4.58 $X2=0 $Y2=0
cc_432 X N_VGND_c_763_n 0.0356028f $X=10.235 $Y=6.76 $X2=0 $Y2=0
cc_433 X N_VGND_c_765_n 0.0326456f $X=10.235 $Y=6.76 $X2=0 $Y2=0
