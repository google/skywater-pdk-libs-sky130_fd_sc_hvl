* File: sky130_fd_sc_hvl__einvp_1.pxi.spice
* Created: Fri Aug 28 09:35:32 2020
* 
x_PM_SKY130_FD_SC_HVL__EINVP_1%VNB N_VNB_M1005_b VNB N_VNB_c_4_p VNB
+ PM_SKY130_FD_SC_HVL__EINVP_1%VNB
x_PM_SKY130_FD_SC_HVL__EINVP_1%VPB N_VPB_M1002_b VPB N_VPB_c_34_p VPB
+ PM_SKY130_FD_SC_HVL__EINVP_1%VPB
x_PM_SKY130_FD_SC_HVL__EINVP_1%TE N_TE_M1005_g N_TE_M1002_g N_TE_c_52_n
+ N_TE_c_53_n N_TE_c_55_n N_TE_M1001_g TE TE N_TE_c_57_n
+ PM_SKY130_FD_SC_HVL__EINVP_1%TE
x_PM_SKY130_FD_SC_HVL__EINVP_1%A_30_189# N_A_30_189#_M1005_s N_A_30_189#_M1002_s
+ N_A_30_189#_M1004_g N_A_30_189#_c_89_n N_A_30_189#_c_90_n N_A_30_189#_c_94_n
+ N_A_30_189#_c_106_n N_A_30_189#_c_91_n N_A_30_189#_c_96_n N_A_30_189#_c_92_n
+ N_A_30_189#_c_98_n N_A_30_189#_c_99_n PM_SKY130_FD_SC_HVL__EINVP_1%A_30_189#
x_PM_SKY130_FD_SC_HVL__EINVP_1%A N_A_M1003_g N_A_M1000_g A A A N_A_c_140_n
+ N_A_c_141_n A PM_SKY130_FD_SC_HVL__EINVP_1%A
x_PM_SKY130_FD_SC_HVL__EINVP_1%VPWR N_VPWR_M1002_d VPWR N_VPWR_c_177_n
+ N_VPWR_c_180_n PM_SKY130_FD_SC_HVL__EINVP_1%VPWR
x_PM_SKY130_FD_SC_HVL__EINVP_1%Z N_Z_M1003_d N_Z_M1000_d N_Z_c_203_n Z Z Z Z Z Z
+ Z N_Z_c_201_n Z PM_SKY130_FD_SC_HVL__EINVP_1%Z
x_PM_SKY130_FD_SC_HVL__EINVP_1%VGND N_VGND_M1005_d VGND N_VGND_c_224_n
+ N_VGND_c_226_n PM_SKY130_FD_SC_HVL__EINVP_1%VGND
cc_1 N_VNB_M1005_b N_TE_M1005_g 0.0623383f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=1.155
cc_2 N_VNB_M1005_b N_TE_c_52_n 0.0978212f $X=-0.33 $Y=-0.265 $X2=1.565 $Y2=0.322
cc_3 N_VNB_M1005_b N_TE_c_53_n 0.0960056f $X=-0.33 $Y=-0.265 $X2=0.935 $Y2=0.322
cc_4 N_VNB_c_4_p N_TE_c_53_n 0.0318307f $X=0.24 $Y=0 $X2=0.935 $Y2=0.322
cc_5 N_VNB_M1005_b N_TE_c_55_n 0.0347561f $X=-0.33 $Y=-0.265 $X2=1.815 $Y2=0.505
cc_6 N_VNB_M1005_b TE 0.0107085f $X=-0.33 $Y=-0.265 $X2=1.115 $Y2=1.58
cc_7 N_VNB_M1005_b N_TE_c_57_n 0.0564291f $X=-0.33 $Y=-0.265 $X2=1.02 $Y2=1.66
cc_8 N_VNB_M1005_b N_A_30_189#_c_89_n 0.00484338f $X=-0.33 $Y=-0.265 $X2=0.935
+ $Y2=0.322
cc_9 N_VNB_M1005_b N_A_30_189#_c_90_n 0.0244824f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.58
cc_10 N_VNB_M1005_b N_A_30_189#_c_91_n 0.00105941f $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=1.627
cc_11 N_VNB_M1005_b N_A_30_189#_c_92_n 0.0311759f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_12 N_VNB_M1005_b N_A_M1003_g 0.0622464f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=1.155
cc_13 N_VNB_c_4_p N_A_M1003_g 5.31052e-19 $X=0.24 $Y=0 $X2=0.685 $Y2=1.155
cc_14 N_VNB_M1005_b N_A_c_140_n 0.0351119f $X=-0.33 $Y=-0.265 $X2=1.02 $Y2=1.66
cc_15 N_VNB_M1005_b N_A_c_141_n 0.00446334f $X=-0.33 $Y=-0.265 $X2=0.81
+ $Y2=1.495
cc_16 N_VNB_M1005_b Z 0.00675384f $X=-0.33 $Y=-0.265 $X2=1.815 $Y2=0.505
cc_17 N_VNB_M1005_b Z 0.0206333f $X=-0.33 $Y=-0.265 $X2=1.815 $Y2=0.99
cc_18 N_VNB_M1005_b N_Z_c_201_n 0.0347331f $X=-0.33 $Y=-0.265 $X2=1.2 $Y2=1.627
cc_19 N_VNB_c_4_p N_Z_c_201_n 5.30181e-19 $X=0.24 $Y=0 $X2=1.2 $Y2=1.627
cc_20 N_VNB_M1005_b N_VGND_c_224_n 0.0727262f $X=-0.33 $Y=-0.265 $X2=0.935
+ $Y2=0.322
cc_21 N_VNB_c_4_p N_VGND_c_224_n 0.356645f $X=0.24 $Y=0 $X2=0.935 $Y2=0.322
cc_22 N_VNB_M1005_b N_VGND_c_226_n 0.101378f $X=-0.33 $Y=-0.265 $X2=1.815
+ $Y2=0.99
cc_23 N_VNB_c_4_p N_VGND_c_226_n 0.00963021f $X=0.24 $Y=0 $X2=1.815 $Y2=0.99
cc_24 N_VPB_M1002_b N_TE_M1002_g 0.043558f $X=-0.33 $Y=1.885 $X2=0.935 $Y2=2.59
cc_25 N_VPB_M1002_b N_TE_c_57_n 0.0309129f $X=-0.33 $Y=1.885 $X2=1.02 $Y2=1.66
cc_26 N_VPB_M1002_b N_A_30_189#_c_90_n 0.00204435f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_27 N_VPB_M1002_b N_A_30_189#_c_94_n 0.0519052f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_28 N_VPB_M1002_b N_A_30_189#_c_91_n 0.00176715f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=1.627
cc_29 N_VPB_M1002_b N_A_30_189#_c_96_n 0.0101855f $X=-0.33 $Y=1.885 $X2=1.2
+ $Y2=1.627
cc_30 N_VPB_M1002_b N_A_30_189#_c_92_n 0.0256162f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_31 N_VPB_M1002_b N_A_30_189#_c_98_n 0.00567684f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_32 N_VPB_M1002_b N_A_30_189#_c_99_n 0.0376268f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_33 VPB N_A_30_189#_c_99_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_34 N_VPB_c_34_p N_A_30_189#_c_99_n 0.0137101f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_35 N_VPB_M1002_b N_A_M1000_g 0.0529589f $X=-0.33 $Y=1.885 $X2=0.935 $Y2=2.59
cc_36 VPB N_A_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.935 $Y2=2.59
cc_37 N_VPB_c_34_p N_A_M1000_g 0.0152014f $X=3.12 $Y=4.07 $X2=0.935 $Y2=2.59
cc_38 N_VPB_M1002_b N_A_c_140_n 0.0161067f $X=-0.33 $Y=1.885 $X2=1.02 $Y2=1.66
cc_39 N_VPB_M1002_b N_A_c_141_n 4.59744e-19 $X=-0.33 $Y=1.885 $X2=0.81 $Y2=1.495
cc_40 N_VPB_M1002_b N_VPWR_c_177_n 0.0313023f $X=-0.33 $Y=1.885 $X2=1.815
+ $Y2=0.505
cc_41 VPB N_VPWR_c_177_n 0.00755533f $X=0 $Y=3.955 $X2=1.815 $Y2=0.505
cc_42 N_VPB_c_34_p N_VPWR_c_177_n 0.100637f $X=3.12 $Y=4.07 $X2=1.815 $Y2=0.505
cc_43 N_VPB_M1002_b N_VPWR_c_180_n 0.0658688f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_44 VPB N_VPWR_c_180_n 0.357555f $X=0 $Y=3.955 $X2=0.635 $Y2=1.58
cc_45 N_VPB_c_34_p N_VPWR_c_180_n 0.0163443f $X=3.12 $Y=4.07 $X2=0.635 $Y2=1.58
cc_46 N_VPB_M1002_b N_Z_c_203_n 0.00675384f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_47 N_VPB_M1002_b Z 0.0115365f $X=-0.33 $Y=1.885 $X2=1.815 $Y2=0.99
cc_48 N_VPB_M1002_b Z 0.0499659f $X=-0.33 $Y=1.885 $X2=0.635 $Y2=1.58
cc_49 VPB Z 7.75439e-19 $X=0 $Y=3.955 $X2=0.635 $Y2=1.58
cc_50 N_VPB_c_34_p Z 0.0133691f $X=3.12 $Y=4.07 $X2=0.635 $Y2=1.58
cc_51 N_TE_M1005_g N_A_30_189#_c_89_n 0.00149905f $X=0.685 $Y=1.155 $X2=0.24
+ $Y2=0
cc_52 N_TE_M1005_g N_A_30_189#_c_90_n 0.0223933f $X=0.685 $Y=1.155 $X2=0 $Y2=0
cc_53 TE N_A_30_189#_c_90_n 0.0194177f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_54 N_TE_M1002_g N_A_30_189#_c_94_n 0.00985499f $X=0.935 $Y=2.59 $X2=3.12
+ $Y2=0
cc_55 N_TE_c_55_n N_A_30_189#_c_106_n 0.00214431f $X=1.815 $Y=0.505 $X2=1.68
+ $Y2=0
cc_56 TE N_A_30_189#_c_106_n 0.00202953f $X=1.115 $Y=1.58 $X2=1.68 $Y2=0
cc_57 N_TE_c_57_n N_A_30_189#_c_106_n 0.00117054f $X=1.02 $Y=1.66 $X2=1.68 $Y2=0
cc_58 TE N_A_30_189#_c_96_n 0.0100739f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_59 N_TE_c_57_n N_A_30_189#_c_96_n 0.0177305f $X=1.02 $Y=1.66 $X2=0 $Y2=0
cc_60 N_TE_c_55_n N_A_30_189#_c_92_n 0.0354262f $X=1.815 $Y=0.505 $X2=0 $Y2=0
cc_61 TE N_A_30_189#_c_92_n 8.23844e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_62 N_TE_c_57_n N_A_30_189#_c_92_n 0.0282711f $X=1.02 $Y=1.66 $X2=0 $Y2=0
cc_63 N_TE_M1002_g N_A_30_189#_c_98_n 0.0124279f $X=0.935 $Y=2.59 $X2=0 $Y2=0
cc_64 TE N_A_30_189#_c_98_n 0.0445331f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_65 N_TE_c_57_n N_A_30_189#_c_98_n 0.0171643f $X=1.02 $Y=1.66 $X2=0 $Y2=0
cc_66 N_TE_M1002_g N_A_30_189#_c_99_n 0.0194804f $X=0.935 $Y=2.59 $X2=0 $Y2=0
cc_67 N_TE_c_52_n N_A_M1003_g 0.0338424f $X=1.565 $Y=0.322 $X2=0 $Y2=0
cc_68 N_TE_c_55_n A 0.00120775f $X=1.815 $Y=0.505 $X2=0 $Y2=0
cc_69 N_TE_M1002_g N_VPWR_c_177_n 0.0639217f $X=0.935 $Y=2.59 $X2=0.24 $Y2=0
cc_70 N_TE_M1002_g N_VPWR_c_180_n 0.00411177f $X=0.935 $Y=2.59 $X2=0 $Y2=0
cc_71 N_TE_M1005_g N_VGND_c_224_n 0.00318443f $X=0.685 $Y=1.155 $X2=0.24 $Y2=0
cc_72 N_TE_c_52_n N_VGND_c_224_n 0.0055897f $X=1.565 $Y=0.322 $X2=0.24 $Y2=0
cc_73 N_TE_c_53_n N_VGND_c_224_n 0.00504778f $X=0.935 $Y=0.322 $X2=0.24 $Y2=0
cc_74 N_TE_M1005_g N_VGND_c_226_n 0.066552f $X=0.685 $Y=1.155 $X2=0 $Y2=0
cc_75 N_TE_c_52_n N_VGND_c_226_n 0.0399241f $X=1.565 $Y=0.322 $X2=0 $Y2=0
cc_76 N_TE_c_53_n N_VGND_c_226_n 0.0129581f $X=0.935 $Y=0.322 $X2=0 $Y2=0
cc_77 N_TE_c_55_n N_VGND_c_226_n 0.0610847f $X=1.815 $Y=0.505 $X2=0 $Y2=0
cc_78 TE N_VGND_c_226_n 0.0578908f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_79 N_TE_c_57_n N_VGND_c_226_n 0.00671392f $X=1.02 $Y=1.66 $X2=0 $Y2=0
cc_80 N_A_30_189#_c_91_n N_A_M1000_g 6.47017e-19 $X=1.9 $Y=1.89 $X2=0 $Y2=0
cc_81 N_A_30_189#_c_92_n N_A_M1000_g 0.0635658f $X=1.56 $Y=1.89 $X2=0 $Y2=0
cc_82 N_A_30_189#_c_91_n N_A_c_140_n 2.83739e-19 $X=1.9 $Y=1.89 $X2=0 $Y2=0
cc_83 N_A_30_189#_c_92_n N_A_c_140_n 0.0163745f $X=1.56 $Y=1.89 $X2=0 $Y2=0
cc_84 N_A_30_189#_c_91_n N_A_c_141_n 0.0159389f $X=1.9 $Y=1.89 $X2=1.68 $Y2=0
cc_85 N_A_30_189#_c_92_n N_A_c_141_n 4.43227e-19 $X=1.56 $Y=1.89 $X2=1.68 $Y2=0
cc_86 N_A_30_189#_c_91_n A 0.00602813f $X=1.9 $Y=1.89 $X2=0 $Y2=0
cc_87 N_A_30_189#_c_92_n A 0.00136166f $X=1.56 $Y=1.89 $X2=0 $Y2=0
cc_88 N_A_30_189#_c_99_n A 2.31883e-19 $X=1.73 $Y=2.105 $X2=0 $Y2=0
cc_89 N_A_30_189#_c_94_n N_VPWR_c_177_n 0.0308168f $X=0.545 $Y=2.34 $X2=0.24
+ $Y2=0
cc_90 N_A_30_189#_c_92_n N_VPWR_c_177_n 0.00393677f $X=1.56 $Y=1.89 $X2=0.24
+ $Y2=0
cc_91 N_A_30_189#_c_98_n N_VPWR_c_177_n 0.089152f $X=1.475 $Y=1.912 $X2=0.24
+ $Y2=0
cc_92 N_A_30_189#_c_99_n N_VPWR_c_177_n 0.100625f $X=1.73 $Y=2.105 $X2=0.24
+ $Y2=0
cc_93 N_A_30_189#_c_94_n N_VPWR_c_180_n 0.0208897f $X=0.545 $Y=2.34 $X2=0 $Y2=0
cc_94 N_A_30_189#_c_99_n N_VPWR_c_180_n 0.00265054f $X=1.73 $Y=2.105 $X2=0 $Y2=0
cc_95 N_A_30_189#_c_89_n N_VGND_c_224_n 0.0103574f $X=0.277 $Y=1.233 $X2=0.24
+ $Y2=0
cc_96 N_A_30_189#_c_89_n N_VGND_c_226_n 0.0196294f $X=0.277 $Y=1.233 $X2=0 $Y2=0
cc_97 N_A_30_189#_c_106_n N_VGND_c_226_n 0.0231198f $X=1.662 $Y=1.912 $X2=0
+ $Y2=0
cc_98 N_A_30_189#_c_92_n N_VGND_c_226_n 0.00515043f $X=1.56 $Y=1.89 $X2=0 $Y2=0
cc_99 N_A_30_189#_c_98_n N_VGND_c_226_n 0.00535328f $X=1.475 $Y=1.912 $X2=0
+ $Y2=0
cc_100 N_A_M1000_g N_VPWR_c_177_n 0.0753079f $X=2.675 $Y=2.965 $X2=0.24 $Y2=0
cc_101 A N_VPWR_c_177_n 0.0512505f $X=2.64 $Y=2.035 $X2=0.24 $Y2=0
cc_102 N_A_M1000_g N_VPWR_c_180_n 0.00858613f $X=2.675 $Y=2.965 $X2=0 $Y2=0
cc_103 N_A_M1000_g N_Z_c_203_n 0.0057757f $X=2.675 $Y=2.965 $X2=0 $Y2=0
cc_104 A N_Z_c_203_n 0.0193751f $X=2.64 $Y=2.035 $X2=0 $Y2=0
cc_105 A Z 0.0148024f $X=2.555 $Y=1.21 $X2=0.24 $Y2=0
cc_106 N_A_M1003_g Z 0.00457212f $X=2.675 $Y=0.99 $X2=0 $Y2=0
cc_107 N_A_M1000_g Z 0.00457212f $X=2.675 $Y=2.965 $X2=0 $Y2=0
cc_108 A Z 0.0105027f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_109 N_A_c_140_n Z 0.00947198f $X=2.78 $Y=1.79 $X2=0 $Y2=0
cc_110 N_A_c_141_n Z 0.0262246f $X=2.78 $Y=1.79 $X2=0 $Y2=0
cc_111 A Z 0.0105027f $X=2.64 $Y=2.035 $X2=0 $Y2=0
cc_112 N_A_M1003_g N_Z_c_201_n 0.0061935f $X=2.675 $Y=0.99 $X2=0 $Y2=0
cc_113 N_A_M1003_g N_VGND_c_224_n 0.00852558f $X=2.675 $Y=0.99 $X2=0.24 $Y2=0
cc_114 A N_VGND_c_224_n 0.00153036f $X=2.555 $Y=1.21 $X2=0.24 $Y2=0
cc_115 N_A_M1003_g N_VGND_c_226_n 0.049015f $X=2.675 $Y=0.99 $X2=0 $Y2=0
cc_116 A N_VGND_c_226_n 0.0426319f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_117 N_A_c_140_n N_VGND_c_226_n 0.00226959f $X=2.78 $Y=1.79 $X2=0 $Y2=0
cc_118 N_A_c_141_n N_VGND_c_226_n 0.00396758f $X=2.78 $Y=1.79 $X2=0 $Y2=0
cc_119 N_VPWR_c_177_n A_413_443# 0.0159386f $X=0.915 $Y=3.59 $X2=0 $Y2=3.985
cc_120 N_VPWR_c_180_n N_Z_M1000_d 0.00221032f $X=2.715 $Y=3.59 $X2=0 $Y2=0
cc_121 N_VPWR_c_177_n Z 0.0450946f $X=0.915 $Y=3.59 $X2=3.12 $Y2=4.07
cc_122 N_VPWR_c_180_n Z 0.0358369f $X=2.715 $Y=3.59 $X2=3.12 $Y2=4.07
cc_123 N_Z_M1003_d N_VGND_c_224_n 0.00221032f $X=2.925 $Y=0.615 $X2=0.24 $Y2=0
cc_124 N_Z_c_201_n N_VGND_c_224_n 0.0224844f $X=3.065 $Y=0.74 $X2=0.24 $Y2=0
cc_125 N_Z_c_201_n N_VGND_c_226_n 0.017742f $X=3.065 $Y=0.74 $X2=0 $Y2=0
cc_126 N_VGND_c_226_n A_413_123# 0.0126427f $X=1.425 $Y=0.74 $X2=0 $Y2=0
