* File: sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1.pex.spice
* Created: Fri Aug 28 09:37:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%VNB 9 11 12 17 43 46
r87 12 29 0.000656703 $w=1.104e-05 $l=5.8e-08 $layer=MET1_cond $X=5.52 $Y=8.082
+ $X2=5.52 $Y2=8.14
r88 12 46 2.26449e-05 $w=1.104e-05 $l=2e-09 $layer=MET1_cond $X=5.52 $Y=8.082
+ $X2=5.52 $Y2=8.08
r89 11 43 3.39674e-05 $w=1.104e-05 $l=3e-09 $layer=MET1_cond $X=5.52 $Y=0.057
+ $X2=5.52 $Y2=0.06
r90 11 17 0.00064538 $w=1.104e-05 $l=5.7e-08 $layer=MET1_cond $X=5.52 $Y=0.057
+ $X2=5.52 $Y2=0
r91 9 29 0.808696 $w=1.7e-07 $l=1.955e-06 $layer=mcon $count=11 $X=10.8 $Y=8.14
+ $X2=10.8 $Y2=8.14
r92 9 29 0.808696 $w=1.7e-07 $l=1.955e-06 $layer=mcon $count=11 $X=0.24 $Y=8.14
+ $X2=0.24 $Y2=8.14
r93 9 17 0.808696 $w=1.7e-07 $l=1.955e-06 $layer=mcon $count=11 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r94 9 17 0.808696 $w=1.7e-07 $l=1.955e-06 $layer=mcon $count=11 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%VPB 10 11 14 17 29 30
c83 30 0 1.93214e-19 $X=10.8 $Y=4.07
r84 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=4.07
+ $X2=10.8 $Y2=4.07
r85 27 29 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.88 $Y=4.07
+ $X2=10.8 $Y2=4.07
r86 24 30 1.53985 $w=2.3e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=4.07 $X2=10.8
+ $Y2=4.07
r87 23 27 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=4.07 $X2=8.88
+ $Y2=4.07
r88 23 24 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=4.07 $X2=8.4
+ $Y2=4.07
r89 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r90 14 24 1.84782 $w=2.3e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=4.07
+ $X2=8.4 $Y2=4.07
r91 14 18 3.38767 $w=2.3e-07 $l=5.28e-06 $layer=MET1_cond $X=5.52 $Y=4.07
+ $X2=0.24 $Y2=4.07
r92 11 29 182 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=1
+ $X=10.56 $Y=3.985 $X2=10.8 $Y2=4.07
r93 11 27 91 $w=1.7e-07 $l=7.26258e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=8.195 $Y=3.985 $X2=8.88 $Y2=4.07
r94 10 17 182 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=1 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%LVPWR 1 7 11 13 19
r55 19 22 4.74802 $w=7.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.73 $Y=3.19
+ $X2=3.73 $Y2=3.485
r56 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.93 $Y=3.19
+ $X2=3.93 $Y2=3.19
r57 17 20 0.179425 $w=2.85e-07 $l=3.6e-07 $layer=MET1_cond $X=3.57 $Y=3.162
+ $X2=3.93 $Y2=3.162
r58 16 19 0.885224 $w=7.58e-07 $l=5.5e-08 $layer=LI1_cond $X=3.73 $Y=3.135
+ $X2=3.73 $Y2=3.19
r59 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.57 $Y=3.135
+ $X2=3.57 $Y2=3.135
r60 13 20 0.792462 $w=2.85e-07 $l=1.59e-06 $layer=MET1_cond $X=5.52 $Y=3.162
+ $X2=3.93 $Y2=3.162
r61 9 16 6.31558 $w=7.58e-07 $l=1.87617e-07 $layer=LI1_cond $X=3.57 $Y=3.075
+ $X2=3.73 $Y2=3.135
r62 9 11 31.7989 $w=2.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.57 $Y=3.075
+ $X2=3.57 $Y2=2.33
r63 7 22 45.5 $w=1.7e-07 $l=7.69756e-07 $layer=licon1_NTAP_notbjt $count=4
+ $X=3.265 $Y=3.305 $X2=3.95 $Y2=3.485
r64 1 11 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=3.43
+ $Y=2.195 $X2=3.57 $Y2=2.33
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A 1 3 5 8 10 11 12 16
r32 16 19 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.66 $Y=1.695
+ $X2=2.66 $Y2=1.87
r33 11 12 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.65 $Y=1.665
+ $X2=2.65 $Y2=2.035
r34 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.66
+ $Y=1.695 $X2=2.66 $Y2=1.695
r35 6 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=2.035
+ $X2=3.355 $Y2=1.87
r36 6 8 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.355 $Y=2.035
+ $X2=3.355 $Y2=2.615
r37 3 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.705
+ $X2=3.355 $Y2=1.87
r38 3 5 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.355 $Y=1.705
+ $X2=3.355 $Y2=1.175
r39 2 19 2.83073 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.825 $Y=1.87
+ $X2=2.66 $Y2=1.87
r40 1 10 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.28 $Y=1.87
+ $X2=3.355 $Y2=1.87
r41 1 2 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=3.28 $Y=1.87
+ $X2=2.825 $Y2=1.87
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_573_897# 1 2 7 8 9 11 12
+ 14 17 19 21 27 30 31 38 43 46 47 50 51
c82 31 0 1.93214e-19 $X=3.03 $Y=4.65
r83 49 50 8.79496 $w=3.78e-07 $l=2.9e-07 $layer=LI1_cond $X=3.075 $Y=2.765
+ $X2=3.075 $Y2=3.055
r84 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.145
+ $Y=1.87 $X2=4.145 $Y2=1.87
r85 44 51 1.88208 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=3.265 $Y=1.87
+ $X2=3.12 $Y2=1.87
r86 44 46 40.566 $w=2.48e-07 $l=8.8e-07 $layer=LI1_cond $X=3.265 $Y=1.87
+ $X2=4.145 $Y2=1.87
r87 43 49 17.2866 $w=2.88e-07 $l=4.35e-07 $layer=LI1_cond $X=3.12 $Y=2.33
+ $X2=3.12 $Y2=2.765
r88 40 51 4.55795 $w=2.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.12 $Y=1.995
+ $X2=3.12 $Y2=1.87
r89 40 43 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=3.12 $Y=1.995
+ $X2=3.12 $Y2=2.33
r90 36 51 4.55795 $w=2.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.12 $Y=1.745
+ $X2=3.12 $Y2=1.87
r91 36 38 33.5798 $w=2.88e-07 $l=8.45e-07 $layer=LI1_cond $X=3.12 $Y=1.745
+ $X2=3.12 $Y2=0.9
r92 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.03
+ $Y=5.33 $X2=3.03 $Y2=5.33
r93 31 34 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=3.03 $Y=4.65
+ $X2=3.03 $Y2=5.33
r94 30 33 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=3.03 $Y=4.65
+ $X2=3.03 $Y2=5.33
r95 30 50 63.3844 $w=2.88e-07 $l=1.595e-06 $layer=LI1_cond $X=3.03 $Y=4.65
+ $X2=3.03 $Y2=3.055
r96 30 31 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.03
+ $Y=4.65 $X2=3.03 $Y2=4.65
r97 26 47 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=3.86 $Y=1.87
+ $X2=4.145 $Y2=1.87
r98 26 27 5.03009 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.86 $Y=1.87
+ $X2=3.75 $Y2=1.87
r99 22 34 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=3.03 $Y=5.665
+ $X2=3.03 $Y2=5.33
r100 19 21 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.61 $Y=5.995 $X2=4.61
+ $Y2=6.855
r101 15 27 37.0704 $w=1.5e-07 $l=1.81659e-07 $layer=POLY_cond $X=3.785 $Y=2.035
+ $X2=3.75 $Y2=1.87
r102 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.785 $Y=2.035
+ $X2=3.785 $Y2=2.615
r103 12 27 37.0704 $w=1.5e-07 $l=1.81659e-07 $layer=POLY_cond $X=3.785 $Y=1.705
+ $X2=3.75 $Y2=1.87
r104 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.785 $Y=1.705
+ $X2=3.785 $Y2=1.175
r105 9 19 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=3.83 $Y=5.83
+ $X2=4.61 $Y2=5.83
r106 9 11 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.83 $Y=5.995 $X2=3.83
+ $Y2=6.855
r107 8 22 26.9307 $w=3.3e-07 $l=2.33345e-07 $layer=POLY_cond $X=3.195 $Y=5.83
+ $X2=3.03 $Y2=5.665
r108 7 9 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.58 $Y=5.83 $X2=3.83
+ $Y2=5.83
r109 7 8 67.3216 $w=3.3e-07 $l=3.85e-07 $layer=POLY_cond $X=3.58 $Y=5.83
+ $X2=3.195 $Y2=5.83
r110 2 43 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=2.195 $X2=3.14 $Y2=2.33
r111 1 38 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=2.985
+ $Y=0.755 $X2=3.14 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_772_151# 1 2 7 9 10 12 15
+ 20 21 26 31 35 37
r50 35 36 23.6688 $w=3.17e-07 $l=6.15e-07 $layer=LI1_cond $X=4.03 $Y=2.31
+ $X2=4.645 $Y2=2.31
r51 34 35 1.15457 $w=3.17e-07 $l=3e-08 $layer=LI1_cond $X=4 $Y=2.31 $X2=4.03
+ $Y2=2.31
r52 29 31 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=4.03 $Y=1.41
+ $X2=4.645 $Y2=1.41
r53 27 37 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.625 $Y=2.31
+ $X2=5.485 $Y2=2.31
r54 26 27 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.625
+ $Y=2.31 $X2=5.625 $Y2=2.31
r55 24 37 94.4251 $w=3.3e-07 $l=5.4e-07 $layer=POLY_cond $X=4.945 $Y=2.31
+ $X2=5.485 $Y2=2.31
r56 23 26 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.945 $Y=2.31
+ $X2=5.625 $Y2=2.31
r57 23 24 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.945
+ $Y=2.31 $X2=4.945 $Y2=2.31
r58 21 36 6.1 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.81 $Y=2.31 $X2=4.645
+ $Y2=2.31
r59 21 23 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=4.81 $Y=2.31
+ $X2=4.945 $Y2=2.31
r60 20 36 0.469914 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=2.145
+ $X2=4.645 $Y2=2.31
r61 19 31 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=1.575
+ $X2=4.645 $Y2=1.41
r62 19 20 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=4.645 $Y=1.575
+ $X2=4.645 $Y2=2.145
r63 13 29 1.09485 $w=3.1e-07 $l=1.65e-07 $layer=LI1_cond $X=4.03 $Y=1.245
+ $X2=4.03 $Y2=1.41
r64 13 15 12.8256 $w=3.08e-07 $l=3.45e-07 $layer=LI1_cond $X=4.03 $Y=1.245
+ $X2=4.03 $Y2=0.9
r65 10 12 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.515 $Y=2.145
+ $X2=6.515 $Y2=1.285
r66 7 10 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=5.735 $Y=2.31
+ $X2=6.515 $Y2=2.31
r67 7 27 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=5.735 $Y=2.31
+ $X2=5.625 $Y2=2.31
r68 7 9 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.735 $Y=2.145 $X2=5.735
+ $Y2=1.285
r69 2 34 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=3.86
+ $Y=2.195 $X2=4 $Y2=2.33
r70 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.86
+ $Y=0.755 $X2=4 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_1400_777# 1 2 10 12 14 21
+ 22 24 25 26 28
r70 28 31 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=8.465 $Y=0.68
+ $X2=8.465 $Y2=1.89
r71 26 34 23.7599 $w=6.29e-07 $l=1.44733e-06 $layer=LI1_cond $X=8.465 $Y=2.495
+ $X2=9.69 $Y2=2.98
r72 26 31 12.2649 $w=5.88e-07 $l=6.05e-07 $layer=LI1_cond $X=8.465 $Y=2.495
+ $X2=8.465 $Y2=1.89
r73 24 26 11.5337 $w=6.29e-07 $l=3.43511e-07 $layer=LI1_cond $X=8.17 $Y=2.6
+ $X2=8.465 $Y2=2.495
r74 24 25 21.3896 $w=2.08e-07 $l=4.05e-07 $layer=LI1_cond $X=8.17 $Y=2.6
+ $X2=7.765 $Y2=2.6
r75 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.6 $Y=4.05
+ $X2=7.6 $Y2=4.05
r76 19 25 9.58248 $w=2.1e-07 $l=3.83927e-07 $layer=LI1_cond $X=7.43 $Y=2.705
+ $X2=7.765 $Y2=2.6
r77 19 21 24.0108 $w=6.68e-07 $l=1.345e-06 $layer=LI1_cond $X=7.43 $Y=2.705
+ $X2=7.43 $Y2=4.05
r78 12 14 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=8.075 $Y=6.055
+ $X2=8.075 $Y2=5.175
r79 11 22 54.642 $w=4.19e-07 $l=4.75e-07 $layer=POLY_cond $X=8.075 $Y=4.117
+ $X2=7.6 $Y2=4.117
r80 11 14 88.2799 $w=5e-07 $l=8.25e-07 $layer=POLY_cond $X=8.075 $Y=4.35
+ $X2=8.075 $Y2=5.175
r81 8 12 144.261 $w=3.3e-07 $l=8.25e-07 $layer=POLY_cond $X=7.25 $Y=6.22
+ $X2=8.075 $Y2=6.22
r82 8 10 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=7.25 $Y=6.055 $X2=7.25
+ $Y2=5.175
r83 7 22 40.2625 $w=4.19e-07 $l=3.5e-07 $layer=POLY_cond $X=7.25 $Y=4.117
+ $X2=7.6 $Y2=4.117
r84 7 10 88.2799 $w=5e-07 $l=8.25e-07 $layer=POLY_cond $X=7.25 $Y=4.35 $X2=7.25
+ $Y2=5.175
r85 2 34 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=9.47
+ $Y=2.815 $X2=9.69 $Y2=2.96
r86 1 31 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=8.325
+ $Y=0.535 $X2=8.465 $Y2=1.89
r87 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.325
+ $Y=0.535 $X2=8.465 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_816_1221# 1 2 3 4 15 19 22
+ 24 25 27 29 31 32 36 40 41 44 47 49 50 51 54 61 65 67 68
c109 29 0 1.38777e-20 $X=8.97 $Y=3.025
c110 24 0 1.38892e-19 $X=9.51 $Y=6.285
r111 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.7
+ $Y=6.45 $X2=8.7 $Y2=6.45
r112 61 63 5.26418 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.795 $Y=4.57
+ $X2=6.795 $Y2=4.735
r113 61 62 5.26418 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.795 $Y=4.57
+ $X2=6.795 $Y2=4.405
r114 54 57 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=8.465 $Y=4.57
+ $X2=8.465 $Y2=5.78
r115 52 67 5.51329 $w=3.05e-07 $l=2.05925e-07 $layer=LI1_cond $X=8.465 $Y=6.285
+ $X2=8.557 $Y2=6.45
r116 52 57 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=8.465 $Y=6.285
+ $X2=8.465 $Y2=5.78
r117 50 67 1.06046 $w=3.3e-07 $l=2.57e-07 $layer=LI1_cond $X=8.3 $Y=6.45
+ $X2=8.557 $Y2=6.45
r118 50 51 44.5262 $w=3.28e-07 $l=1.275e-06 $layer=LI1_cond $X=8.3 $Y=6.45
+ $X2=7.025 $Y2=6.45
r119 49 51 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=6.86 $Y=6.285
+ $X2=7.025 $Y2=6.45
r120 48 65 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.86 $Y=5.995
+ $X2=6.86 $Y2=5.83
r121 48 49 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=6.86 $Y=5.995
+ $X2=6.86 $Y2=6.285
r122 47 65 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.86 $Y=5.665
+ $X2=6.86 $Y2=5.83
r123 47 63 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=6.86 $Y=5.665
+ $X2=6.86 $Y2=4.735
r124 44 62 50.463 $w=3.28e-07 $l=1.445e-06 $layer=LI1_cond $X=6.73 $Y=2.96
+ $X2=6.73 $Y2=4.405
r125 40 65 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=5.83
+ $X2=6.86 $Y2=5.83
r126 40 41 80.671 $w=3.28e-07 $l=2.31e-06 $layer=LI1_cond $X=6.695 $Y=5.83
+ $X2=4.385 $Y2=5.83
r127 36 38 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=4.22 $Y=6.25
+ $X2=4.22 $Y2=7.46
r128 34 41 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=4.22 $Y=5.995
+ $X2=4.385 $Y2=5.83
r129 34 36 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.22 $Y=5.995
+ $X2=4.22 $Y2=6.25
r130 29 30 19.4957 $w=1.162e-06 $l=4.7e-07 $layer=POLY_cond $X=8.97 $Y=3.307
+ $X2=9.44 $Y2=3.307
r131 25 33 51.2401 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=9.55 $Y=6.975
+ $X2=9.55 $Y2=6.45
r132 25 27 24.582 $w=5e-07 $l=2.55e-07 $layer=POLY_cond $X=9.55 $Y=6.975
+ $X2=9.55 $Y2=7.23
r133 24 33 18.0037 $w=4.48e-07 $l=1.83916e-07 $layer=POLY_cond $X=9.51 $Y=6.285
+ $X2=9.55 $Y2=6.45
r134 24 32 30.456 $w=4.2e-07 $l=2.3e-07 $layer=POLY_cond $X=9.51 $Y=6.285
+ $X2=9.51 $Y2=6.055
r135 20 32 28.2776 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=9.55 $Y=5.805
+ $X2=9.55 $Y2=6.055
r136 20 22 67.4137 $w=5e-07 $l=6.3e-07 $layer=POLY_cond $X=9.55 $Y=5.805
+ $X2=9.55 $Y2=5.175
r137 19 31 37.0268 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=9.55 $Y=4.535
+ $X2=9.55 $Y2=4.285
r138 19 22 68.4838 $w=5e-07 $l=6.4e-07 $layer=POLY_cond $X=9.55 $Y=4.535
+ $X2=9.55 $Y2=5.175
r139 17 30 37.0314 $w=2.8e-07 $l=6.23e-07 $layer=POLY_cond $X=9.44 $Y=3.93
+ $X2=9.44 $Y2=3.307
r140 17 31 76.0548 $w=2.8e-07 $l=3.55e-07 $layer=POLY_cond $X=9.44 $Y=3.93
+ $X2=9.44 $Y2=4.285
r141 16 68 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.865 $Y=6.45
+ $X2=8.7 $Y2=6.45
r142 15 33 9.99217 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=9.3 $Y=6.45
+ $X2=9.55 $Y2=6.45
r143 15 16 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=9.3 $Y=6.45
+ $X2=8.865 $Y2=6.45
r144 4 57 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=8.325
+ $Y=4.425 $X2=8.465 $Y2=5.78
r145 4 54 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.325
+ $Y=4.425 $X2=8.465 $Y2=4.57
r146 3 44 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=6.665
+ $Y=2.815 $X2=6.81 $Y2=2.96
r147 2 65 300 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_PDIFF $count=2 $X=6.735
+ $Y=4.425 $X2=6.86 $Y2=5.78
r148 2 61 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=6.735
+ $Y=4.425 $X2=6.86 $Y2=4.57
r149 1 38 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=4.08
+ $Y=6.105 $X2=4.22 $Y2=7.46
r150 1 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.08
+ $Y=6.105 $X2=4.22 $Y2=6.25
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_1406_429# 1 2 7 9 10 12 13
+ 14 16 18 22 25 28 33 39 43 44 46
c99 46 0 1.38892e-19 $X=9.16 $Y=6.39
c100 7 0 6.01901e-20 $X=8.075 $Y=2.145
r101 44 49 16.3371 $w=6.95e-07 $l=1.65e-07 $layer=POLY_cond $X=10.277 $Y=6.39
+ $X2=10.277 $Y2=6.555
r102 44 48 16.3371 $w=6.95e-07 $l=1.65e-07 $layer=POLY_cond $X=10.277 $Y=6.39
+ $X2=10.277 $Y2=6.225
r103 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.435
+ $Y=6.39 $X2=10.435 $Y2=6.39
r104 41 46 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.325 $Y=6.39
+ $X2=9.16 $Y2=6.39
r105 41 43 38.764 $w=3.28e-07 $l=1.11e-06 $layer=LI1_cond $X=9.325 $Y=6.39
+ $X2=10.435 $Y2=6.39
r106 37 46 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.16 $Y=6.555
+ $X2=9.16 $Y2=6.39
r107 37 39 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=9.16 $Y=6.555
+ $X2=9.16 $Y2=7
r108 33 36 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=9.16 $Y=4.57
+ $X2=9.16 $Y2=5.78
r109 31 46 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.16 $Y=6.225
+ $X2=9.16 $Y2=6.39
r110 31 36 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=9.16 $Y=6.225
+ $X2=9.16 $Y2=5.78
r111 25 49 72.229 $w=5e-07 $l=6.75e-07 $layer=POLY_cond $X=10.375 $Y=7.23
+ $X2=10.375 $Y2=6.555
r112 22 48 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=10.375 $Y=5.175
+ $X2=10.375 $Y2=6.225
r113 19 22 88.2799 $w=5e-07 $l=8.25e-07 $layer=POLY_cond $X=10.375 $Y=4.35
+ $X2=10.375 $Y2=5.175
r114 16 19 37.6298 $w=5.7e-07 $l=5.41941e-07 $layer=POLY_cond $X=10.16 $Y=3.905
+ $X2=10.375 $Y2=4.35
r115 16 18 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=10.16 $Y=3.905
+ $X2=10.16 $Y2=3.025
r116 15 18 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=10.16 $Y=2.475
+ $X2=10.16 $Y2=3.025
r117 13 15 28.4267 $w=3.3e-07 $l=3.22102e-07 $layer=POLY_cond $X=9.91 $Y=2.31
+ $X2=10.16 $Y2=2.475
r118 13 14 140.763 $w=3.3e-07 $l=8.05e-07 $layer=POLY_cond $X=9.91 $Y=2.31
+ $X2=9.105 $Y2=2.31
r119 10 14 31.5386 $w=7.58e-07 $l=3.22102e-07 $layer=POLY_cond $X=8.855 $Y=2.145
+ $X2=9.105 $Y2=2.31
r120 10 12 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.855 $Y=2.145
+ $X2=8.855 $Y2=1.285
r121 7 10 49.5989 $w=7.58e-07 $l=7.8e-07 $layer=POLY_cond $X=8.075 $Y=2.145
+ $X2=8.855 $Y2=2.145
r122 7 28 34.6557 $w=7.58e-07 $l=1.01143e-06 $layer=POLY_cond $X=8.075 $Y=2.145
+ $X2=7.53 $Y2=2.92
r123 7 9 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.075 $Y=2.145 $X2=8.075
+ $Y2=1.285
r124 2 36 300 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_PDIFF $count=2 $X=9.035
+ $Y=4.425 $X2=9.16 $Y2=5.78
r125 2 33 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=9.035
+ $Y=4.425 $X2=9.16 $Y2=4.57
r126 1 39 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=9.035
+ $Y=6.855 $X2=9.16 $Y2=7
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%VPWR 1 2 3 4 13 14 18 27 34
+ 38 43 47
r86 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.6 $Y=3.56
+ $X2=10.6 $Y2=3.56
r87 43 46 12.1635 $w=5.88e-07 $l=6e-07 $layer=LI1_cond $X=10.42 $Y=2.96
+ $X2=10.42 $Y2=3.56
r88 37 40 24.327 $w=5.88e-07 $l=1.2e-06 $layer=LI1_cond $X=9.985 $Y=4.58
+ $X2=9.985 $Y2=5.78
r89 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.165 $Y=4.58
+ $X2=10.165 $Y2=4.58
r90 34 37 0.202725 $w=5.88e-07 $l=1e-08 $layer=LI1_cond $X=9.985 $Y=4.57
+ $X2=9.985 $Y2=4.58
r91 31 47 0.833075 $w=3.7e-07 $l=2.17e-06 $layer=MET1_cond $X=8.43 $Y=3.63
+ $X2=10.6 $Y2=3.63
r92 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.43 $Y=3.56
+ $X2=8.43 $Y2=3.56
r93 27 30 12.1635 $w=5.88e-07 $l=6e-07 $layer=LI1_cond $X=8.25 $Y=2.96 $X2=8.25
+ $Y2=3.56
r94 22 38 0.882982 $w=3.7e-07 $l=2.3e-06 $layer=MET1_cond $X=7.865 $Y=4.51
+ $X2=10.165 $Y2=4.51
r95 21 24 24.327 $w=5.88e-07 $l=1.2e-06 $layer=LI1_cond $X=7.685 $Y=4.58
+ $X2=7.685 $Y2=5.78
r96 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.865 $Y=4.58
+ $X2=7.865 $Y2=4.58
r97 18 21 0.202725 $w=5.88e-07 $l=1e-08 $layer=LI1_cond $X=7.685 $Y=4.57
+ $X2=7.685 $Y2=4.58
r98 14 22 0.900258 $w=3.7e-07 $l=2.345e-06 $layer=MET1_cond $X=5.52 $Y=4.51
+ $X2=7.865 $Y2=4.51
r99 13 31 1.11716 $w=3.7e-07 $l=2.91e-06 $layer=MET1_cond $X=5.52 $Y=3.63
+ $X2=8.43 $Y2=3.63
r100 4 43 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=10.41
+ $Y=2.815 $X2=10.63 $Y2=2.96
r101 3 40 300 $w=1.7e-07 $l=1.44454e-06 $layer=licon1_PDIFF $count=2 $X=9.8
+ $Y=4.425 $X2=9.985 $Y2=5.78
r102 3 34 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=9.8
+ $Y=4.425 $X2=9.985 $Y2=4.57
r103 2 27 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=8.03
+ $Y=2.815 $X2=8.25 $Y2=2.96
r104 1 24 300 $w=1.7e-07 $l=1.44454e-06 $layer=licon1_PDIFF $count=2 $X=7.5
+ $Y=4.425 $X2=7.685 $Y2=5.78
r105 1 18 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=7.5
+ $Y=4.425 $X2=7.685 $Y2=4.57
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%X 1 2 7 8 9 10 11 21 31 45
r17 35 45 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=10.765 $Y=6.89
+ $X2=10.765 $Y2=6.845
r18 31 41 2.40092 $w=2.38e-07 $l=5e-08 $layer=LI1_cond $X=10.81 $Y=6.105
+ $X2=10.81 $Y2=6.055
r19 11 45 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=10.765 $Y=6.825
+ $X2=10.765 $Y2=6.845
r20 11 43 4.36998 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=10.765 $Y=6.825
+ $X2=10.765 $Y2=6.725
r21 11 38 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=10.765 $Y=6.91
+ $X2=10.765 $Y2=7
r22 11 35 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=10.765 $Y=6.91
+ $X2=10.765 $Y2=6.89
r23 10 43 12.0046 $w=2.38e-07 $l=2.5e-07 $layer=LI1_cond $X=10.81 $Y=6.475
+ $X2=10.81 $Y2=6.725
r24 9 41 1.50633 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=10.765 $Y=6.037
+ $X2=10.765 $Y2=6.055
r25 9 19 5.13361 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=10.765 $Y=6.037
+ $X2=10.765 $Y2=5.89
r26 9 10 16.9505 $w=2.38e-07 $l=3.53e-07 $layer=LI1_cond $X=10.81 $Y=6.122
+ $X2=10.81 $Y2=6.475
r27 9 31 0.816314 $w=2.38e-07 $l=1.7e-08 $layer=LI1_cond $X=10.81 $Y=6.122
+ $X2=10.81 $Y2=6.105
r28 8 19 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=10.765 $Y=5.735
+ $X2=10.765 $Y2=5.89
r29 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.765 $Y=5.365
+ $X2=10.765 $Y2=5.735
r30 7 21 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=10.765 $Y=5.365
+ $X2=10.765 $Y2=4.57
r31 2 8 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=10.625
+ $Y=4.425 $X2=10.765 $Y2=5.78
r32 2 21 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=10.625
+ $Y=4.425 $X2=10.765 $Y2=4.57
r33 1 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.625
+ $Y=6.855 $X2=10.765 $Y2=7
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%VGND 1 2 3 4 5 6 21 23 24 25
+ 26 31 32 35 41 50 54 62 70 71 78 82 85
c96 25 0 6.01901e-20 $X=6.61 $Y=0.34
r97 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.57 $Y=0.51
+ $X2=3.57 $Y2=0.51
r98 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.165 $Y=7.63
+ $X2=10.165 $Y2=7.63
r99 78 81 12.7717 $w=5.88e-07 $l=6.3e-07 $layer=LI1_cond $X=9.985 $Y=7 $X2=9.985
+ $Y2=7.63
r100 73 75 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=6.905 $Y=0.68
+ $X2=6.905 $Y2=1.89
r101 70 73 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=6.905 $Y=0.51
+ $X2=6.905 $Y2=0.68
r102 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.085 $Y=0.51
+ $X2=7.085 $Y2=0.51
r103 65 67 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=5.345 $Y=0.68
+ $X2=5.345 $Y2=1.89
r104 62 65 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=5.345 $Y=0.51
+ $X2=5.345 $Y2=0.68
r105 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.18 $Y=7.63
+ $X2=5.18 $Y2=7.63
r106 57 59 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=5 $Y=7.46 $X2=5
+ $Y2=7.63
r107 54 57 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=5 $Y=6.25 $X2=5
+ $Y2=7.46
r108 51 86 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=3.93 $Y=0.44
+ $X2=3.57 $Y2=0.44
r109 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.93 $Y=0.45
+ $X2=3.93 $Y2=0.45
r110 48 85 5.89082 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=3.705 $Y=0.45
+ $X2=3.57 $Y2=0.45
r111 48 50 11.2739 $w=2.28e-07 $l=2.25e-07 $layer=LI1_cond $X=3.705 $Y=0.45
+ $X2=3.93 $Y2=0.45
r112 47 60 0.598892 $w=3.7e-07 $l=1.56e-06 $layer=MET1_cond $X=3.62 $Y=7.7
+ $X2=5.18 $Y2=7.7
r113 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.62 $Y=7.63
+ $X2=3.62 $Y2=7.63
r114 44 46 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=3.44 $Y=7.46
+ $X2=3.44 $Y2=7.63
r115 41 44 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=3.44 $Y=6.25
+ $X2=3.44 $Y2=7.46
r116 38 86 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=3.21 $Y=0.44
+ $X2=3.57 $Y2=0.44
r117 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.21 $Y=0.45
+ $X2=3.21 $Y2=0.45
r118 35 85 5.89082 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=3.435 $Y=0.45
+ $X2=3.57 $Y2=0.45
r119 35 37 11.2739 $w=2.28e-07 $l=2.25e-07 $layer=LI1_cond $X=3.435 $Y=0.45
+ $X2=3.21 $Y2=0.45
r120 32 82 1.78324 $w=3.7e-07 $l=4.645e-06 $layer=MET1_cond $X=5.52 $Y=7.7
+ $X2=10.165 $Y2=7.7
r121 32 60 0.130528 $w=3.7e-07 $l=3.4e-07 $layer=MET1_cond $X=5.52 $Y=7.7
+ $X2=5.18 $Y2=7.7
r122 31 71 0.600812 $w=3.7e-07 $l=1.565e-06 $layer=MET1_cond $X=5.52 $Y=0.44
+ $X2=7.085 $Y2=0.44
r123 31 51 0.61041 $w=3.7e-07 $l=1.59e-06 $layer=MET1_cond $X=5.52 $Y=0.44
+ $X2=3.93 $Y2=0.44
r124 31 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.525 $Y=0.51
+ $X2=5.525 $Y2=0.51
r125 30 70 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=0.425
+ $X2=6.905 $Y2=0.51
r126 29 62 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=5.345 $Y=0.425
+ $X2=5.345 $Y2=0.51
r127 28 59 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=7.715 $X2=5
+ $Y2=7.63
r128 27 46 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=7.715
+ $X2=3.44 $Y2=7.63
r129 26 29 9.96617 $w=1.7e-07 $l=3.34813e-07 $layer=LI1_cond $X=5.64 $Y=0.34
+ $X2=5.345 $Y2=0.425
r130 25 30 9.96617 $w=1.7e-07 $l=3.34813e-07 $layer=LI1_cond $X=6.61 $Y=0.34
+ $X2=6.905 $Y2=0.425
r131 25 26 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=6.61 $Y=0.34
+ $X2=5.64 $Y2=0.34
r132 24 27 9.96617 $w=1.7e-07 $l=3.34813e-07 $layer=LI1_cond $X=3.735 $Y=7.8
+ $X2=3.44 $Y2=7.715
r133 23 28 9.96617 $w=1.7e-07 $l=3.34813e-07 $layer=LI1_cond $X=4.705 $Y=7.8
+ $X2=5 $Y2=7.715
r134 23 24 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=4.705 $Y=7.8
+ $X2=3.735 $Y2=7.8
r135 19 85 0.77205 $w=2.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.57 $Y=0.565
+ $X2=3.57 $Y2=0.45
r136 19 21 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.57 $Y=0.565
+ $X2=3.57 $Y2=0.88
r137 6 78 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=9.8
+ $Y=6.855 $X2=9.985 $Y2=7
r138 5 75 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.535 $X2=6.905 $Y2=1.89
r139 5 73 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.535 $X2=6.905 $Y2=0.68
r140 4 67 91 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.535 $X2=5.345 $Y2=1.89
r141 4 65 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.535 $X2=5.345 $Y2=0.68
r142 3 57 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=4.86
+ $Y=6.105 $X2=5 $Y2=7.46
r143 3 54 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.86
+ $Y=6.105 $X2=5 $Y2=6.25
r144 2 21 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.43
+ $Y=0.755 $X2=3.57 $Y2=0.88
r145 1 44 91 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_NDIFF $count=2 $X=3.315
+ $Y=6.105 $X2=3.44 $Y2=7.46
r146 1 41 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=3.315
+ $Y=6.105 $X2=3.44 $Y2=6.25
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_SYMMETRIC_1%A_1197_107# 1 2 3 12 16 17
+ 21 24 25 28
c38 28 0 1.38777e-20 $X=9.245 $Y=0.68
r39 28 30 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=9.245 $Y=0.68
+ $X2=9.245 $Y2=1.89
r40 26 28 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=9.245 $Y=0.425
+ $X2=9.245 $Y2=0.68
r41 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.08 $Y=0.34
+ $X2=9.245 $Y2=0.425
r42 24 25 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=9.08 $Y=0.34
+ $X2=7.85 $Y2=0.34
r43 21 23 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=7.685 $Y=0.68
+ $X2=7.685 $Y2=1.89
r44 19 23 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.685 $Y=2.145
+ $X2=7.685 $Y2=1.89
r45 18 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.685 $Y=0.425
+ $X2=7.85 $Y2=0.34
r46 18 21 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.685 $Y=0.425
+ $X2=7.685 $Y2=0.68
r47 16 19 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=7.52 $Y=2.235
+ $X2=7.685 $Y2=2.145
r48 16 17 75.7879 $w=1.78e-07 $l=1.23e-06 $layer=LI1_cond $X=7.52 $Y=2.235
+ $X2=6.29 $Y2=2.235
r49 12 15 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=6.125 $Y=0.68
+ $X2=6.125 $Y2=1.89
r50 10 17 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=6.125 $Y=2.145
+ $X2=6.29 $Y2=2.235
r51 10 15 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.125 $Y=2.145
+ $X2=6.125 $Y2=1.89
r52 3 30 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=9.105
+ $Y=0.535 $X2=9.245 $Y2=1.89
r53 3 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.105
+ $Y=0.535 $X2=9.245 $Y2=0.68
r54 2 23 91 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_NDIFF $count=2 $X=7.56
+ $Y=0.535 $X2=7.685 $Y2=1.89
r55 2 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=7.56
+ $Y=0.535 $X2=7.685 $Y2=0.68
r56 1 15 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=5.985
+ $Y=0.535 $X2=6.125 $Y2=1.89
r57 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.985
+ $Y=0.535 $X2=6.125 $Y2=0.68
.ends

