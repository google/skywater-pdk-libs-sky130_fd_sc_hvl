* File: sky130_fd_sc_hvl__nor3_1.pxi.spice
* Created: Fri Aug 28 09:38:18 2020
* 
x_PM_SKY130_FD_SC_HVL__NOR3_1%VNB N_VNB_M1003_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__NOR3_1%VNB
x_PM_SKY130_FD_SC_HVL__NOR3_1%VPB N_VPB_M1000_b VPB N_VPB_c_25_p N_VPB_c_26_p
+ VPB PM_SKY130_FD_SC_HVL__NOR3_1%VPB
x_PM_SKY130_FD_SC_HVL__NOR3_1%A N_A_M1003_g N_A_M1000_g A A N_A_c_48_n
+ PM_SKY130_FD_SC_HVL__NOR3_1%A
x_PM_SKY130_FD_SC_HVL__NOR3_1%B B B B N_B_M1005_g N_B_M1001_g
+ PM_SKY130_FD_SC_HVL__NOR3_1%B
x_PM_SKY130_FD_SC_HVL__NOR3_1%C N_C_M1002_g N_C_M1004_g C C C C N_C_c_102_n
+ N_C_c_110_n N_C_c_104_n PM_SKY130_FD_SC_HVL__NOR3_1%C
x_PM_SKY130_FD_SC_HVL__NOR3_1%VPWR N_VPWR_M1000_s VPWR N_VPWR_c_129_n VPWR
+ PM_SKY130_FD_SC_HVL__NOR3_1%VPWR
x_PM_SKY130_FD_SC_HVL__NOR3_1%Y N_Y_M1003_d N_Y_M1004_d N_Y_M1002_d N_Y_c_148_n
+ N_Y_c_150_n N_Y_c_151_n N_Y_c_152_n Y Y Y Y Y Y PM_SKY130_FD_SC_HVL__NOR3_1%Y
x_PM_SKY130_FD_SC_HVL__NOR3_1%VGND N_VGND_M1003_s N_VGND_M1005_d VGND
+ N_VGND_c_186_n N_VGND_c_188_n N_VGND_c_190_n VGND
+ PM_SKY130_FD_SC_HVL__NOR3_1%VGND
cc_1 N_VNB_M1003_b N_A_M1003_g 0.0497587f $X=-0.33 $Y=-0.265 $X2=0.705 $Y2=0.91
cc_2 N_VNB_c_2_p N_A_M1003_g 0.00128467f $X=3.12 $Y=0 $X2=0.705 $Y2=0.91
cc_3 N_VNB_M1003_b N_A_c_48_n 0.0883861f $X=-0.33 $Y=-0.265 $X2=0.775 $Y2=1.665
cc_4 N_VNB_M1003_b B 0.0032323f $X=-0.33 $Y=-0.265 $X2=0.705 $Y2=0.91
cc_5 N_VNB_M1003_b N_B_M1005_g 0.0797958f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_c_2_p N_B_M1005_g 5.86481e-19 $X=3.12 $Y=0 $X2=0 $Y2=0
cc_7 N_VNB_M1003_b N_C_M1004_g 0.0653582f $X=-0.33 $Y=-0.265 $X2=0.775 $Y2=2.965
cc_8 N_VNB_c_2_p N_C_M1004_g 9.58849e-19 $X=3.12 $Y=0 $X2=0.775 $Y2=2.965
cc_9 N_VNB_M1003_b N_C_c_102_n 0.0314103f $X=-0.33 $Y=-0.265 $X2=0.705 $Y2=1.665
cc_10 N_VNB_M1003_b N_Y_c_148_n 0.00995666f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_11 N_VNB_c_2_p N_Y_c_148_n 6.32535e-19 $X=3.12 $Y=0 $X2=0 $Y2=0
cc_12 N_VNB_M1003_b N_Y_c_150_n 0.0112009f $X=-0.33 $Y=-0.265 $X2=0.29 $Y2=1.69
cc_13 N_VNB_M1003_b N_Y_c_151_n 0.00148421f $X=-0.33 $Y=-0.265 $X2=0.29 $Y2=1.69
cc_14 N_VNB_M1003_b N_Y_c_152_n 0.0149107f $X=-0.33 $Y=-0.265 $X2=0.775
+ $Y2=1.665
cc_15 N_VNB_c_2_p N_Y_c_152_n 6.67688e-19 $X=3.12 $Y=0 $X2=0.775 $Y2=1.665
cc_16 N_VNB_M1003_b Y 0.00730093f $X=-0.33 $Y=-0.265 $X2=0.275 $Y2=1.665
cc_17 N_VNB_M1003_b Y 0.0111156f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_18 N_VNB_M1003_b N_VGND_c_186_n 0.0675832f $X=-0.33 $Y=-0.265 $X2=0.155
+ $Y2=1.95
cc_19 N_VNB_c_2_p N_VGND_c_186_n 0.00166879f $X=3.12 $Y=0 $X2=0.155 $Y2=1.95
cc_20 N_VNB_M1003_b N_VGND_c_188_n 0.0470117f $X=-0.33 $Y=-0.265 $X2=0.705
+ $Y2=1.665
cc_21 N_VNB_c_2_p N_VGND_c_188_n 0.00269049f $X=3.12 $Y=0 $X2=0.705 $Y2=1.665
cc_22 N_VNB_M1003_b N_VGND_c_190_n 0.093576f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_23 N_VNB_c_2_p N_VGND_c_190_n 0.35939f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_24 N_VPB_M1000_b N_A_M1000_g 0.0556136f $X=-0.33 $Y=1.885 $X2=0.775 $Y2=2.965
cc_25 N_VPB_c_25_p N_A_M1000_g 0.0137101f $X=3.12 $Y=4.07 $X2=0.775 $Y2=2.965
cc_26 N_VPB_c_26_p N_A_M1000_g 0.00970178f $X=3.12 $Y=4.07 $X2=0.775 $Y2=2.965
cc_27 N_VPB_M1000_b A 0.0118924f $X=-0.33 $Y=1.885 $X2=0.155 $Y2=1.58
cc_28 N_VPB_M1000_b N_A_c_48_n 0.0170594f $X=-0.33 $Y=1.885 $X2=0.775 $Y2=1.665
cc_29 N_VPB_M1000_b B 0.00501275f $X=-0.33 $Y=1.885 $X2=0.705 $Y2=0.91
cc_30 N_VPB_M1000_b N_B_M1005_g 0.0483363f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_31 N_VPB_c_25_p N_B_M1005_g 0.0137101f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_32 N_VPB_c_26_p N_B_M1005_g 0.00970178f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_33 N_VPB_M1000_b N_C_c_102_n 0.0265187f $X=-0.33 $Y=1.885 $X2=0.705 $Y2=1.665
cc_34 N_VPB_M1000_b N_C_c_104_n 0.0365691f $X=-0.33 $Y=1.885 $X2=0.275 $Y2=1.665
cc_35 N_VPB_c_25_p N_C_c_104_n 0.0196751f $X=3.12 $Y=4.07 $X2=0.275 $Y2=1.665
cc_36 N_VPB_c_26_p N_C_c_104_n 0.00970178f $X=3.12 $Y=4.07 $X2=0.275 $Y2=1.665
cc_37 N_VPB_M1000_b VPWR 0.0684523f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_38 N_VPB_c_25_p VPWR 0.0173213f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_39 N_VPB_c_26_p VPWR 0.356869f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_40 N_VPB_M1000_b N_VPWR_c_129_n 0.0639637f $X=-0.33 $Y=1.885 $X2=0.775
+ $Y2=2.965
cc_41 N_VPB_c_25_p N_VPWR_c_129_n 0.0841836f $X=3.12 $Y=4.07 $X2=0.775 $Y2=2.965
cc_42 N_VPB_c_26_p N_VPWR_c_129_n 0.00684647f $X=3.12 $Y=4.07 $X2=0.775
+ $Y2=2.965
cc_43 N_VPB_M1000_b Y 0.0653471f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_44 N_VPB_c_25_p Y 0.0138976f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_45 N_VPB_c_26_p Y 8.06088e-19 $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_46 N_A_M1000_g B 0.0174876f $X=0.775 $Y=2.965 $X2=0 $Y2=0
cc_47 A B 0.0267563f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_48 N_A_c_48_n B 0.0240431f $X=0.775 $Y=1.665 $X2=0 $Y2=0
cc_49 N_A_M1003_g N_B_M1005_g 0.0171339f $X=0.705 $Y=0.91 $X2=0 $Y2=0
cc_50 N_A_c_48_n N_B_M1005_g 0.164643f $X=0.775 $Y=1.665 $X2=0 $Y2=0
cc_51 N_A_M1000_g VPWR 0.00233065f $X=0.775 $Y=2.965 $X2=0 $Y2=0
cc_52 N_A_M1000_g N_VPWR_c_129_n 0.0959019f $X=0.775 $Y=2.965 $X2=0 $Y2=0
cc_53 A N_VPWR_c_129_n 0.0262091f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_54 N_A_c_48_n N_VPWR_c_129_n 0.00499082f $X=0.775 $Y=1.665 $X2=0 $Y2=0
cc_55 N_A_M1003_g N_Y_c_148_n 0.0219702f $X=0.705 $Y=0.91 $X2=0 $Y2=0
cc_56 N_A_c_48_n N_Y_c_148_n 0.00230731f $X=0.775 $Y=1.665 $X2=0 $Y2=0
cc_57 A N_Y_c_151_n 0.0022759f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_58 N_A_c_48_n N_Y_c_151_n 0.0115313f $X=0.775 $Y=1.665 $X2=0 $Y2=0
cc_59 N_A_M1003_g N_VGND_c_186_n 0.0523043f $X=0.705 $Y=0.91 $X2=0.24 $Y2=0
cc_60 A N_VGND_c_186_n 0.0232634f $X=0.155 $Y=1.58 $X2=0.24 $Y2=0
cc_61 N_A_c_48_n N_VGND_c_186_n 0.0111074f $X=0.775 $Y=1.665 $X2=0.24 $Y2=0
cc_62 N_A_M1003_g N_VGND_c_188_n 0.00110089f $X=0.705 $Y=0.91 $X2=3.12 $Y2=0
cc_63 N_A_M1003_g N_VGND_c_190_n 0.0153388f $X=0.705 $Y=0.91 $X2=0.24 $Y2=0
cc_64 N_B_M1005_g N_C_M1004_g 0.0278295f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_65 B N_C_c_102_n 0.00238952f $X=1.595 $Y=1.95 $X2=3.12 $Y2=0
cc_66 N_B_M1005_g N_C_c_102_n 0.151092f $X=1.485 $Y=0.91 $X2=3.12 $Y2=0
cc_67 B N_C_c_110_n 0.0276703f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_68 N_B_M1005_g N_C_c_110_n 0.00270278f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_69 N_B_M1005_g VPWR 0.00178648f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_70 B N_VPWR_c_129_n 0.0839418f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_71 N_B_M1005_g N_VPWR_c_129_n 0.0943249f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_72 N_B_M1005_g N_Y_c_148_n 0.00472529f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_73 B N_Y_c_150_n 0.0429816f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_74 N_B_M1005_g N_Y_c_150_n 0.0293191f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_75 B N_Y_c_151_n 0.0204336f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_76 B N_VGND_c_186_n 0.00268541f $X=1.595 $Y=1.95 $X2=0.24 $Y2=0
cc_77 N_B_M1005_g N_VGND_c_186_n 8.41089e-19 $X=1.485 $Y=0.91 $X2=0.24 $Y2=0
cc_78 N_B_M1005_g N_VGND_c_188_n 0.050898f $X=1.485 $Y=0.91 $X2=3.12 $Y2=0
cc_79 N_B_M1005_g N_VGND_c_190_n 0.00778503f $X=1.485 $Y=0.91 $X2=0.24 $Y2=0
cc_80 N_C_c_110_n VPWR 0.0158931f $X=2.14 $Y=1.89 $X2=0 $Y2=0
cc_81 N_C_c_104_n VPWR 0.0230278f $X=2.23 $Y=2.105 $X2=0 $Y2=0
cc_82 N_C_c_104_n N_VPWR_c_129_n 0.00724412f $X=2.23 $Y=2.105 $X2=0 $Y2=0
cc_83 N_C_M1004_g N_Y_c_150_n 0.0337297f $X=2.265 $Y=0.91 $X2=0 $Y2=0
cc_84 N_C_c_102_n N_Y_c_150_n 0.00278092f $X=2.14 $Y=1.89 $X2=0 $Y2=0
cc_85 N_C_c_110_n N_Y_c_150_n 0.0240062f $X=2.14 $Y=1.89 $X2=0 $Y2=0
cc_86 N_C_M1004_g N_Y_c_152_n 0.024718f $X=2.265 $Y=0.91 $X2=0 $Y2=0
cc_87 N_C_M1004_g Y 0.00365193f $X=2.265 $Y=0.91 $X2=0 $Y2=0
cc_88 N_C_M1004_g Y 5.02484e-19 $X=2.265 $Y=0.91 $X2=0 $Y2=0
cc_89 N_C_c_102_n Y 0.0236175f $X=2.14 $Y=1.89 $X2=0 $Y2=0
cc_90 N_C_c_110_n Y 0.0673558f $X=2.14 $Y=1.89 $X2=0 $Y2=0
cc_91 N_C_c_104_n Y 0.009101f $X=2.23 $Y=2.105 $X2=0 $Y2=0
cc_92 N_C_M1004_g N_VGND_c_188_n 0.0469268f $X=2.265 $Y=0.91 $X2=3.12 $Y2=0
cc_93 N_C_M1004_g N_VGND_c_190_n 0.0118525f $X=2.265 $Y=0.91 $X2=0.24 $Y2=0
cc_94 N_VPWR_c_129_n A_205_443# 0.00109099f $X=0.385 $Y=2.385 $X2=0 $Y2=3.985
cc_95 VPWR A_347_443# 0.00767357f $X=0 $Y=3.445 $X2=0 $Y2=3.985
cc_96 VPWR N_Y_M1002_d 0.00179328f $X=0 $Y=3.445 $X2=0 $Y2=0
cc_97 VPWR Y 0.046643f $X=0 $Y=3.445 $X2=0 $Y2=0
cc_98 N_Y_c_148_n N_VGND_c_186_n 0.0451007f $X=1.095 $Y=0.66 $X2=0.24 $Y2=0
cc_99 N_Y_c_148_n N_VGND_c_188_n 0.0316828f $X=1.095 $Y=0.66 $X2=3.12 $Y2=0
cc_100 N_Y_c_150_n N_VGND_c_188_n 0.0658158f $X=2.49 $Y=1.51 $X2=3.12 $Y2=0
cc_101 N_Y_c_152_n N_VGND_c_188_n 0.0542931f $X=2.655 $Y=0.68 $X2=3.12 $Y2=0
cc_102 N_Y_M1003_d N_VGND_c_190_n 0.00221032f $X=0.955 $Y=0.535 $X2=0.24 $Y2=0
cc_103 N_Y_M1004_d N_VGND_c_190_n 0.00108431f $X=2.515 $Y=0.535 $X2=0.24 $Y2=0
cc_104 N_Y_c_148_n N_VGND_c_190_n 0.0247302f $X=1.095 $Y=0.66 $X2=0.24 $Y2=0
cc_105 N_Y_c_152_n N_VGND_c_190_n 0.0282633f $X=2.655 $Y=0.68 $X2=0.24 $Y2=0
