# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
SITE unithvdbl
    SYMMETRY y  ;
    CLASS CORE  ;
    SIZE  0.480 BY 8.140 ;
END unithvdbl
MACRO sky130_fd_sc_hvl__buf_32
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  33.60000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  11.25000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.220000 1.580000 4.630000 1.815000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  10.08000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.950000 2.290000 32.640000 2.520000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 33.600000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 33.600000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 33.600000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 33.600000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 33.600000 0.085000 ;
      RECT  0.000000  3.985000 33.600000 4.155000 ;
      RECT  0.110000  0.425000  0.645000 1.410000 ;
      RECT  0.110000  2.175000  0.680000 3.755000 ;
      RECT  0.815000  0.755000  1.170000 1.195000 ;
      RECT  0.815000  1.195000  7.410000 1.410000 ;
      RECT  0.850000  1.985000  7.410000 2.265000 ;
      RECT  0.850000  2.265000  1.160000 3.755000 ;
      RECT  1.340000  0.415000  2.230000 1.025000 ;
      RECT  1.340000  2.445000  2.230000 3.675000 ;
      RECT  2.400000  0.730000  2.790000 1.195000 ;
      RECT  2.400000  2.265000  2.710000 3.755000 ;
      RECT  2.880000  2.445000  3.770000 3.675000 ;
      RECT  2.960000  0.425000  3.855000 1.025000 ;
      RECT  3.940000  2.265000  4.290000 3.755000 ;
      RECT  4.025000  0.730000  4.270000 1.195000 ;
      RECT  4.440000  0.425000  5.330000 1.025000 ;
      RECT  4.460000  2.445000  5.350000 3.675000 ;
      RECT  4.800000  1.410000  7.410000 1.985000 ;
      RECT  5.520000  0.730000  5.910000 1.195000 ;
      RECT  5.520000  2.265000  5.830000 3.755000 ;
      RECT  6.000000  2.445000  6.890000 3.675000 ;
      RECT  6.080000  0.425000  6.975000 1.025000 ;
      RECT  7.060000  2.265000  7.410000 3.755000 ;
      RECT  7.145000  0.730000  7.390000 1.195000 ;
      RECT  7.560000  0.425000  8.480000 1.025000 ;
      RECT  7.580000  1.025000  8.480000 1.395000 ;
      RECT  7.580000  2.235000  8.480000 3.675000 ;
      RECT  8.930000  0.790000  9.260000 3.755000 ;
      RECT  9.430000  0.425000 10.320000 1.395000 ;
      RECT  9.430000  2.175000 10.320000 3.755000 ;
      RECT  9.520000  1.565000 10.190000 1.895000 ;
      RECT 10.490000  0.790000 10.820000 3.755000 ;
      RECT 10.990000  0.425000 11.880000 1.395000 ;
      RECT 10.990000  2.175000 11.880000 3.755000 ;
      RECT 11.080000  1.565000 11.750000 1.895000 ;
      RECT 12.050000  0.790000 12.380000 3.755000 ;
      RECT 12.550000  0.425000 13.440000 1.395000 ;
      RECT 12.550000  2.175000 13.440000 3.755000 ;
      RECT 12.640000  1.565000 13.310000 1.895000 ;
      RECT 13.610000  0.790000 13.940000 3.755000 ;
      RECT 14.110000  0.425000 15.000000 1.395000 ;
      RECT 14.110000  2.175000 15.000000 3.755000 ;
      RECT 14.200000  1.565000 14.870000 1.895000 ;
      RECT 15.170000  0.790000 15.500000 3.755000 ;
      RECT 15.670000  0.425000 16.560000 1.395000 ;
      RECT 15.670000  2.175000 16.560000 3.755000 ;
      RECT 15.760000  1.565000 16.430000 1.895000 ;
      RECT 16.730000  0.790000 17.060000 3.755000 ;
      RECT 17.230000  0.425000 18.120000 1.395000 ;
      RECT 17.230000  2.175000 18.120000 3.755000 ;
      RECT 17.320000  1.565000 17.990000 1.895000 ;
      RECT 18.290000  0.790000 18.620000 3.755000 ;
      RECT 18.790000  0.425000 19.680000 1.395000 ;
      RECT 18.790000  2.175000 19.680000 3.755000 ;
      RECT 18.880000  1.565000 19.550000 1.895000 ;
      RECT 19.850000  0.790000 20.260000 3.755000 ;
      RECT 20.430000  0.425000 20.960000 1.395000 ;
      RECT 20.430000  1.565000 21.100000 1.895000 ;
      RECT 20.430000  2.175000 20.960000 3.755000 ;
      RECT 21.410000  0.790000 21.740000 3.755000 ;
      RECT 21.910000  0.425000 22.800000 1.395000 ;
      RECT 21.910000  2.175000 22.800000 3.755000 ;
      RECT 22.000000  1.565000 22.670000 1.895000 ;
      RECT 22.970000  0.790000 23.300000 3.755000 ;
      RECT 23.470000  0.425000 24.360000 1.395000 ;
      RECT 23.470000  2.175000 24.360000 3.755000 ;
      RECT 23.560000  1.565000 24.230000 1.895000 ;
      RECT 24.530000  0.790000 24.860000 3.755000 ;
      RECT 25.030000  0.425000 25.920000 1.395000 ;
      RECT 25.030000  2.175000 25.920000 3.755000 ;
      RECT 25.120000  1.565000 25.790000 1.895000 ;
      RECT 26.090000  0.790000 26.420000 3.755000 ;
      RECT 26.590000  0.425000 27.480000 1.395000 ;
      RECT 26.590000  2.175000 27.480000 3.755000 ;
      RECT 26.680000  1.565000 27.350000 1.895000 ;
      RECT 27.650000  0.790000 27.980000 3.755000 ;
      RECT 28.150000  0.425000 29.040000 1.395000 ;
      RECT 28.150000  2.175000 29.040000 3.755000 ;
      RECT 28.240000  1.565000 28.910000 1.895000 ;
      RECT 29.210000  0.790000 29.540000 3.755000 ;
      RECT 29.710000  0.425000 30.600000 1.395000 ;
      RECT 29.710000  2.175000 30.600000 3.755000 ;
      RECT 29.800000  1.565000 30.470000 1.895000 ;
      RECT 30.770000  0.790000 31.100000 3.755000 ;
      RECT 31.270000  0.425000 32.160000 1.395000 ;
      RECT 31.270000  2.175000 32.160000 3.755000 ;
      RECT 31.360000  1.565000 32.030000 1.895000 ;
      RECT 32.330000  0.790000 32.740000 3.755000 ;
      RECT 32.910000  0.425000 33.440000 1.495000 ;
      RECT 32.910000  2.175000 33.440000 3.755000 ;
    LAYER mcon ;
      RECT  0.115000  0.425000  0.285000 0.595000 ;
      RECT  0.150000  3.475000  0.320000 3.645000 ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.475000  0.425000  0.645000 0.595000 ;
      RECT  0.510000  3.475000  0.680000 3.645000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.340000  0.425000  1.510000 0.595000 ;
      RECT  1.340000  3.475000  1.510000 3.645000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  1.700000  0.425000  1.870000 0.595000 ;
      RECT  1.700000  3.475000  1.870000 3.645000 ;
      RECT  2.060000  0.425000  2.230000 0.595000 ;
      RECT  2.060000  3.475000  2.230000 3.645000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.880000  3.475000  3.050000 3.645000 ;
      RECT  2.960000  0.425000  3.130000 0.595000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.240000  3.475000  3.410000 3.645000 ;
      RECT  3.320000  0.425000  3.490000 0.595000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.600000  3.475000  3.770000 3.645000 ;
      RECT  3.680000  0.425000  3.850000 0.595000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.440000  0.425000  4.610000 0.595000 ;
      RECT  4.460000  3.475000  4.630000 3.645000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.800000  0.425000  4.970000 0.595000 ;
      RECT  4.820000  3.475000  4.990000 3.645000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.020000  1.580000  5.190000 1.750000 ;
      RECT  5.160000  0.425000  5.330000 0.595000 ;
      RECT  5.180000  3.475000  5.350000 3.645000 ;
      RECT  5.380000  1.580000  5.550000 1.750000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.740000  1.580000  5.910000 1.750000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.000000  3.475000  6.170000 3.645000 ;
      RECT  6.080000  0.425000  6.250000 0.595000 ;
      RECT  6.100000  1.580000  6.270000 1.750000 ;
      RECT  6.360000  3.475000  6.530000 3.645000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.440000  0.425000  6.610000 0.595000 ;
      RECT  6.460000  1.580000  6.630000 1.750000 ;
      RECT  6.720000  3.475000  6.890000 3.645000 ;
      RECT  6.800000  0.425000  6.970000 0.595000 ;
      RECT  6.820000  1.580000  6.990000 1.750000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.180000  1.580000  7.350000 1.750000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.560000  0.425000  7.730000 0.595000 ;
      RECT  7.580000  3.475000  7.750000 3.645000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  7.920000  0.425000  8.090000 0.595000 ;
      RECT  7.940000  3.475000  8.110000 3.645000 ;
      RECT  8.280000  0.425000  8.450000 0.595000 ;
      RECT  8.300000  3.475000  8.470000 3.645000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.010000  2.320000  9.180000 2.490000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.430000  0.425000  9.600000 0.595000 ;
      RECT  9.430000  3.475000  9.600000 3.645000 ;
      RECT  9.590000  1.580000  9.760000 1.750000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.790000  0.425000  9.960000 0.595000 ;
      RECT  9.790000  3.475000  9.960000 3.645000 ;
      RECT  9.950000  1.580000 10.120000 1.750000 ;
      RECT 10.150000  0.425000 10.320000 0.595000 ;
      RECT 10.150000  3.475000 10.320000 3.645000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.570000  2.320000 10.740000 2.490000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.990000  0.425000 11.160000 0.595000 ;
      RECT 10.990000  3.475000 11.160000 3.645000 ;
      RECT 11.150000  1.580000 11.320000 1.750000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.350000  0.425000 11.520000 0.595000 ;
      RECT 11.350000  3.475000 11.520000 3.645000 ;
      RECT 11.510000  1.580000 11.680000 1.750000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 11.710000  0.425000 11.880000 0.595000 ;
      RECT 11.710000  3.475000 11.880000 3.645000 ;
      RECT 12.130000  2.320000 12.300000 2.490000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.550000  0.425000 12.720000 0.595000 ;
      RECT 12.550000  3.475000 12.720000 3.645000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 12.710000  1.580000 12.880000 1.750000 ;
      RECT 12.910000  0.425000 13.080000 0.595000 ;
      RECT 12.910000  3.475000 13.080000 3.645000 ;
      RECT 13.070000  1.580000 13.240000 1.750000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.270000  0.425000 13.440000 0.595000 ;
      RECT 13.270000  3.475000 13.440000 3.645000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.690000  2.320000 13.860000 2.490000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.110000  0.425000 14.280000 0.595000 ;
      RECT 14.110000  3.475000 14.280000 3.645000 ;
      RECT 14.270000  1.580000 14.440000 1.750000 ;
      RECT 14.470000  0.425000 14.640000 0.595000 ;
      RECT 14.470000  3.475000 14.640000 3.645000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.630000  1.580000 14.800000 1.750000 ;
      RECT 14.830000  0.425000 15.000000 0.595000 ;
      RECT 14.830000  3.475000 15.000000 3.645000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.250000  2.320000 15.420000 2.490000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.670000  0.425000 15.840000 0.595000 ;
      RECT 15.670000  3.475000 15.840000 3.645000 ;
      RECT 15.830000  1.580000 16.000000 1.750000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.030000  0.425000 16.200000 0.595000 ;
      RECT 16.030000  3.475000 16.200000 3.645000 ;
      RECT 16.190000  1.580000 16.360000 1.750000 ;
      RECT 16.390000  0.425000 16.560000 0.595000 ;
      RECT 16.390000  3.475000 16.560000 3.645000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.810000  2.320000 16.980000 2.490000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 17.230000  0.425000 17.400000 0.595000 ;
      RECT 17.230000  3.475000 17.400000 3.645000 ;
      RECT 17.390000  1.580000 17.560000 1.750000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
      RECT 17.590000  0.425000 17.760000 0.595000 ;
      RECT 17.590000  3.475000 17.760000 3.645000 ;
      RECT 17.750000  1.580000 17.920000 1.750000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.985000 18.085000 4.155000 ;
      RECT 17.950000  0.425000 18.120000 0.595000 ;
      RECT 17.950000  3.475000 18.120000 3.645000 ;
      RECT 18.370000  2.320000 18.540000 2.490000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.985000 18.565000 4.155000 ;
      RECT 18.790000  0.425000 18.960000 0.595000 ;
      RECT 18.790000  3.475000 18.960000 3.645000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  3.985000 19.045000 4.155000 ;
      RECT 18.950000  1.580000 19.120000 1.750000 ;
      RECT 19.150000  0.425000 19.320000 0.595000 ;
      RECT 19.150000  3.475000 19.320000 3.645000 ;
      RECT 19.310000  1.580000 19.480000 1.750000 ;
      RECT 19.355000 -0.085000 19.525000 0.085000 ;
      RECT 19.355000  3.985000 19.525000 4.155000 ;
      RECT 19.510000  0.425000 19.680000 0.595000 ;
      RECT 19.510000  3.475000 19.680000 3.645000 ;
      RECT 19.835000 -0.085000 20.005000 0.085000 ;
      RECT 19.835000  3.985000 20.005000 4.155000 ;
      RECT 19.930000  2.320000 20.100000 2.490000 ;
      RECT 20.315000 -0.085000 20.485000 0.085000 ;
      RECT 20.315000  3.985000 20.485000 4.155000 ;
      RECT 20.430000  0.425000 20.600000 0.595000 ;
      RECT 20.430000  3.475000 20.600000 3.645000 ;
      RECT 20.500000  1.580000 20.670000 1.750000 ;
      RECT 20.790000  0.425000 20.960000 0.595000 ;
      RECT 20.790000  3.475000 20.960000 3.645000 ;
      RECT 20.795000 -0.085000 20.965000 0.085000 ;
      RECT 20.795000  3.985000 20.965000 4.155000 ;
      RECT 20.860000  1.580000 21.030000 1.750000 ;
      RECT 21.275000 -0.085000 21.445000 0.085000 ;
      RECT 21.275000  3.985000 21.445000 4.155000 ;
      RECT 21.490000  2.320000 21.660000 2.490000 ;
      RECT 21.755000 -0.085000 21.925000 0.085000 ;
      RECT 21.755000  3.985000 21.925000 4.155000 ;
      RECT 21.910000  0.425000 22.080000 0.595000 ;
      RECT 21.910000  3.475000 22.080000 3.645000 ;
      RECT 22.070000  1.580000 22.240000 1.750000 ;
      RECT 22.235000 -0.085000 22.405000 0.085000 ;
      RECT 22.235000  3.985000 22.405000 4.155000 ;
      RECT 22.270000  0.425000 22.440000 0.595000 ;
      RECT 22.270000  3.475000 22.440000 3.645000 ;
      RECT 22.430000  1.580000 22.600000 1.750000 ;
      RECT 22.630000  0.425000 22.800000 0.595000 ;
      RECT 22.630000  3.475000 22.800000 3.645000 ;
      RECT 22.715000 -0.085000 22.885000 0.085000 ;
      RECT 22.715000  3.985000 22.885000 4.155000 ;
      RECT 23.050000  2.320000 23.220000 2.490000 ;
      RECT 23.195000 -0.085000 23.365000 0.085000 ;
      RECT 23.195000  3.985000 23.365000 4.155000 ;
      RECT 23.470000  0.425000 23.640000 0.595000 ;
      RECT 23.470000  3.475000 23.640000 3.645000 ;
      RECT 23.630000  1.580000 23.800000 1.750000 ;
      RECT 23.675000 -0.085000 23.845000 0.085000 ;
      RECT 23.675000  3.985000 23.845000 4.155000 ;
      RECT 23.830000  0.425000 24.000000 0.595000 ;
      RECT 23.830000  3.475000 24.000000 3.645000 ;
      RECT 23.990000  1.580000 24.160000 1.750000 ;
      RECT 24.155000 -0.085000 24.325000 0.085000 ;
      RECT 24.155000  3.985000 24.325000 4.155000 ;
      RECT 24.190000  0.425000 24.360000 0.595000 ;
      RECT 24.190000  3.475000 24.360000 3.645000 ;
      RECT 24.610000  2.320000 24.780000 2.490000 ;
      RECT 24.635000 -0.085000 24.805000 0.085000 ;
      RECT 24.635000  3.985000 24.805000 4.155000 ;
      RECT 25.030000  0.425000 25.200000 0.595000 ;
      RECT 25.030000  3.475000 25.200000 3.645000 ;
      RECT 25.115000 -0.085000 25.285000 0.085000 ;
      RECT 25.115000  3.985000 25.285000 4.155000 ;
      RECT 25.190000  1.580000 25.360000 1.750000 ;
      RECT 25.390000  0.425000 25.560000 0.595000 ;
      RECT 25.390000  3.475000 25.560000 3.645000 ;
      RECT 25.550000  1.580000 25.720000 1.750000 ;
      RECT 25.595000 -0.085000 25.765000 0.085000 ;
      RECT 25.595000  3.985000 25.765000 4.155000 ;
      RECT 25.750000  0.425000 25.920000 0.595000 ;
      RECT 25.750000  3.475000 25.920000 3.645000 ;
      RECT 26.075000 -0.085000 26.245000 0.085000 ;
      RECT 26.075000  3.985000 26.245000 4.155000 ;
      RECT 26.170000  2.320000 26.340000 2.490000 ;
      RECT 26.555000 -0.085000 26.725000 0.085000 ;
      RECT 26.555000  3.985000 26.725000 4.155000 ;
      RECT 26.590000  0.425000 26.760000 0.595000 ;
      RECT 26.590000  3.475000 26.760000 3.645000 ;
      RECT 26.750000  1.580000 26.920000 1.750000 ;
      RECT 26.950000  0.425000 27.120000 0.595000 ;
      RECT 26.950000  3.475000 27.120000 3.645000 ;
      RECT 27.035000 -0.085000 27.205000 0.085000 ;
      RECT 27.035000  3.985000 27.205000 4.155000 ;
      RECT 27.110000  1.580000 27.280000 1.750000 ;
      RECT 27.310000  0.425000 27.480000 0.595000 ;
      RECT 27.310000  3.475000 27.480000 3.645000 ;
      RECT 27.515000 -0.085000 27.685000 0.085000 ;
      RECT 27.515000  3.985000 27.685000 4.155000 ;
      RECT 27.730000  2.320000 27.900000 2.490000 ;
      RECT 27.995000 -0.085000 28.165000 0.085000 ;
      RECT 27.995000  3.985000 28.165000 4.155000 ;
      RECT 28.150000  0.425000 28.320000 0.595000 ;
      RECT 28.150000  3.475000 28.320000 3.645000 ;
      RECT 28.310000  1.580000 28.480000 1.750000 ;
      RECT 28.475000 -0.085000 28.645000 0.085000 ;
      RECT 28.475000  3.985000 28.645000 4.155000 ;
      RECT 28.510000  0.425000 28.680000 0.595000 ;
      RECT 28.510000  3.475000 28.680000 3.645000 ;
      RECT 28.670000  1.580000 28.840000 1.750000 ;
      RECT 28.870000  0.425000 29.040000 0.595000 ;
      RECT 28.870000  3.475000 29.040000 3.645000 ;
      RECT 28.955000 -0.085000 29.125000 0.085000 ;
      RECT 28.955000  3.985000 29.125000 4.155000 ;
      RECT 29.290000  2.320000 29.460000 2.490000 ;
      RECT 29.435000 -0.085000 29.605000 0.085000 ;
      RECT 29.435000  3.985000 29.605000 4.155000 ;
      RECT 29.710000  0.425000 29.880000 0.595000 ;
      RECT 29.710000  3.475000 29.880000 3.645000 ;
      RECT 29.870000  1.580000 30.040000 1.750000 ;
      RECT 29.915000 -0.085000 30.085000 0.085000 ;
      RECT 29.915000  3.985000 30.085000 4.155000 ;
      RECT 30.070000  0.425000 30.240000 0.595000 ;
      RECT 30.070000  3.475000 30.240000 3.645000 ;
      RECT 30.230000  1.580000 30.400000 1.750000 ;
      RECT 30.395000 -0.085000 30.565000 0.085000 ;
      RECT 30.395000  3.985000 30.565000 4.155000 ;
      RECT 30.430000  0.425000 30.600000 0.595000 ;
      RECT 30.430000  3.475000 30.600000 3.645000 ;
      RECT 30.850000  2.320000 31.020000 2.490000 ;
      RECT 30.875000 -0.085000 31.045000 0.085000 ;
      RECT 30.875000  3.985000 31.045000 4.155000 ;
      RECT 31.270000  0.425000 31.440000 0.595000 ;
      RECT 31.270000  3.475000 31.440000 3.645000 ;
      RECT 31.355000 -0.085000 31.525000 0.085000 ;
      RECT 31.355000  3.985000 31.525000 4.155000 ;
      RECT 31.430000  1.580000 31.600000 1.750000 ;
      RECT 31.630000  0.425000 31.800000 0.595000 ;
      RECT 31.630000  3.475000 31.800000 3.645000 ;
      RECT 31.790000  1.580000 31.960000 1.750000 ;
      RECT 31.835000 -0.085000 32.005000 0.085000 ;
      RECT 31.835000  3.985000 32.005000 4.155000 ;
      RECT 31.990000  0.425000 32.160000 0.595000 ;
      RECT 31.990000  3.475000 32.160000 3.645000 ;
      RECT 32.315000 -0.085000 32.485000 0.085000 ;
      RECT 32.315000  3.985000 32.485000 4.155000 ;
      RECT 32.410000  2.320000 32.580000 2.490000 ;
      RECT 32.795000 -0.085000 32.965000 0.085000 ;
      RECT 32.795000  3.985000 32.965000 4.155000 ;
      RECT 32.910000  0.425000 33.080000 0.595000 ;
      RECT 32.910000  3.475000 33.080000 3.645000 ;
      RECT 33.270000  0.425000 33.440000 0.595000 ;
      RECT 33.270000  3.475000 33.440000 3.645000 ;
      RECT 33.275000 -0.085000 33.445000 0.085000 ;
      RECT 33.275000  3.985000 33.445000 4.155000 ;
    LAYER met1 ;
      RECT 4.960000 1.550000 32.090000 1.780000 ;
  END
END sky130_fd_sc_hvl__buf_32
END LIBRARY
