* File: sky130_fd_sc_hvl__einvn_1.pxi.spice
* Created: Fri Aug 28 09:35:25 2020
* 
x_PM_SKY130_FD_SC_HVL__EINVN_1%VNB N_VNB_M1001_b VNB N_VNB_c_12_p VNB
+ PM_SKY130_FD_SC_HVL__EINVN_1%VNB
x_PM_SKY130_FD_SC_HVL__EINVN_1%VPB N_VPB_M1005_b VPB N_VPB_c_24_p VPB
+ PM_SKY130_FD_SC_HVL__EINVN_1%VPB
x_PM_SKY130_FD_SC_HVL__EINVN_1%TE_B N_TE_B_M1001_g N_TE_B_M1005_g N_TE_B_c_47_n
+ N_TE_B_c_48_n N_TE_B_M1004_g TE_B TE_B TE_B N_TE_B_c_45_n N_TE_B_c_56_p
+ PM_SKY130_FD_SC_HVL__EINVN_1%TE_B
x_PM_SKY130_FD_SC_HVL__EINVN_1%A_30_173# N_A_30_173#_M1001_s N_A_30_173#_M1005_s
+ N_A_30_173#_c_88_n N_A_30_173#_M1002_g N_A_30_173#_c_89_n N_A_30_173#_c_90_n
+ N_A_30_173#_c_91_n N_A_30_173#_c_92_n N_A_30_173#_c_93_n N_A_30_173#_c_95_n
+ PM_SKY130_FD_SC_HVL__EINVN_1%A_30_173#
x_PM_SKY130_FD_SC_HVL__EINVN_1%A N_A_M1000_g A A A A N_A_M1003_g N_A_c_133_n A A
+ PM_SKY130_FD_SC_HVL__EINVN_1%A
x_PM_SKY130_FD_SC_HVL__EINVN_1%VPWR N_VPWR_M1005_d VPWR N_VPWR_c_166_n
+ N_VPWR_c_169_n PM_SKY130_FD_SC_HVL__EINVN_1%VPWR
x_PM_SKY130_FD_SC_HVL__EINVN_1%Z N_Z_M1003_d N_Z_M1000_d Z Z Z Z Z Z Z
+ N_Z_c_193_n PM_SKY130_FD_SC_HVL__EINVN_1%Z
x_PM_SKY130_FD_SC_HVL__EINVN_1%VGND N_VGND_M1001_d VGND N_VGND_c_206_n
+ N_VGND_c_208_n PM_SKY130_FD_SC_HVL__EINVN_1%VGND
cc_1 N_VNB_M1001_b N_TE_B_M1001_g 0.0698509f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=1.075
cc_2 N_VNB_M1001_b TE_B 0.00501792f $X=-0.33 $Y=-0.265 $X2=1.595 $Y2=1.95
cc_3 N_VNB_M1001_b N_TE_B_c_45_n 0.0466027f $X=-0.33 $Y=-0.265 $X2=1.185
+ $Y2=1.855
cc_4 N_VNB_M1001_b N_A_30_173#_c_88_n 0.0420434f $X=-0.33 $Y=-0.265 $X2=0.76
+ $Y2=2.61
cc_5 N_VNB_M1001_b N_A_30_173#_c_89_n 0.0217245f $X=-0.33 $Y=-0.265 $X2=1.815
+ $Y2=2.965
cc_6 N_VNB_M1001_b N_A_30_173#_c_90_n 0.0121912f $X=-0.33 $Y=-0.265 $X2=1.115
+ $Y2=1.95
cc_7 N_VNB_M1001_b N_A_30_173#_c_91_n 0.00710377f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=1.855
cc_8 N_VNB_M1001_b N_A_30_173#_c_92_n 0.0622851f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_M1001_b N_A_30_173#_c_93_n 0.0110756f $X=-0.33 $Y=-0.265 $X2=1.02
+ $Y2=1.855
cc_10 N_VNB_M1001_b A 0.00330514f $X=-0.33 $Y=-0.265 $X2=0.76 $Y2=2.61
cc_11 N_VNB_M1001_b N_A_M1003_g 0.0745362f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_12 N_VNB_c_12_p N_A_M1003_g 5.81826e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_13 N_VNB_M1001_b N_A_c_133_n 0.0250732f $X=-0.33 $Y=-0.265 $X2=1.02 $Y2=1.855
cc_14 N_VNB_M1001_b N_Z_c_193_n 0.0693798f $X=-0.33 $Y=-0.265 $X2=0.76 $Y2=1.855
cc_15 N_VNB_c_12_p N_Z_c_193_n 6.63219e-19 $X=0.24 $Y=0 $X2=0.76 $Y2=1.855
cc_16 N_VNB_M1001_b N_VGND_c_206_n 0.0746313f $X=-0.33 $Y=-0.265 $X2=1.185
+ $Y2=2.022
cc_17 N_VNB_c_12_p N_VGND_c_206_n 0.359247f $X=0.24 $Y=0 $X2=1.185 $Y2=2.022
cc_18 N_VNB_M1001_b N_VGND_c_208_n 0.12837f $X=-0.33 $Y=-0.265 $X2=1.815
+ $Y2=2.965
cc_19 N_VNB_c_12_p N_VGND_c_208_n 0.00662201f $X=0.24 $Y=0 $X2=1.815 $Y2=2.965
cc_20 N_VPB_M1005_b N_TE_B_M1005_g 0.0459093f $X=-0.33 $Y=1.885 $X2=0.76
+ $Y2=2.61
cc_21 N_VPB_M1005_b N_TE_B_c_47_n 0.0413175f $X=-0.33 $Y=1.885 $X2=1.565
+ $Y2=2.022
cc_22 N_VPB_M1005_b N_TE_B_c_48_n 0.0376535f $X=-0.33 $Y=1.885 $X2=1.815
+ $Y2=2.105
cc_23 VPB N_TE_B_c_48_n 0.00970178f $X=0 $Y=3.955 $X2=1.815 $Y2=2.105
cc_24 N_VPB_c_24_p N_TE_B_c_48_n 0.0137101f $X=3.12 $Y=4.07 $X2=1.815 $Y2=2.105
cc_25 N_VPB_M1005_b TE_B 0.00582731f $X=-0.33 $Y=1.885 $X2=1.595 $Y2=1.95
cc_26 N_VPB_M1005_b N_TE_B_c_45_n 0.0299585f $X=-0.33 $Y=1.885 $X2=1.185
+ $Y2=1.855
cc_27 N_VPB_M1005_b N_A_30_173#_c_90_n 0.0161622f $X=-0.33 $Y=1.885 $X2=1.115
+ $Y2=1.95
cc_28 N_VPB_M1005_b N_A_30_173#_c_95_n 0.0452329f $X=-0.33 $Y=1.885 $X2=1.02
+ $Y2=1.91
cc_29 N_VPB_M1005_b N_A_M1000_g 0.0415498f $X=-0.33 $Y=1.885 $X2=0.665 $Y2=1.075
cc_30 VPB N_A_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.665 $Y2=1.075
cc_31 N_VPB_c_24_p N_A_M1000_g 0.0152014f $X=3.12 $Y=4.07 $X2=0.665 $Y2=1.075
cc_32 N_VPB_M1005_b N_A_c_133_n 0.0224936f $X=-0.33 $Y=1.885 $X2=1.02 $Y2=1.855
cc_33 N_VPB_M1005_b A 0.00166534f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_34 N_VPB_M1005_b N_VPWR_c_166_n 0.031636f $X=-0.33 $Y=1.885 $X2=1.815
+ $Y2=2.105
cc_35 VPB N_VPWR_c_166_n 0.00773923f $X=0 $Y=3.955 $X2=1.815 $Y2=2.105
cc_36 N_VPB_c_24_p N_VPWR_c_166_n 0.103807f $X=3.12 $Y=4.07 $X2=1.815 $Y2=2.105
cc_37 N_VPB_M1005_b N_VPWR_c_169_n 0.0608255f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.95
cc_38 VPB N_VPWR_c_169_n 0.357529f $X=0 $Y=3.955 $X2=0.635 $Y2=1.95
cc_39 N_VPB_c_24_p N_VPWR_c_169_n 0.0159797f $X=3.12 $Y=4.07 $X2=0.635 $Y2=1.95
cc_40 N_VPB_M1005_b N_Z_c_193_n 0.0711858f $X=-0.33 $Y=1.885 $X2=0.76 $Y2=1.855
cc_41 VPB N_Z_c_193_n 8.67388e-19 $X=0 $Y=3.955 $X2=0.76 $Y2=1.855
cc_42 N_VPB_c_24_p N_Z_c_193_n 0.0149544f $X=3.12 $Y=4.07 $X2=0.76 $Y2=1.855
cc_43 N_TE_B_M1001_g N_A_30_173#_c_89_n 0.0174876f $X=0.665 $Y=1.075 $X2=0 $Y2=0
cc_44 N_TE_B_M1005_g N_A_30_173#_c_90_n 0.00346525f $X=0.76 $Y=2.61 $X2=0 $Y2=0
cc_45 N_TE_B_c_45_n N_A_30_173#_c_90_n 0.0171643f $X=1.185 $Y=1.855 $X2=0 $Y2=0
cc_46 N_TE_B_c_56_p N_A_30_173#_c_90_n 0.0216659f $X=0.93 $Y=1.972 $X2=0 $Y2=0
cc_47 N_TE_B_M1001_g N_A_30_173#_c_91_n 0.0230969f $X=0.665 $Y=1.075 $X2=0 $Y2=0
cc_48 N_TE_B_c_47_n N_A_30_173#_c_91_n 0.00261282f $X=1.565 $Y=2.022 $X2=0 $Y2=0
cc_49 TE_B N_A_30_173#_c_91_n 0.0628791f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_50 N_TE_B_c_45_n N_A_30_173#_c_91_n 0.0193301f $X=1.185 $Y=1.855 $X2=0 $Y2=0
cc_51 N_TE_B_c_56_p N_A_30_173#_c_91_n 0.0284976f $X=0.93 $Y=1.972 $X2=0 $Y2=0
cc_52 N_TE_B_M1001_g N_A_30_173#_c_92_n 0.00492567f $X=0.665 $Y=1.075 $X2=1.68
+ $Y2=0
cc_53 N_TE_B_c_47_n N_A_30_173#_c_92_n 0.0451892f $X=1.565 $Y=2.022 $X2=1.68
+ $Y2=0
cc_54 TE_B N_A_30_173#_c_92_n 0.00273599f $X=1.595 $Y=1.95 $X2=1.68 $Y2=0
cc_55 N_TE_B_c_45_n N_A_30_173#_c_92_n 0.00970155f $X=1.185 $Y=1.855 $X2=1.68
+ $Y2=0
cc_56 N_TE_B_M1001_g N_A_30_173#_c_93_n 0.00409122f $X=0.665 $Y=1.075 $X2=1.68
+ $Y2=0.057
cc_57 N_TE_B_c_45_n N_A_30_173#_c_93_n 0.00149451f $X=1.185 $Y=1.855 $X2=1.68
+ $Y2=0.057
cc_58 N_TE_B_M1005_g N_A_30_173#_c_95_n 0.0189913f $X=0.76 $Y=2.61 $X2=1.68
+ $Y2=0.058
cc_59 N_TE_B_c_45_n N_A_30_173#_c_95_n 0.00145162f $X=1.185 $Y=1.855 $X2=1.68
+ $Y2=0.058
cc_60 N_TE_B_c_56_p N_A_30_173#_c_95_n 0.001051f $X=0.93 $Y=1.972 $X2=1.68
+ $Y2=0.058
cc_61 N_TE_B_c_47_n N_A_M1000_g 0.0664946f $X=1.565 $Y=2.022 $X2=0 $Y2=0
cc_62 N_TE_B_c_47_n A 5.38795e-19 $X=1.565 $Y=2.022 $X2=0 $Y2=0
cc_63 TE_B A 0.0111101f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_64 N_TE_B_c_47_n N_A_c_133_n 0.00817559f $X=1.565 $Y=2.022 $X2=1.68 $Y2=0.057
cc_65 TE_B N_A_c_133_n 0.00272508f $X=1.595 $Y=1.95 $X2=1.68 $Y2=0.057
cc_66 N_TE_B_c_47_n A 0.00544628f $X=1.565 $Y=2.022 $X2=0 $Y2=0
cc_67 N_TE_B_c_48_n A 8.46551e-19 $X=1.815 $Y=2.105 $X2=0 $Y2=0
cc_68 N_TE_B_M1005_g N_VPWR_c_166_n 0.0623823f $X=0.76 $Y=2.61 $X2=0.24 $Y2=0
cc_69 N_TE_B_c_48_n N_VPWR_c_166_n 0.0979109f $X=1.815 $Y=2.105 $X2=0.24 $Y2=0
cc_70 TE_B N_VPWR_c_166_n 0.0642361f $X=1.595 $Y=1.95 $X2=0.24 $Y2=0
cc_71 N_TE_B_c_45_n N_VPWR_c_166_n 0.00284873f $X=1.185 $Y=1.855 $X2=0.24 $Y2=0
cc_72 N_TE_B_c_56_p N_VPWR_c_166_n 0.0144384f $X=0.93 $Y=1.972 $X2=0.24 $Y2=0
cc_73 N_TE_B_M1005_g N_VPWR_c_169_n 0.00659903f $X=0.76 $Y=2.61 $X2=0 $Y2=0
cc_74 N_TE_B_c_48_n N_VPWR_c_169_n 0.00262016f $X=1.815 $Y=2.105 $X2=0 $Y2=0
cc_75 N_TE_B_M1001_g N_VGND_c_206_n 8.16601e-19 $X=0.665 $Y=1.075 $X2=0.24 $Y2=0
cc_76 N_TE_B_M1001_g N_VGND_c_208_n 0.0560884f $X=0.665 $Y=1.075 $X2=0 $Y2=0
cc_77 N_TE_B_c_45_n N_VGND_c_208_n 0.00126795f $X=1.185 $Y=1.855 $X2=0 $Y2=0
cc_78 N_A_30_173#_c_88_n A 0.00144272f $X=1.935 $Y=1.395 $X2=-0.33 $Y2=-0.265
cc_79 N_A_30_173#_c_91_n A 0.00793179f $X=1.9 $Y=1.56 $X2=-0.33 $Y2=-0.265
cc_80 N_A_30_173#_c_92_n A 6.11791e-19 $X=1.9 $Y=1.56 $X2=-0.33 $Y2=-0.265
cc_81 N_A_30_173#_c_88_n N_A_M1003_g 0.0737549f $X=1.935 $Y=1.395 $X2=3.12 $Y2=0
cc_82 N_A_30_173#_c_91_n N_A_M1003_g 8.85892e-19 $X=1.9 $Y=1.56 $X2=3.12 $Y2=0
cc_83 N_A_30_173#_c_92_n N_A_M1003_g 0.00856358f $X=1.9 $Y=1.56 $X2=3.12 $Y2=0
cc_84 N_A_30_173#_c_92_n N_A_c_133_n 3.73923e-19 $X=1.9 $Y=1.56 $X2=1.68
+ $Y2=0.057
cc_85 N_A_30_173#_c_91_n N_VPWR_c_166_n 0.0067663f $X=1.9 $Y=1.56 $X2=0.24 $Y2=0
cc_86 N_A_30_173#_c_92_n N_VPWR_c_166_n 6.93292e-19 $X=1.9 $Y=1.56 $X2=0.24
+ $Y2=0
cc_87 N_A_30_173#_c_95_n N_VPWR_c_166_n 0.0509129f $X=0.37 $Y=2.36 $X2=0.24
+ $Y2=0
cc_88 N_A_30_173#_c_95_n N_VPWR_c_169_n 0.0198345f $X=0.37 $Y=2.36 $X2=0 $Y2=0
cc_89 N_A_30_173#_c_89_n N_VGND_c_206_n 0.0176561f $X=0.275 $Y=1.075 $X2=0.24
+ $Y2=0
cc_90 N_A_30_173#_c_88_n N_VGND_c_208_n 0.0704198f $X=1.935 $Y=1.395 $X2=0 $Y2=0
cc_91 N_A_30_173#_c_89_n N_VGND_c_208_n 0.0268555f $X=0.275 $Y=1.075 $X2=0 $Y2=0
cc_92 N_A_30_173#_c_91_n N_VGND_c_208_n 0.106793f $X=1.9 $Y=1.56 $X2=0 $Y2=0
cc_93 N_A_30_173#_c_92_n N_VGND_c_208_n 0.00680039f $X=1.9 $Y=1.56 $X2=0 $Y2=0
cc_94 N_A_M1000_g N_VPWR_c_166_n 0.0660853f $X=2.645 $Y=2.965 $X2=0.24 $Y2=0
cc_95 N_A_c_133_n N_VPWR_c_166_n 2.89617e-19 $X=2.44 $Y=1.89 $X2=0.24 $Y2=0
cc_96 A N_VPWR_c_166_n 0.0373341f $X=2.64 $Y=2.035 $X2=0.24 $Y2=0
cc_97 N_A_M1000_g N_VPWR_c_169_n 0.00857457f $X=2.645 $Y=2.965 $X2=0 $Y2=0
cc_98 A A_413_443# 0.00394495f $X=2.64 $Y=2.035 $X2=0 $Y2=0
cc_99 A N_Z_c_193_n 0.0908993f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_100 N_A_M1003_g N_Z_c_193_n 0.033719f $X=2.645 $Y=0.91 $X2=0 $Y2=0
cc_101 A N_VGND_c_206_n 0.00147299f $X=2.555 $Y=1.21 $X2=0.24 $Y2=0
cc_102 N_A_M1003_g N_VGND_c_206_n 0.00841297f $X=2.645 $Y=0.91 $X2=0.24 $Y2=0
cc_103 A N_VGND_c_208_n 0.0212421f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_104 A N_VGND_c_208_n 0.00229459f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_105 N_A_M1003_g N_VGND_c_208_n 0.0474117f $X=2.645 $Y=0.91 $X2=0 $Y2=0
cc_106 N_A_c_133_n N_VGND_c_208_n 3.98931e-19 $X=2.44 $Y=1.89 $X2=0 $Y2=0
cc_107 N_VPWR_c_166_n A_413_443# 0.00758262f $X=0.855 $Y=3.59 $X2=0 $Y2=3.985
cc_108 N_VPWR_c_169_n N_Z_M1000_d 0.00221032f $X=2.655 $Y=3.59 $X2=0 $Y2=0
cc_109 N_VPWR_c_166_n N_Z_c_193_n 0.0451154f $X=0.855 $Y=3.59 $X2=1.68 $Y2=4.07
cc_110 N_VPWR_c_169_n N_Z_c_193_n 0.0387829f $X=2.655 $Y=3.59 $X2=1.68 $Y2=4.07
cc_111 N_Z_M1003_d N_VGND_c_206_n 0.00221032f $X=2.895 $Y=0.535 $X2=0.24 $Y2=0
cc_112 N_Z_c_193_n N_VGND_c_206_n 0.0294061f $X=3.035 $Y=0.66 $X2=0.24 $Y2=0
cc_113 N_Z_c_193_n N_VGND_c_208_n 0.0179684f $X=3.035 $Y=0.66 $X2=0 $Y2=0
cc_114 N_VGND_c_208_n A_437_107# 0.00694399f $X=1.545 $Y=0.66 $X2=0 $Y2=0
