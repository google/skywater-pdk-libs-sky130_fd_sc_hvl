* File: sky130_fd_sc_hvl__probe_p_8.pex.spice
* Created: Wed Sep  2 09:09:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__PROBE_P_8%VNB 5 7 11 25
r41 7 25 1.30208e-05 $w=9.6e-06 $l=1e-09 $layer=MET1_cond $X=4.8 $Y=0.057
+ $X2=4.8 $Y2=0.058
r42 7 11 0.000742187 $w=9.6e-06 $l=5.7e-08 $layer=MET1_cond $X=4.8 $Y=0.057
+ $X2=4.8 $Y2=0
r43 5 11 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r44 5 11 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBE_P_8%VPB 4 6 14 21
r82 10 21 0.000742187 $w=9.6e-06 $l=5.7e-08 $layer=MET1_cond $X=4.8 $Y=4.07
+ $X2=4.8 $Y2=4.013
r83 10 14 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=9.36 $Y=4.07
+ $X2=9.36 $Y2=4.07
r84 9 14 594.995 $w=1.68e-07 $l=9.12e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=9.36 $Y2=4.07
r85 9 10 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r86 6 21 1.30208e-05 $w=9.6e-06 $l=1e-09 $layer=MET1_cond $X=4.8 $Y=4.012
+ $X2=4.8 $Y2=4.013
r87 4 14 18.2 $w=1.7e-07 $l=9.4024e-06 $layer=licon1_NTAP_notbjt $count=10 $X=0
+ $Y=3.985 $X2=9.36 $Y2=4.07
r88 4 9 18.2 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=10 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBE_P_8%A 3 5 7 8 10 12 15 17 19 22 24 25 26 27
+ 28 37
c74 15 0 1.75696e-19 $X=1.82 $Y=2.965
r75 36 37 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.82 $Y=1.815 $X2=2.6
+ $Y2=1.815
r76 34 36 9.0955 $w=5e-07 $l=8.5e-08 $layer=POLY_cond $X=1.735 $Y=1.815 $X2=1.82
+ $Y2=1.815
r77 27 28 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.697
+ $X2=2.16 $Y2=1.697
r78 27 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.735
+ $Y=1.73 $X2=1.735 $Y2=1.73
r79 26 27 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.697
+ $X2=1.68 $Y2=1.697
r80 25 26 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.697
+ $X2=1.2 $Y2=1.697
r81 20 37 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.6 $Y=2.065 $X2=2.6
+ $Y2=1.815
r82 20 22 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=2.6 $Y=2.065 $X2=2.6
+ $Y2=2.965
r83 17 37 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.6 $Y=1.565 $X2=2.6
+ $Y2=1.815
r84 17 19 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.6 $Y=1.565 $X2=2.6
+ $Y2=1.08
r85 13 36 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.82 $Y=2.065 $X2=1.82
+ $Y2=1.815
r86 13 15 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=1.82 $Y=2.065 $X2=1.82
+ $Y2=2.965
r87 10 36 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.82 $Y=1.565 $X2=1.82
+ $Y2=1.815
r88 10 12 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.82 $Y=1.565 $X2=1.82
+ $Y2=1.08
r89 9 24 5.30422 $w=5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.03 $Y=1.815 $X2=0.77
+ $Y2=1.815
r90 8 34 17.656 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.815 $X2=1.735
+ $Y2=1.815
r91 8 9 57.7832 $w=5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.57 $Y=1.815 $X2=1.03
+ $Y2=1.815
r92 5 24 20.4101 $w=5e-07 $l=2.54951e-07 $layer=POLY_cond $X=0.78 $Y=1.565
+ $X2=0.77 $Y2=1.815
r93 5 7 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.78 $Y=1.565 $X2=0.78
+ $Y2=1.08
r94 1 24 20.4101 $w=5e-07 $l=2.54951e-07 $layer=POLY_cond $X=0.76 $Y=2.065
+ $X2=0.77 $Y2=1.815
r95 1 3 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=0.76 $Y=2.065 $X2=0.76
+ $Y2=2.965
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBE_P_8%A_45_443# 1 2 3 4 15 17 19 22 24 26 29 31
+ 33 36 38 40 43 45 47 50 52 54 57 59 61 64 66 68 71 74 77 81 85 91 94 96 99 102
+ 103 104 107 109 119
c266 107 0 1.68957e-19 $X=2.51 $Y=1.315
c267 96 0 1.75696e-19 $X=2.51 $Y=2.095
c268 59 0 1.51336e-19 $X=8.06 $Y=2.105
c269 57 0 1.2129e-19 $X=8.06 $Y=1.08
c270 31 0 2.63163e-20 $X=4.94 $Y=2.105
r271 118 119 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=8.06 $Y=1.855
+ $X2=8.84 $Y2=1.855
r272 117 118 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.28 $Y=1.855
+ $X2=8.06 $Y2=1.855
r273 116 117 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=6.5 $Y=1.855
+ $X2=7.28 $Y2=1.855
r274 115 116 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=5.72 $Y=1.855
+ $X2=6.5 $Y2=1.855
r275 114 115 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=4.94 $Y=1.855
+ $X2=5.72 $Y2=1.855
r276 113 114 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=4.16 $Y=1.855
+ $X2=4.94 $Y2=1.855
r277 112 113 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.38 $Y=1.855
+ $X2=4.16 $Y2=1.855
r278 100 112 9.0955 $w=5e-07 $l=8.5e-08 $layer=POLY_cond $X=3.295 $Y=1.855
+ $X2=3.38 $Y2=1.855
r279 99 100 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.295
+ $Y=1.79 $X2=3.295 $Y2=1.79
r280 97 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.79
+ $X2=2.51 $Y2=1.79
r281 97 99 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.595 $Y=1.79
+ $X2=3.295 $Y2=1.79
r282 96 104 2.66603 $w=3.6e-07 $l=2.28583e-07 $layer=LI1_cond $X=2.51 $Y=2.095
+ $X2=2.32 $Y2=2.18
r283 95 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=1.955
+ $X2=2.51 $Y2=1.79
r284 95 96 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.51 $Y=1.955
+ $X2=2.51 $Y2=2.095
r285 94 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=1.625
+ $X2=2.51 $Y2=1.79
r286 93 107 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=1.4
+ $X2=2.51 $Y2=1.315
r287 93 94 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.51 $Y=1.4
+ $X2=2.51 $Y2=1.625
r288 89 107 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.21 $Y=1.315
+ $X2=2.51 $Y2=1.315
r289 89 91 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=2.21 $Y=1.23
+ $X2=2.21 $Y2=0.895
r290 85 87 22.1818 $w=5.48e-07 $l=1.02e-06 $layer=LI1_cond $X=2.32 $Y=2.34
+ $X2=2.32 $Y2=3.36
r291 83 104 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.32 $Y=2.265
+ $X2=2.32 $Y2=2.18
r292 83 85 1.63102 $w=5.48e-07 $l=7.5e-08 $layer=LI1_cond $X=2.32 $Y=2.265
+ $X2=2.32 $Y2=2.34
r293 82 103 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.435 $Y=2.18
+ $X2=0.34 $Y2=2.18
r294 81 104 4.14084 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.045 $Y=2.18
+ $X2=2.32 $Y2=2.18
r295 81 82 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=2.045 $Y=2.18
+ $X2=0.435 $Y2=2.18
r296 77 79 59.5407 $w=1.88e-07 $l=1.02e-06 $layer=LI1_cond $X=0.34 $Y=2.36
+ $X2=0.34 $Y2=3.38
r297 75 103 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.34 $Y=2.265
+ $X2=0.34 $Y2=2.18
r298 75 77 5.54545 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=0.34 $Y=2.265
+ $X2=0.34 $Y2=2.36
r299 74 103 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.34 $Y=2.095
+ $X2=0.34 $Y2=2.18
r300 74 102 36.1914 $w=1.88e-07 $l=6.2e-07 $layer=LI1_cond $X=0.34 $Y=2.095
+ $X2=0.34 $Y2=1.475
r301 69 102 5.66915 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=0.35 $Y=1.37
+ $X2=0.35 $Y2=1.475
r302 69 71 21.1255 $w=2.08e-07 $l=4e-07 $layer=LI1_cond $X=0.35 $Y=1.37 $X2=0.35
+ $Y2=0.97
r303 66 119 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.84 $Y=2.105
+ $X2=8.84 $Y2=1.855
r304 66 68 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.84 $Y=2.105 $X2=8.84
+ $Y2=2.965
r305 62 119 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.84 $Y=1.605
+ $X2=8.84 $Y2=1.855
r306 62 64 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=8.84 $Y=1.605
+ $X2=8.84 $Y2=1.08
r307 59 118 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.06 $Y=2.105
+ $X2=8.06 $Y2=1.855
r308 59 61 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.06 $Y=2.105 $X2=8.06
+ $Y2=2.965
r309 55 118 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.06 $Y=1.605
+ $X2=8.06 $Y2=1.855
r310 55 57 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=8.06 $Y=1.605
+ $X2=8.06 $Y2=1.08
r311 52 117 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.28 $Y=2.105
+ $X2=7.28 $Y2=1.855
r312 52 54 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.28 $Y=2.105 $X2=7.28
+ $Y2=2.965
r313 48 117 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.28 $Y=1.605
+ $X2=7.28 $Y2=1.855
r314 48 50 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=7.28 $Y=1.605
+ $X2=7.28 $Y2=1.08
r315 45 116 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.5 $Y=2.105 $X2=6.5
+ $Y2=1.855
r316 45 47 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.5 $Y=2.105 $X2=6.5
+ $Y2=2.965
r317 41 116 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.5 $Y=1.605 $X2=6.5
+ $Y2=1.855
r318 41 43 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=6.5 $Y=1.605 $X2=6.5
+ $Y2=1.08
r319 38 115 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.72 $Y=2.105
+ $X2=5.72 $Y2=1.855
r320 38 40 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.72 $Y=2.105 $X2=5.72
+ $Y2=2.965
r321 34 115 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.72 $Y=1.605
+ $X2=5.72 $Y2=1.855
r322 34 36 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=5.72 $Y=1.605
+ $X2=5.72 $Y2=1.08
r323 31 114 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.94 $Y=2.105
+ $X2=4.94 $Y2=1.855
r324 31 33 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.94 $Y=2.105 $X2=4.94
+ $Y2=2.965
r325 27 114 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.94 $Y=1.605
+ $X2=4.94 $Y2=1.855
r326 27 29 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.94 $Y=1.605
+ $X2=4.94 $Y2=1.08
r327 24 113 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.16 $Y=2.105
+ $X2=4.16 $Y2=1.855
r328 24 26 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.16 $Y=2.105 $X2=4.16
+ $Y2=2.965
r329 20 113 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.16 $Y=1.605
+ $X2=4.16 $Y2=1.855
r330 20 22 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.16 $Y=1.605
+ $X2=4.16 $Y2=1.08
r331 17 112 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.38 $Y=2.105
+ $X2=3.38 $Y2=1.855
r332 17 19 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.38 $Y=2.105 $X2=3.38
+ $Y2=2.965
r333 13 112 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.38 $Y=1.605
+ $X2=3.38 $Y2=1.855
r334 13 15 56.1781 $w=5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.38 $Y=1.605
+ $X2=3.38 $Y2=1.08
r335 4 87 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=2.07
+ $Y=2.215 $X2=2.21 $Y2=3.36
r336 4 85 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.07
+ $Y=2.215 $X2=2.21 $Y2=2.34
r337 3 79 300 $w=1.7e-07 $l=1.22591e-06 $layer=licon1_PDIFF $count=2 $X=0.225
+ $Y=2.215 $X2=0.35 $Y2=3.38
r338 3 77 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.225
+ $Y=2.215 $X2=0.35 $Y2=2.36
r339 2 91 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=2.07
+ $Y=0.705 $X2=2.21 $Y2=0.895
r340 1 71 91 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=2 $X=0.245
+ $Y=0.705 $X2=0.37 $Y2=0.97
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBE_P_8%VPWR 1 2 3 4 5 6 19 21 23 25 29 31 36 38
+ 40 42 43 46 56 68 80 90 105 108
r140 104 105 14.2225 $w=3.18e-07 $l=3.25e-07 $layer=LI1_cond $X=9.23 $Y=3.635
+ $X2=8.905 $Y2=3.635
r141 100 101 1.3664 $w=1.248e-06 $l=1.4e-07 $layer=LI1_cond $X=1.24 $Y=3.57
+ $X2=1.24 $Y2=3.71
r142 96 98 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=1.42 $Y=3.63
+ $X2=1.78 $Y2=3.63
r143 94 96 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.7 $Y=3.63
+ $X2=1.42 $Y2=3.63
r144 93 100 0.0976 $w=1.248e-06 $l=1e-08 $layer=LI1_cond $X=1.24 $Y=3.56
+ $X2=1.24 $Y2=3.57
r145 93 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.78 $Y=3.56
+ $X2=1.78 $Y2=3.56
r146 93 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.42 $Y=3.56
+ $X2=1.42 $Y2=3.56
r147 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.7 $Y=3.56
+ $X2=0.7 $Y2=3.56
r148 90 93 9.8576 $w=1.248e-06 $l=1.01e-06 $layer=LI1_cond $X=1.24 $Y=2.55
+ $X2=1.24 $Y2=3.56
r149 86 108 0.506755 $w=3.7e-07 $l=1.32e-06 $layer=MET1_cond $X=8.03 $Y=3.63
+ $X2=9.35 $Y2=3.63
r150 84 86 0.274492 $w=3.7e-07 $l=7.15e-07 $layer=MET1_cond $X=7.315 $Y=3.63
+ $X2=8.03 $Y2=3.63
r151 83 88 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=7.67 $Y=3.56
+ $X2=7.67 $Y2=3.57
r152 83 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.03 $Y=3.56
+ $X2=8.03 $Y2=3.56
r153 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.315 $Y=3.56
+ $X2=7.315 $Y2=3.56
r154 80 83 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=7.67 $Y=2.55
+ $X2=7.67 $Y2=3.56
r155 76 84 0.3244 $w=3.7e-07 $l=8.45e-07 $layer=MET1_cond $X=6.47 $Y=3.63
+ $X2=7.315 $Y2=3.63
r156 74 76 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=6.11 $Y=3.63
+ $X2=6.47 $Y2=3.63
r157 72 74 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=5.75 $Y=3.63
+ $X2=6.11 $Y2=3.63
r158 71 78 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=6.11 $Y=3.56
+ $X2=6.11 $Y2=3.57
r159 71 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.47 $Y=3.56
+ $X2=6.47 $Y2=3.56
r160 71 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.11 $Y=3.56
+ $X2=6.11 $Y2=3.56
r161 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=3.56
+ $X2=5.75 $Y2=3.56
r162 68 71 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=6.11 $Y=2.55
+ $X2=6.11 $Y2=3.56
r163 64 72 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=4.91 $Y=3.63
+ $X2=5.75 $Y2=3.63
r164 60 62 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=4.19 $Y=3.63
+ $X2=4.55 $Y2=3.63
r165 59 66 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=4.55 $Y=3.56
+ $X2=4.55 $Y2=3.57
r166 59 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.91 $Y=3.56
+ $X2=4.91 $Y2=3.56
r167 59 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.55 $Y=3.56
+ $X2=4.55 $Y2=3.56
r168 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.19 $Y=3.56
+ $X2=4.19 $Y2=3.56
r169 56 59 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=4.55 $Y=2.55
+ $X2=4.55 $Y2=3.56
r170 52 60 0.374308 $w=3.7e-07 $l=9.75e-07 $layer=MET1_cond $X=3.215 $Y=3.63
+ $X2=4.19 $Y2=3.63
r171 50 52 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=2.855 $Y=3.63
+ $X2=3.215 $Y2=3.63
r172 50 98 0.412698 $w=3.7e-07 $l=1.075e-06 $layer=MET1_cond $X=2.855 $Y=3.63
+ $X2=1.78 $Y2=3.63
r173 49 54 0.178519 $w=6.68e-07 $l=1e-08 $layer=LI1_cond $X=3.1 $Y=3.56 $X2=3.1
+ $Y2=3.57
r174 49 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.215 $Y=3.56
+ $X2=3.215 $Y2=3.56
r175 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.855 $Y=3.56
+ $X2=2.855 $Y2=3.56
r176 46 49 18.0304 $w=6.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.1 $Y=2.55
+ $X2=3.1 $Y2=3.56
r177 43 64 0.0422296 $w=3.7e-07 $l=1.1e-07 $layer=MET1_cond $X=4.8 $Y=3.63
+ $X2=4.91 $Y2=3.63
r178 43 62 0.0959764 $w=3.7e-07 $l=2.5e-07 $layer=MET1_cond $X=4.8 $Y=3.63
+ $X2=4.55 $Y2=3.63
r179 41 88 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=7.67 $Y=3.625
+ $X2=7.67 $Y2=3.57
r180 41 42 3.33002 $w=8.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.67 $Y=3.625
+ $X2=7.67 $Y2=3.71
r181 39 78 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6.11 $Y=3.625
+ $X2=6.11 $Y2=3.57
r182 39 40 3.33002 $w=8.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.11 $Y=3.625
+ $X2=6.11 $Y2=3.71
r183 37 66 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=4.55 $Y=3.625
+ $X2=4.55 $Y2=3.57
r184 37 38 3.33002 $w=8.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=3.625
+ $X2=4.55 $Y2=3.71
r185 35 54 0.981855 $w=6.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.1 $Y=3.625
+ $X2=3.1 $Y2=3.57
r186 35 36 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=3.625 $X2=3.1
+ $Y2=3.71
r187 31 34 21.18 $w=3.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.32 $Y=2.55 $X2=9.32
+ $Y2=3.23
r188 29 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.35 $Y=3.56
+ $X2=9.35 $Y2=3.56
r189 29 104 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=9.32 $Y=3.635
+ $X2=9.23 $Y2=3.635
r190 29 34 7.63104 $w=3.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.32 $Y=3.475
+ $X2=9.32 $Y2=3.23
r191 28 42 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=8.115 $Y=3.71
+ $X2=7.67 $Y2=3.71
r192 28 105 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.115 $Y=3.71
+ $X2=8.905 $Y2=3.71
r193 26 40 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=6.555 $Y=3.71
+ $X2=6.11 $Y2=3.71
r194 25 42 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=7.225 $Y=3.71
+ $X2=7.67 $Y2=3.71
r195 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.225 $Y=3.71
+ $X2=6.555 $Y2=3.71
r196 24 38 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=4.995 $Y=3.71
+ $X2=4.55 $Y2=3.71
r197 23 40 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=5.665 $Y=3.71
+ $X2=6.11 $Y2=3.71
r198 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.665 $Y=3.71
+ $X2=4.995 $Y2=3.71
r199 22 36 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.435 $Y=3.71
+ $X2=3.1 $Y2=3.71
r200 21 38 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=4.105 $Y=3.71
+ $X2=4.55 $Y2=3.71
r201 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.105 $Y=3.71
+ $X2=3.435 $Y2=3.71
r202 20 101 13.277 $w=1.7e-07 $l=6.25e-07 $layer=LI1_cond $X=1.865 $Y=3.71
+ $X2=1.24 $Y2=3.71
r203 19 36 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.765 $Y=3.71
+ $X2=3.1 $Y2=3.71
r204 19 20 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.765 $Y=3.71
+ $X2=1.865 $Y2=3.71
r205 6 104 600 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=1 $X=9.09
+ $Y=2.215 $X2=9.23 $Y2=3.57
r206 6 34 400 $w=1.7e-07 $l=1.08274e-06 $layer=licon1_PDIFF $count=1 $X=9.09
+ $Y=2.215 $X2=9.23 $Y2=3.23
r207 6 31 400 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=9.09
+ $Y=2.215 $X2=9.23 $Y2=2.55
r208 5 88 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=7.53
+ $Y=2.215 $X2=7.67 $Y2=3.57
r209 5 80 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=7.53
+ $Y=2.215 $X2=7.67 $Y2=2.55
r210 4 78 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=5.97
+ $Y=2.215 $X2=6.11 $Y2=3.57
r211 4 68 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=5.97
+ $Y=2.215 $X2=6.11 $Y2=2.55
r212 3 66 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=4.41
+ $Y=2.215 $X2=4.55 $Y2=3.57
r213 3 56 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=4.41
+ $Y=2.215 $X2=4.55 $Y2=2.55
r214 2 54 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=2.85
+ $Y=2.215 $X2=2.99 $Y2=3.57
r215 2 46 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=2.85
+ $Y=2.215 $X2=2.99 $Y2=2.55
r216 1 100 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=2.215 $X2=1.15 $Y2=3.57
r217 1 90 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=2.215 $X2=1.15 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBE_P_8%noxref_6 1 2 3 4 5 6 7 8 27 33 35 36 37
+ 38 41 47 49 51 55 61 63 66 68 69 70 71 74 75 76 78 79 80 81 88 91 92 94 95 98
+ 100 109
c168 109 0 9.10144e-21 $X=6.025 $Y=2.05
c169 98 0 7.9949e-21 $X=6.025 $Y=2.05
c170 94 0 2.93855e-19 $X=5.6 $Y=1.945
c171 91 0 9.21995e-21 $X=6.015 $Y=2.105
c172 88 0 1.51336e-19 $X=7.17 $Y=2.12
r173 105 109 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=5.985 $Y=2.105
+ $X2=5.985 $Y2=2.105
r174 98 109 1.705 $w=2e-07 $l=4e-07 $layer=via2 $count=2 $X=6.025 $Y=2.05
+ $X2=6.025 $Y2=2.05
r175 95 100 0.00650012 $w=3.02e-06 $l=6.75e-07 $layer=MET5_cond $X=4.8 $Y=1.945
+ $X2=4.8 $Y2=2.62
r176 94 98 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=6.025 $Y=2.05
+ $X2=6.025 $Y2=2.05
r177 94 95 0.19 $w=8e-07 $l=1.6e-06 $layer=via4_notcap2m $count=2 $X=5.6
+ $Y=1.945 $X2=5.6 $Y2=1.945
r178 91 105 0.0170272 $w=2.6e-07 $l=3e-08 $layer=MET1_cond $X=6.015 $Y=2.105
+ $X2=5.985 $Y2=2.105
r179 91 92 0.076112 $w=2.6e-07 $l=1.3e-07 $layer=MET1_cond $X=6.015 $Y=2.105
+ $X2=6.145 $Y2=2.105
r180 88 92 0.657644 $w=2.3e-07 $l=1.025e-06 $layer=MET1_cond $X=7.17 $Y=2.12
+ $X2=6.145 $Y2=2.12
r181 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.17 $Y=2.12
+ $X2=7.17 $Y2=2.12
r182 80 89 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=8.285 $Y=2.12
+ $X2=7.17 $Y2=2.12
r183 80 81 5.03717 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=8.285 $Y=2.12
+ $X2=8.625 $Y2=2.12
r184 77 89 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.055 $Y=2.12
+ $X2=7.17 $Y2=2.12
r185 77 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.055 $Y=2.12
+ $X2=6.89 $Y2=2.12
r186 74 81 2.14437 $w=4.55e-07 $l=2.64102e-07 $layer=LI1_cond $X=8.85 $Y=2.035
+ $X2=8.625 $Y2=2.12
r187 73 74 53.1126 $w=2.28e-07 $l=1.06e-06 $layer=LI1_cond $X=8.85 $Y=0.975
+ $X2=8.85 $Y2=2.035
r188 72 85 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.555 $Y=0.89
+ $X2=8.45 $Y2=0.89
r189 71 73 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=8.735 $Y=0.89
+ $X2=8.85 $Y2=0.975
r190 71 72 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.735 $Y=0.89
+ $X2=8.555 $Y2=0.89
r191 69 85 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=0.975
+ $X2=8.45 $Y2=0.89
r192 69 70 34.329 $w=2.08e-07 $l=6.5e-07 $layer=LI1_cond $X=8.45 $Y=0.975
+ $X2=8.45 $Y2=1.625
r193 66 83 8.67899 $w=6.8e-07 $l=4.7e-07 $layer=LI1_cond $X=8.625 $Y=2.89
+ $X2=8.625 $Y2=3.36
r194 66 68 9.67416 $w=6.78e-07 $l=5.5e-07 $layer=LI1_cond $X=8.625 $Y=2.89
+ $X2=8.625 $Y2=2.34
r195 65 81 2.14437 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=8.625 $Y=2.205
+ $X2=8.625 $Y2=2.12
r196 65 68 2.37457 $w=6.78e-07 $l=1.35e-07 $layer=LI1_cond $X=8.625 $Y=2.205
+ $X2=8.625 $Y2=2.34
r197 64 79 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.995 $Y=1.71
+ $X2=6.89 $Y2=1.71
r198 63 70 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.345 $Y=1.71
+ $X2=8.45 $Y2=1.625
r199 63 64 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=8.345 $Y=1.71
+ $X2=6.995 $Y2=1.71
r200 59 79 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.625
+ $X2=6.89 $Y2=1.71
r201 59 61 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=6.89 $Y=1.625
+ $X2=6.89 $Y2=0.97
r202 55 57 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=6.89 $Y=2.34
+ $X2=6.89 $Y2=3.36
r203 53 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=2.205
+ $X2=6.89 $Y2=2.12
r204 53 55 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.89 $Y=2.205
+ $X2=6.89 $Y2=2.34
r205 52 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.495 $Y=2.12
+ $X2=5.33 $Y2=2.12
r206 51 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=2.12
+ $X2=6.89 $Y2=2.12
r207 51 52 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=6.725 $Y=2.12
+ $X2=5.495 $Y2=2.12
r208 50 76 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.435 $Y=1.71
+ $X2=5.33 $Y2=1.71
r209 49 79 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.785 $Y=1.71
+ $X2=6.89 $Y2=1.71
r210 49 50 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=6.785 $Y=1.71
+ $X2=5.435 $Y2=1.71
r211 45 76 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.33 $Y=1.625
+ $X2=5.33 $Y2=1.71
r212 45 47 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=5.33 $Y=1.625
+ $X2=5.33 $Y2=0.97
r213 41 43 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=5.33 $Y=2.34
+ $X2=5.33 $Y2=3.36
r214 39 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.33 $Y=2.205
+ $X2=5.33 $Y2=2.12
r215 39 41 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.33 $Y=2.205
+ $X2=5.33 $Y2=2.34
r216 37 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=2.12
+ $X2=5.33 $Y2=2.12
r217 37 38 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=5.165 $Y=2.12
+ $X2=3.935 $Y2=2.12
r218 35 76 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.225 $Y=1.71
+ $X2=5.33 $Y2=1.71
r219 35 36 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=5.225 $Y=1.71
+ $X2=3.875 $Y2=1.71
r220 31 36 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.77 $Y=1.625
+ $X2=3.875 $Y2=1.71
r221 31 33 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=3.77 $Y=1.625
+ $X2=3.77 $Y2=0.97
r222 27 29 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3.77 $Y=2.34
+ $X2=3.77 $Y2=3.36
r223 25 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.77 $Y=2.205
+ $X2=3.935 $Y2=2.12
r224 25 27 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.77 $Y=2.205
+ $X2=3.77 $Y2=2.34
r225 8 83 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=8.31
+ $Y=2.215 $X2=8.45 $Y2=3.36
r226 8 68 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=8.31
+ $Y=2.215 $X2=8.45 $Y2=2.34
r227 7 57 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=6.75
+ $Y=2.215 $X2=6.89 $Y2=3.36
r228 7 55 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=6.75
+ $Y=2.215 $X2=6.89 $Y2=2.34
r229 6 43 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=5.19
+ $Y=2.215 $X2=5.33 $Y2=3.36
r230 6 41 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=5.19
+ $Y=2.215 $X2=5.33 $Y2=2.34
r231 5 29 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=3.63
+ $Y=2.215 $X2=3.77 $Y2=3.36
r232 5 27 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=3.63
+ $Y=2.215 $X2=3.77 $Y2=2.34
r233 4 85 91 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=2 $X=8.31
+ $Y=0.705 $X2=8.45 $Y2=0.97
r234 3 61 91 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=2 $X=6.75
+ $Y=0.705 $X2=6.89 $Y2=0.97
r235 2 47 91 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=2 $X=5.19
+ $Y=0.705 $X2=5.33 $Y2=0.97
r236 1 33 91 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=2 $X=3.63
+ $Y=0.705 $X2=3.77 $Y2=0.97
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBE_P_8%VGND 1 2 3 4 5 6 19 31 33 44 46 55 61 65
+ 71 75 81 83 85 86
c97 85 0 1.2129e-19 $X=9.42 $Y=0.465
c98 4 0 1.24898e-19 $X=5.97 $Y=0.705
r99 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.42 $Y=0.465
+ $X2=9.42 $Y2=0.465
r100 81 83 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=8.175 $Y=0.465
+ $X2=8.975 $Y2=0.465
r101 80 86 0.529789 $w=3.7e-07 $l=1.38e-06 $layer=MET1_cond $X=8.04 $Y=0.44
+ $X2=9.42 $Y2=0.44
r102 79 81 12.8638 $w=1.063e-06 $l=1.35e-07 $layer=LI1_cond $X=8.04 $Y=0.912
+ $X2=8.175 $Y2=0.912
r103 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.04 $Y=0.465
+ $X2=8.04 $Y2=0.465
r104 77 79 4.2385 $w=1.063e-06 $l=3.7e-07 $layer=LI1_cond $X=7.67 $Y=0.912
+ $X2=8.04 $Y2=0.912
r105 74 80 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.32 $Y=0.44
+ $X2=8.04 $Y2=0.44
r106 73 77 4.00939 $w=1.063e-06 $l=3.5e-07 $layer=LI1_cond $X=7.32 $Y=0.912
+ $X2=7.67 $Y2=0.912
r107 73 75 13.0929 $w=1.063e-06 $l=1.55e-07 $layer=LI1_cond $X=7.32 $Y=0.912
+ $X2=7.165 $Y2=0.912
r108 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.32 $Y=0.465
+ $X2=7.32 $Y2=0.465
r109 71 75 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.615 $Y=0.465
+ $X2=7.165 $Y2=0.465
r110 70 74 0.3244 $w=3.7e-07 $l=8.45e-07 $layer=MET1_cond $X=6.475 $Y=0.44
+ $X2=7.32 $Y2=0.44
r111 69 71 12.9211 $w=1.063e-06 $l=1.4e-07 $layer=LI1_cond $X=6.475 $Y=0.912
+ $X2=6.615 $Y2=0.912
r112 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.475 $Y=0.465
+ $X2=6.475 $Y2=0.465
r113 67 69 4.18122 $w=1.063e-06 $l=3.65e-07 $layer=LI1_cond $X=6.11 $Y=0.912
+ $X2=6.475 $Y2=0.912
r114 64 70 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.755 $Y=0.44
+ $X2=6.475 $Y2=0.44
r115 63 67 4.06667 $w=1.063e-06 $l=3.55e-07 $layer=LI1_cond $X=5.755 $Y=0.912
+ $X2=6.11 $Y2=0.912
r116 63 65 13.0357 $w=1.063e-06 $l=1.5e-07 $layer=LI1_cond $X=5.755 $Y=0.912
+ $X2=5.605 $Y2=0.912
r117 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.755 $Y=0.465
+ $X2=5.755 $Y2=0.465
r118 61 65 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.055 $Y=0.465
+ $X2=5.605 $Y2=0.465
r119 59 61 13.3793 $w=1.063e-06 $l=1.8e-07 $layer=LI1_cond $X=4.875 $Y=0.912
+ $X2=5.055 $Y2=0.912
r120 57 59 3.723 $w=1.063e-06 $l=3.25e-07 $layer=LI1_cond $X=4.55 $Y=0.912
+ $X2=4.875 $Y2=0.912
r121 53 57 4.52488 $w=1.063e-06 $l=3.95e-07 $layer=LI1_cond $X=4.155 $Y=0.912
+ $X2=4.55 $Y2=0.912
r122 53 55 12.5774 $w=1.063e-06 $l=1.1e-07 $layer=LI1_cond $X=4.155 $Y=0.912
+ $X2=4.045 $Y2=0.912
r123 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.155 $Y=0.465
+ $X2=4.155 $Y2=0.465
r124 49 54 0.28601 $w=3.7e-07 $l=7.45e-07 $layer=MET1_cond $X=3.41 $Y=0.44
+ $X2=4.155 $Y2=0.44
r125 47 49 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.69 $Y=0.44
+ $X2=3.41 $Y2=0.44
r126 46 51 7.36341 $w=7.87e-07 $l=4.75e-07 $layer=LI1_cond $X=3.05 $Y=0.465
+ $X2=3.05 $Y2=0.94
r127 46 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.41 $Y=0.465
+ $X2=3.41 $Y2=0.465
r128 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.69 $Y=0.465
+ $X2=2.69 $Y2=0.465
r129 43 47 0.32632 $w=3.7e-07 $l=8.5e-07 $layer=MET1_cond $X=1.84 $Y=0.44
+ $X2=2.69 $Y2=0.44
r130 42 44 11.907 $w=1.003e-06 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=0.882
+ $X2=1.925 $Y2=0.882
r131 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.84 $Y=0.465
+ $X2=1.84 $Y2=0.465
r132 40 42 7.64776 $w=1.003e-06 $l=6.3e-07 $layer=LI1_cond $X=1.21 $Y=0.882
+ $X2=1.84 $Y2=0.882
r133 37 43 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=0.76 $Y=0.44
+ $X2=1.84 $Y2=0.44
r134 36 40 5.46269 $w=1.003e-06 $l=4.5e-07 $layer=LI1_cond $X=0.76 $Y=0.882
+ $X2=1.21 $Y2=0.882
r135 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.76 $Y=0.465
+ $X2=0.76 $Y2=0.465
r136 33 64 0.36663 $w=3.7e-07 $l=9.55e-07 $layer=MET1_cond $X=4.8 $Y=0.44
+ $X2=5.755 $Y2=0.44
r137 33 54 0.247619 $w=3.7e-07 $l=6.45e-07 $layer=MET1_cond $X=4.8 $Y=0.44
+ $X2=4.155 $Y2=0.44
r138 33 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.875 $Y=0.465
+ $X2=4.875 $Y2=0.465
r139 29 85 5.23838 $w=2.18e-07 $l=1e-07 $layer=LI1_cond $X=9.32 $Y=0.49 $X2=9.42
+ $Y2=0.49
r140 29 83 18.6977 $w=2.18e-07 $l=3.45e-07 $layer=LI1_cond $X=9.32 $Y=0.49
+ $X2=8.975 $Y2=0.49
r141 29 31 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.32 $Y=0.6 $X2=9.32
+ $Y2=0.94
r142 22 46 10.0992 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=3.495 $Y=0.465
+ $X2=3.05 $Y2=0.465
r143 22 55 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.495 $Y=0.465
+ $X2=4.045 $Y2=0.465
r144 19 46 10.0992 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=2.605 $Y=0.465
+ $X2=3.05 $Y2=0.465
r145 19 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.605 $Y=0.465
+ $X2=1.925 $Y2=0.465
r146 6 31 91 $w=1.7e-07 $l=3.04672e-07 $layer=licon1_NDIFF $count=2 $X=9.09
+ $Y=0.705 $X2=9.25 $Y2=0.94
r147 5 77 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=7.53
+ $Y=0.705 $X2=7.67 $Y2=0.94
r148 4 67 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=5.97
+ $Y=0.705 $X2=6.11 $Y2=0.94
r149 3 57 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=4.41
+ $Y=0.705 $X2=4.55 $Y2=0.94
r150 2 51 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.705 $X2=2.99 $Y2=0.94
r151 1 40 91 $w=1.7e-07 $l=3.1229e-07 $layer=licon1_NDIFF $count=2 $X=1.03
+ $Y=0.705 $X2=1.21 $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_HVL__PROBE_P_8%X 1 3
r12 1 3 0.00103039 $w=3.02e-06 $l=1.07e-07 $layer=MET5_cond $X=4.8 $Y=2.732
+ $X2=4.8 $Y2=2.625
.ends

