* File: sky130_fd_sc_hvl__xnor2_1.pxi.spice
* Created: Fri Aug 28 09:40:51 2020
* 
x_PM_SKY130_FD_SC_HVL__XNOR2_1%VNB N_VNB_M1004_b VNB N_VNB_c_4_p VNB
+ PM_SKY130_FD_SC_HVL__XNOR2_1%VNB
x_PM_SKY130_FD_SC_HVL__XNOR2_1%VPB N_VPB_M1009_b VPB N_VPB_c_36_p VPB
+ PM_SKY130_FD_SC_HVL__XNOR2_1%VPB
x_PM_SKY130_FD_SC_HVL__XNOR2_1%B N_B_M1004_g N_B_M1009_g N_B_c_83_n N_B_c_84_n
+ N_B_c_77_n B B B B N_B_M1006_g N_B_M1001_g PM_SKY130_FD_SC_HVL__XNOR2_1%B
x_PM_SKY130_FD_SC_HVL__XNOR2_1%A N_A_M1005_g N_A_M1003_g N_A_M1008_g N_A_M1000_g
+ A A N_A_c_147_n N_A_c_148_n PM_SKY130_FD_SC_HVL__XNOR2_1%A
x_PM_SKY130_FD_SC_HVL__XNOR2_1%A_30_107# N_A_30_107#_M1004_s N_A_30_107#_M1009_d
+ N_A_30_107#_M1007_g N_A_30_107#_c_191_n N_A_30_107#_M1002_g
+ N_A_30_107#_c_193_n N_A_30_107#_c_195_n N_A_30_107#_c_214_n
+ N_A_30_107#_c_204_n N_A_30_107#_c_196_n N_A_30_107#_c_222_n
+ N_A_30_107#_c_205_n N_A_30_107#_c_197_n N_A_30_107#_c_198_n
+ N_A_30_107#_c_226_n N_A_30_107#_c_228_n N_A_30_107#_c_199_n
+ PM_SKY130_FD_SC_HVL__XNOR2_1%A_30_107#
x_PM_SKY130_FD_SC_HVL__XNOR2_1%VPWR N_VPWR_M1009_s N_VPWR_M1003_d N_VPWR_M1007_d
+ VPWR N_VPWR_c_279_n N_VPWR_c_282_n N_VPWR_c_285_n N_VPWR_c_288_n
+ PM_SKY130_FD_SC_HVL__XNOR2_1%VPWR
x_PM_SKY130_FD_SC_HVL__XNOR2_1%Y N_Y_M1002_d N_Y_M1001_d N_Y_c_327_n Y Y Y
+ N_Y_c_325_n PM_SKY130_FD_SC_HVL__XNOR2_1%Y
x_PM_SKY130_FD_SC_HVL__XNOR2_1%VGND N_VGND_M1005_d N_VGND_M1006_d VGND
+ N_VGND_c_351_n N_VGND_c_353_n N_VGND_c_355_n PM_SKY130_FD_SC_HVL__XNOR2_1%VGND
x_PM_SKY130_FD_SC_HVL__XNOR2_1%A_523_107# N_A_523_107#_M1008_d
+ N_A_523_107#_M1002_s N_A_523_107#_c_386_n N_A_523_107#_c_388_n
+ N_A_523_107#_c_389_n N_A_523_107#_c_390_n
+ PM_SKY130_FD_SC_HVL__XNOR2_1%A_523_107#
cc_1 N_VNB_M1004_b N_B_M1004_g 0.0404146f $X=-0.33 $Y=-0.265 $X2=0.86 $Y2=0.91
cc_2 N_VNB_M1004_b N_B_c_77_n 0.0480321f $X=-0.33 $Y=-0.265 $X2=0.74 $Y2=1.89
cc_3 N_VNB_M1004_b N_B_M1006_g 0.0895439f $X=-0.33 $Y=-0.265 $X2=3.155 $Y2=0.91
cc_4 N_VNB_c_4_p N_B_M1006_g 9.12303e-19 $X=0.24 $Y=0 $X2=3.155 $Y2=0.91
cc_5 N_VNB_M1004_b N_A_M1005_g 0.0367658f $X=-0.33 $Y=-0.265 $X2=0.86 $Y2=0.91
cc_6 N_VNB_M1004_b N_A_M1008_g 0.0431152f $X=-0.33 $Y=-0.265 $X2=0.74 $Y2=1.89
cc_7 N_VNB_c_4_p N_A_M1008_g 9.54195e-19 $X=0.24 $Y=0 $X2=0.74 $Y2=1.89
cc_8 N_VNB_M1004_b N_A_c_147_n 0.00393347f $X=-0.33 $Y=-0.265 $X2=3.155 $Y2=0.91
cc_9 N_VNB_M1004_b N_A_c_148_n 0.0871769f $X=-0.33 $Y=-0.265 $X2=3.155 $Y2=1.89
cc_10 N_VNB_M1004_b N_A_30_107#_c_191_n 0.0572854f $X=-0.33 $Y=-0.265 $X2=0.74
+ $Y2=1.89
cc_11 N_VNB_c_4_p N_A_30_107#_c_191_n 0.00222193f $X=0.24 $Y=0 $X2=0.74 $Y2=1.89
cc_12 N_VNB_M1004_b N_A_30_107#_c_193_n 0.0373001f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_c_4_p N_A_30_107#_c_193_n 7.68678e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_14 N_VNB_M1004_b N_A_30_107#_c_195_n 0.0262533f $X=-0.33 $Y=-0.265 $X2=2.555
+ $Y2=1.95
cc_15 N_VNB_M1004_b N_A_30_107#_c_196_n 0.00898042f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_16 N_VNB_M1004_b N_A_30_107#_c_197_n 0.0101886f $X=-0.33 $Y=-0.265 $X2=3.155
+ $Y2=1.89
cc_17 N_VNB_M1004_b N_A_30_107#_c_198_n 0.0116243f $X=-0.33 $Y=-0.265 $X2=3.09
+ $Y2=1.89
cc_18 N_VNB_M1004_b N_A_30_107#_c_199_n 0.0908536f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_19 N_VNB_M1004_b Y 0.0164354f $X=-0.33 $Y=-0.265 $X2=0.74 $Y2=2.015
cc_20 N_VNB_M1004_b N_Y_c_325_n 0.0535592f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_21 N_VNB_c_4_p N_Y_c_325_n 9.44604e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_22 N_VNB_M1004_b N_VGND_c_351_n 0.0893487f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_23 N_VNB_c_4_p N_VGND_c_351_n 0.00510042f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_24 N_VNB_M1004_b N_VGND_c_353_n 0.0285222f $X=-0.33 $Y=-0.265 $X2=3.035
+ $Y2=1.95
cc_25 N_VNB_c_4_p N_VGND_c_353_n 0.00150311f $X=0.24 $Y=0 $X2=3.035 $Y2=1.95
cc_26 N_VNB_M1004_b N_VGND_c_355_n 0.0970287f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_27 N_VNB_c_4_p N_VGND_c_355_n 0.564754f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_28 N_VNB_M1004_b N_A_523_107#_c_386_n 0.0110898f $X=-0.33 $Y=-0.265 $X2=1.565
+ $Y2=2.015
cc_29 N_VNB_c_4_p N_A_523_107#_c_386_n 8.49965e-19 $X=0.24 $Y=0 $X2=1.565
+ $Y2=2.015
cc_30 N_VNB_M1004_b N_A_523_107#_c_388_n 0.00805263f $X=-0.33 $Y=-0.265 $X2=0.74
+ $Y2=1.89
cc_31 N_VNB_M1004_b N_A_523_107#_c_389_n 0.00157567f $X=-0.33 $Y=-0.265 $X2=0.74
+ $Y2=1.89
cc_32 N_VNB_M1004_b N_A_523_107#_c_390_n 0.016955f $X=-0.33 $Y=-0.265 $X2=0.74
+ $Y2=2.015
cc_33 N_VNB_c_4_p N_A_523_107#_c_390_n 7.78491e-19 $X=0.24 $Y=0 $X2=0.74
+ $Y2=2.015
cc_34 N_VPB_M1009_b N_B_M1009_g 0.0392003f $X=-0.33 $Y=1.885 $X2=0.86 $Y2=2.965
cc_35 VPB N_B_M1009_g 0.00970178f $X=0 $Y=3.955 $X2=0.86 $Y2=2.965
cc_36 N_VPB_c_36_p N_B_M1009_g 0.0152133f $X=5.04 $Y=4.07 $X2=0.86 $Y2=2.965
cc_37 N_VPB_M1009_b N_B_c_83_n 0.00637064f $X=-0.33 $Y=1.885 $X2=1.565 $Y2=2.015
cc_38 N_VPB_M1009_b N_B_c_84_n 4.73761e-19 $X=-0.33 $Y=1.885 $X2=0.74 $Y2=1.89
cc_39 N_VPB_M1009_b N_B_c_77_n 0.021356f $X=-0.33 $Y=1.885 $X2=0.74 $Y2=1.89
cc_40 N_VPB_M1009_b B 0.010289f $X=-0.33 $Y=1.885 $X2=3.035 $Y2=1.95
cc_41 N_VPB_M1009_b N_B_M1006_g 0.0558512f $X=-0.33 $Y=1.885 $X2=3.155 $Y2=0.91
cc_42 VPB N_B_M1006_g 0.00970178f $X=0 $Y=3.955 $X2=3.155 $Y2=0.91
cc_43 N_VPB_c_36_p N_B_M1006_g 0.013715f $X=5.04 $Y=4.07 $X2=3.155 $Y2=0.91
cc_44 N_VPB_M1009_b N_A_M1003_g 0.0491254f $X=-0.33 $Y=1.885 $X2=0.86 $Y2=2.965
cc_45 VPB N_A_M1003_g 0.00970178f $X=0 $Y=3.955 $X2=0.86 $Y2=2.965
cc_46 N_VPB_c_36_p N_A_M1003_g 0.015205f $X=5.04 $Y=4.07 $X2=0.86 $Y2=2.965
cc_47 N_VPB_M1009_b N_A_M1000_g 0.0476289f $X=-0.33 $Y=1.885 $X2=0.74 $Y2=2.015
cc_48 VPB N_A_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.74 $Y2=2.015
cc_49 N_VPB_c_36_p N_A_M1000_g 0.013715f $X=5.04 $Y=4.07 $X2=0.74 $Y2=2.015
cc_50 N_VPB_M1009_b N_A_c_148_n 0.0102004f $X=-0.33 $Y=1.885 $X2=3.155 $Y2=1.89
cc_51 N_VPB_M1009_b N_A_30_107#_M1007_g 0.0465814f $X=-0.33 $Y=1.885 $X2=1.565
+ $Y2=2.015
cc_52 VPB N_A_30_107#_M1007_g 0.00970178f $X=0 $Y=3.955 $X2=1.565 $Y2=2.015
cc_53 N_VPB_c_36_p N_A_30_107#_M1007_g 0.0160007f $X=5.04 $Y=4.07 $X2=1.565
+ $Y2=2.015
cc_54 N_VPB_M1009_b N_A_30_107#_c_195_n 0.0203691f $X=-0.33 $Y=1.885 $X2=2.555
+ $Y2=1.95
cc_55 N_VPB_M1009_b N_A_30_107#_c_204_n 0.0103208f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_56 N_VPB_M1009_b N_A_30_107#_c_205_n 0.00127492f $X=-0.33 $Y=1.885 $X2=3.155
+ $Y2=0.91
cc_57 VPB N_A_30_107#_c_205_n 5.14916e-19 $X=0 $Y=3.955 $X2=3.155 $Y2=0.91
cc_58 N_VPB_c_36_p N_A_30_107#_c_205_n 0.00887752f $X=5.04 $Y=4.07 $X2=3.155
+ $Y2=0.91
cc_59 N_VPB_M1009_b N_A_30_107#_c_199_n 0.056491f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_60 N_VPB_M1009_b N_VPWR_c_279_n 0.0522351f $X=-0.33 $Y=1.885 $X2=0.74
+ $Y2=1.89
cc_61 VPB N_VPWR_c_279_n 0.00338384f $X=0 $Y=3.955 $X2=0.74 $Y2=1.89
cc_62 N_VPB_c_36_p N_VPWR_c_279_n 0.0457121f $X=5.04 $Y=4.07 $X2=0.74 $Y2=1.89
cc_63 N_VPB_M1009_b N_VPWR_c_282_n 0.00479569f $X=-0.33 $Y=1.885 $X2=3.09
+ $Y2=1.89
cc_64 VPB N_VPWR_c_282_n 0.0095202f $X=0 $Y=3.955 $X2=3.09 $Y2=1.89
cc_65 N_VPB_c_36_p N_VPWR_c_282_n 0.117146f $X=5.04 $Y=4.07 $X2=3.09 $Y2=1.89
cc_66 N_VPB_M1009_b N_VPWR_c_285_n 0.0543731f $X=-0.33 $Y=1.885 $X2=0.832
+ $Y2=1.89
cc_67 VPB N_VPWR_c_285_n 0.00229469f $X=0 $Y=3.955 $X2=0.832 $Y2=1.89
cc_68 N_VPB_c_36_p N_VPWR_c_285_n 0.0299474f $X=5.04 $Y=4.07 $X2=0.832 $Y2=1.89
cc_69 N_VPB_M1009_b N_VPWR_c_288_n 0.0532065f $X=-0.33 $Y=1.885 $X2=2.16
+ $Y2=1.962
cc_70 VPB N_VPWR_c_288_n 0.56024f $X=0 $Y=3.955 $X2=2.16 $Y2=1.962
cc_71 N_VPB_c_36_p N_VPWR_c_288_n 0.0223375f $X=5.04 $Y=4.07 $X2=2.16 $Y2=1.962
cc_72 N_VPB_M1009_b N_Y_c_327_n 0.00314504f $X=-0.33 $Y=1.885 $X2=1.565
+ $Y2=2.015
cc_73 VPB N_Y_c_327_n 8.01732e-19 $X=0 $Y=3.955 $X2=1.565 $Y2=2.015
cc_74 N_VPB_c_36_p N_Y_c_327_n 0.0130099f $X=5.04 $Y=4.07 $X2=1.565 $Y2=2.015
cc_75 N_VPB_M1009_b Y 0.0159279f $X=-0.33 $Y=1.885 $X2=0.74 $Y2=2.015
cc_76 N_B_M1004_g N_A_M1005_g 0.0529419f $X=0.86 $Y=0.91 $X2=0 $Y2=0
cc_77 N_B_c_83_n N_A_M1003_g 0.0134617f $X=1.565 $Y=2.015 $X2=0 $Y2=0
cc_78 N_B_c_77_n N_A_M1003_g 0.0246503f $X=0.74 $Y=1.89 $X2=0 $Y2=0
cc_79 B N_A_M1003_g 0.0178095f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_80 N_B_M1006_g N_A_M1008_g 0.0179528f $X=3.155 $Y=0.91 $X2=0.24 $Y2=0
cc_81 B N_A_M1000_g 0.0298754f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_82 N_B_c_83_n N_A_c_147_n 0.0329006f $X=1.565 $Y=2.015 $X2=0 $Y2=0
cc_83 N_B_c_84_n N_A_c_147_n 0.00182946f $X=0.74 $Y=1.89 $X2=0 $Y2=0
cc_84 N_B_c_77_n N_A_c_147_n 0.0100565f $X=0.74 $Y=1.89 $X2=0 $Y2=0
cc_85 B N_A_c_147_n 0.0331482f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_86 N_B_c_83_n N_A_c_148_n 0.00222753f $X=1.565 $Y=2.015 $X2=0 $Y2=0
cc_87 N_B_c_84_n N_A_c_148_n 8.43184e-19 $X=0.74 $Y=1.89 $X2=0 $Y2=0
cc_88 N_B_c_77_n N_A_c_148_n 0.0529419f $X=0.74 $Y=1.89 $X2=0 $Y2=0
cc_89 B N_A_c_148_n 0.00502263f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_90 N_B_M1006_g N_A_c_148_n 0.166218f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_91 N_B_M1004_g N_A_30_107#_c_193_n 0.0116495f $X=0.86 $Y=0.91 $X2=5.04 $Y2=0
cc_92 N_B_M1004_g N_A_30_107#_c_195_n 5.29197e-19 $X=0.86 $Y=0.91 $X2=0 $Y2=0
cc_93 N_B_M1009_g N_A_30_107#_c_195_n 0.00687793f $X=0.86 $Y=2.965 $X2=0 $Y2=0
cc_94 N_B_c_84_n N_A_30_107#_c_195_n 0.0244176f $X=0.74 $Y=1.89 $X2=0 $Y2=0
cc_95 N_B_c_77_n N_A_30_107#_c_195_n 0.02159f $X=0.74 $Y=1.89 $X2=0 $Y2=0
cc_96 N_B_M1009_g N_A_30_107#_c_214_n 0.0294576f $X=0.86 $Y=2.965 $X2=0 $Y2=0
cc_97 N_B_c_83_n N_A_30_107#_c_214_n 0.0152291f $X=1.565 $Y=2.015 $X2=0 $Y2=0
cc_98 N_B_c_84_n N_A_30_107#_c_214_n 0.0217551f $X=0.74 $Y=1.89 $X2=0 $Y2=0
cc_99 N_B_M1004_g N_A_30_107#_c_196_n 0.0309237f $X=0.86 $Y=0.91 $X2=0 $Y2=0
cc_100 N_B_c_83_n N_A_30_107#_c_196_n 0.00480923f $X=1.565 $Y=2.015 $X2=0 $Y2=0
cc_101 N_B_c_84_n N_A_30_107#_c_196_n 0.014256f $X=0.74 $Y=1.89 $X2=0 $Y2=0
cc_102 N_B_c_77_n N_A_30_107#_c_196_n 0.00216274f $X=0.74 $Y=1.89 $X2=0 $Y2=0
cc_103 B N_A_30_107#_c_196_n 0.00557851f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_104 N_B_c_83_n N_A_30_107#_c_222_n 0.0133106f $X=1.565 $Y=2.015 $X2=2.64
+ $Y2=0.058
cc_105 N_B_M1009_g N_A_30_107#_c_205_n 6.0217e-19 $X=0.86 $Y=2.965 $X2=0 $Y2=0
cc_106 B N_A_30_107#_c_197_n 0.0463162f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_107 N_B_M1006_g N_A_30_107#_c_197_n 0.0272882f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_108 B N_A_30_107#_c_226_n 0.00773858f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_109 N_B_M1006_g N_A_30_107#_c_226_n 8.43373e-19 $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_110 N_B_M1006_g N_A_30_107#_c_228_n 8.06536e-19 $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_111 B N_A_30_107#_c_199_n 0.00154768f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_112 N_B_M1006_g N_A_30_107#_c_199_n 0.0440141f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_113 N_B_M1009_g N_VPWR_c_279_n 0.0579667f $X=0.86 $Y=2.965 $X2=0 $Y2=0
cc_114 N_B_c_83_n N_VPWR_c_282_n 0.0032986f $X=1.565 $Y=2.015 $X2=0 $Y2=0
cc_115 B N_VPWR_c_282_n 0.118377f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_116 N_B_M1006_g N_VPWR_c_282_n 0.125699f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_117 N_B_M1009_g N_VPWR_c_288_n 0.00830782f $X=0.86 $Y=2.965 $X2=0 $Y2=0
cc_118 N_B_M1006_g N_VPWR_c_288_n 0.00250239f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_119 N_B_M1006_g N_Y_c_327_n 0.00976924f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_120 N_B_M1006_g Y 5.86585e-19 $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_121 N_B_M1004_g N_VGND_c_351_n 0.0519432f $X=0.86 $Y=0.91 $X2=5.04 $Y2=0
cc_122 N_B_M1006_g N_VGND_c_351_n 8.71685e-19 $X=3.155 $Y=0.91 $X2=5.04 $Y2=0
cc_123 N_B_M1006_g N_VGND_c_353_n 0.0337409f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_124 N_B_M1004_g N_VGND_c_355_n 0.00317371f $X=0.86 $Y=0.91 $X2=2.64 $Y2=0
cc_125 N_B_M1006_g N_VGND_c_355_n 0.00523812f $X=3.155 $Y=0.91 $X2=2.64 $Y2=0
cc_126 N_B_M1006_g N_A_523_107#_c_386_n 0.0161185f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_127 N_B_M1006_g N_A_523_107#_c_388_n 0.0273143f $X=3.155 $Y=0.91 $X2=0.24
+ $Y2=0
cc_128 N_B_M1006_g N_A_523_107#_c_389_n 4.40238e-19 $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_129 N_B_M1006_g N_A_523_107#_c_390_n 0.00591433f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_130 N_A_M1005_g N_A_30_107#_c_196_n 0.0256177f $X=1.57 $Y=0.91 $X2=0 $Y2=0
cc_131 N_A_M1008_g N_A_30_107#_c_196_n 0.00988482f $X=2.365 $Y=0.91 $X2=0 $Y2=0
cc_132 N_A_c_147_n N_A_30_107#_c_196_n 0.0656243f $X=1.895 $Y=1.665 $X2=0 $Y2=0
cc_133 N_A_c_148_n N_A_30_107#_c_196_n 0.00355667f $X=2.445 $Y=1.665 $X2=0 $Y2=0
cc_134 N_A_M1003_g N_A_30_107#_c_205_n 6.14203e-19 $X=1.64 $Y=2.965 $X2=0 $Y2=0
cc_135 N_A_c_148_n N_A_30_107#_c_197_n 0.0207124f $X=2.445 $Y=1.665 $X2=0 $Y2=0
cc_136 N_A_M1008_g N_A_30_107#_c_226_n 0.00895757f $X=2.365 $Y=0.91 $X2=0 $Y2=0
cc_137 N_A_c_147_n N_A_30_107#_c_226_n 0.00320067f $X=1.895 $Y=1.665 $X2=0 $Y2=0
cc_138 N_A_c_148_n N_A_30_107#_c_226_n 0.015755f $X=2.445 $Y=1.665 $X2=0 $Y2=0
cc_139 N_A_M1003_g N_VPWR_c_282_n 0.0702236f $X=1.64 $Y=2.965 $X2=0 $Y2=0
cc_140 N_A_M1000_g N_VPWR_c_282_n 0.0921962f $X=2.445 $Y=2.965 $X2=0 $Y2=0
cc_141 N_A_M1003_g N_VPWR_c_288_n 0.00780691f $X=1.64 $Y=2.965 $X2=0 $Y2=0
cc_142 N_A_M1000_g N_VPWR_c_288_n 0.00189571f $X=2.445 $Y=2.965 $X2=0 $Y2=0
cc_143 N_A_M1005_g N_VGND_c_351_n 0.0541955f $X=1.57 $Y=0.91 $X2=5.04 $Y2=0
cc_144 N_A_M1008_g N_VGND_c_351_n 0.0386531f $X=2.365 $Y=0.91 $X2=5.04 $Y2=0
cc_145 N_A_M1008_g N_VGND_c_353_n 8.27856e-19 $X=2.365 $Y=0.91 $X2=0 $Y2=0
cc_146 N_A_M1008_g N_VGND_c_355_n 0.0108997f $X=2.365 $Y=0.91 $X2=2.64 $Y2=0
cc_147 N_A_M1008_g N_A_523_107#_c_386_n 0.0129777f $X=2.365 $Y=0.91 $X2=0 $Y2=0
cc_148 N_A_M1008_g N_A_523_107#_c_389_n 0.00763703f $X=2.365 $Y=0.91 $X2=0 $Y2=0
cc_149 N_A_c_148_n N_A_523_107#_c_389_n 0.00209717f $X=2.445 $Y=1.665 $X2=0
+ $Y2=0
cc_150 N_A_30_107#_c_195_n N_VPWR_M1009_s 9.46537e-19 $X=0.235 $Y=2.28 $X2=0
+ $Y2=0
cc_151 N_A_30_107#_c_214_n N_VPWR_M1009_s 0.010058f $X=1.165 $Y=2.365 $X2=0
+ $Y2=0
cc_152 N_A_30_107#_c_204_n N_VPWR_M1009_s 7.14809e-19 $X=0.36 $Y=2.365 $X2=0
+ $Y2=0
cc_153 N_A_30_107#_c_214_n N_VPWR_c_279_n 0.0421028f $X=1.165 $Y=2.365 $X2=0
+ $Y2=0
cc_154 N_A_30_107#_c_204_n N_VPWR_c_279_n 0.0222745f $X=0.36 $Y=2.365 $X2=0
+ $Y2=0
cc_155 N_A_30_107#_c_205_n N_VPWR_c_279_n 0.0480001f $X=1.25 $Y=3.59 $X2=0 $Y2=0
cc_156 N_A_30_107#_M1007_g N_VPWR_c_282_n 0.00304668f $X=4.5 $Y=2.965 $X2=0
+ $Y2=0
cc_157 N_A_30_107#_c_205_n N_VPWR_c_282_n 0.0554137f $X=1.25 $Y=3.59 $X2=0 $Y2=0
cc_158 N_A_30_107#_c_197_n N_VPWR_c_282_n 0.010003f $X=3.65 $Y=1.54 $X2=0 $Y2=0
cc_159 N_A_30_107#_c_228_n N_VPWR_c_282_n 0.00607681f $X=3.815 $Y=1.54 $X2=0
+ $Y2=0
cc_160 N_A_30_107#_c_199_n N_VPWR_c_282_n 0.00661542f $X=4.525 $Y=1.76 $X2=0
+ $Y2=0
cc_161 N_A_30_107#_M1007_g N_VPWR_c_285_n 0.0687044f $X=4.5 $Y=2.965 $X2=0 $Y2=0
cc_162 N_A_30_107#_M1009_d N_VPWR_c_288_n 0.00442064f $X=1.11 $Y=2.215 $X2=0
+ $Y2=0
cc_163 N_A_30_107#_M1007_g N_VPWR_c_288_n 0.0116593f $X=4.5 $Y=2.965 $X2=0 $Y2=0
cc_164 N_A_30_107#_c_205_n N_VPWR_c_288_n 0.0229098f $X=1.25 $Y=3.59 $X2=0 $Y2=0
cc_165 N_A_30_107#_M1007_g N_Y_c_327_n 0.03589f $X=4.5 $Y=2.965 $X2=0 $Y2=0
cc_166 N_A_30_107#_c_199_n N_Y_c_327_n 0.00639846f $X=4.525 $Y=1.76 $X2=0 $Y2=0
cc_167 N_A_30_107#_c_228_n Y 0.00635261f $X=3.815 $Y=1.54 $X2=0 $Y2=0
cc_168 N_A_30_107#_c_199_n Y 0.0937999f $X=4.525 $Y=1.76 $X2=0 $Y2=0
cc_169 N_A_30_107#_c_191_n N_Y_c_325_n 0.031999f $X=4.525 $Y=1.435 $X2=2.64
+ $Y2=0
cc_170 N_A_30_107#_c_199_n N_Y_c_325_n 0.00789037f $X=4.525 $Y=1.76 $X2=2.64
+ $Y2=0
cc_171 N_A_30_107#_c_196_n A_222_107# 0.00103377f $X=2.24 $Y=1.315 $X2=0 $Y2=0
cc_172 N_A_30_107#_c_196_n N_VGND_M1005_d 0.00194908f $X=2.24 $Y=1.315 $X2=0
+ $Y2=0
cc_173 N_A_30_107#_c_193_n N_VGND_c_351_n 0.043841f $X=0.275 $Y=0.68 $X2=5.04
+ $Y2=0
cc_174 N_A_30_107#_c_196_n N_VGND_c_351_n 0.100407f $X=2.24 $Y=1.315 $X2=5.04
+ $Y2=0
cc_175 N_A_30_107#_c_226_n N_VGND_c_351_n 0.0126365f $X=2.325 $Y=1.315 $X2=5.04
+ $Y2=0
cc_176 N_A_30_107#_c_191_n N_VGND_c_353_n 0.00214126f $X=4.525 $Y=1.435 $X2=0
+ $Y2=0
cc_177 N_A_30_107#_M1004_s N_VGND_c_355_n 0.00243945f $X=0.15 $Y=0.535 $X2=2.64
+ $Y2=0
cc_178 N_A_30_107#_c_191_n N_VGND_c_355_n 0.030681f $X=4.525 $Y=1.435 $X2=2.64
+ $Y2=0
cc_179 N_A_30_107#_c_193_n N_VGND_c_355_n 0.0331385f $X=0.275 $Y=0.68 $X2=2.64
+ $Y2=0
cc_180 N_A_30_107#_c_196_n N_VGND_c_355_n 0.0106026f $X=2.24 $Y=1.315 $X2=2.64
+ $Y2=0
cc_181 N_A_30_107#_c_226_n N_VGND_c_355_n 5.35774e-19 $X=2.325 $Y=1.315 $X2=2.64
+ $Y2=0
cc_182 N_A_30_107#_c_191_n N_A_523_107#_c_388_n 0.00559092f $X=4.525 $Y=1.435
+ $X2=0.24 $Y2=0
cc_183 N_A_30_107#_c_197_n N_A_523_107#_c_388_n 0.04902f $X=3.65 $Y=1.54
+ $X2=0.24 $Y2=0
cc_184 N_A_30_107#_c_228_n N_A_523_107#_c_388_n 0.0244981f $X=3.815 $Y=1.54
+ $X2=0.24 $Y2=0
cc_185 N_A_30_107#_c_199_n N_A_523_107#_c_388_n 0.0194162f $X=4.525 $Y=1.76
+ $X2=0.24 $Y2=0
cc_186 N_A_30_107#_c_197_n N_A_523_107#_c_389_n 0.0215256f $X=3.65 $Y=1.54 $X2=0
+ $Y2=0
cc_187 N_A_30_107#_c_226_n N_A_523_107#_c_389_n 0.00400084f $X=2.325 $Y=1.315
+ $X2=0 $Y2=0
cc_188 N_A_30_107#_c_191_n N_A_523_107#_c_390_n 0.0174943f $X=4.525 $Y=1.435
+ $X2=0 $Y2=0
cc_189 N_VPWR_c_282_n A_539_443# 0.00109099f $X=3.76 $Y=3.59 $X2=0 $Y2=3.985
cc_190 N_VPWR_c_282_n N_Y_M1001_d 0.0398088f $X=3.76 $Y=3.59 $X2=0 $Y2=0
cc_191 N_VPWR_c_288_n N_Y_M1001_d 0.00754845f $X=4.94 $Y=3.59 $X2=0 $Y2=0
cc_192 N_VPWR_c_282_n N_Y_c_327_n 0.112155f $X=3.76 $Y=3.59 $X2=0.24 $Y2=4.07
cc_193 N_VPWR_c_285_n N_Y_c_327_n 0.101684f $X=4.89 $Y=2.34 $X2=0.24 $Y2=4.07
cc_194 N_VPWR_c_288_n N_Y_c_327_n 0.0305238f $X=4.94 $Y=3.59 $X2=0.24 $Y2=4.07
cc_195 N_VPWR_c_285_n Y 0.0467424f $X=4.89 $Y=2.34 $X2=5.04 $Y2=4.07
cc_196 N_Y_c_325_n N_VGND_c_355_n 0.0381427f $X=4.915 $Y=0.7 $X2=2.64 $Y2=0
cc_197 Y N_A_523_107#_c_388_n 0.00748492f $X=4.955 $Y=1.58 $X2=0.24 $Y2=0
cc_198 N_Y_c_325_n N_A_523_107#_c_388_n 0.00660897f $X=4.915 $Y=0.7 $X2=0.24
+ $Y2=0
cc_199 N_Y_c_325_n N_A_523_107#_c_390_n 0.0183017f $X=4.915 $Y=0.7 $X2=0 $Y2=0
cc_200 A_222_107# N_VGND_c_351_n 0.00109373f $X=1.11 $Y=0.535 $X2=0.275 $Y2=0.68
cc_201 N_VGND_c_351_n N_A_523_107#_c_386_n 0.0403541f $X=2.325 $Y=0.48 $X2=0
+ $Y2=0
cc_202 N_VGND_c_353_n N_A_523_107#_c_386_n 0.0302885f $X=3.545 $Y=0.48 $X2=0
+ $Y2=0
cc_203 N_VGND_c_355_n N_A_523_107#_c_386_n 0.0311904f $X=3.545 $Y=0.48 $X2=0
+ $Y2=0
cc_204 N_VGND_M1006_d N_A_523_107#_c_388_n 0.00614146f $X=3.405 $Y=0.535
+ $X2=0.24 $Y2=0
cc_205 N_VGND_c_353_n N_A_523_107#_c_388_n 0.0333386f $X=3.545 $Y=0.48 $X2=0.24
+ $Y2=0
cc_206 N_VGND_c_355_n N_A_523_107#_c_388_n 0.0201501f $X=3.545 $Y=0.48 $X2=0.24
+ $Y2=0
cc_207 N_VGND_c_353_n N_A_523_107#_c_390_n 0.0186295f $X=3.545 $Y=0.48 $X2=0
+ $Y2=0
cc_208 N_VGND_c_355_n N_A_523_107#_c_390_n 0.0310636f $X=3.545 $Y=0.48 $X2=0
+ $Y2=0
