* File: sky130_fd_sc_hvl__decap_8.pxi.spice
* Created: Fri Aug 28 09:33:52 2020
* 
x_PM_SKY130_FD_SC_HVL__DECAP_8%VNB N_VNB_M1001_b VNB N_VNB_c_6_p VNB
+ PM_SKY130_FD_SC_HVL__DECAP_8%VNB
x_PM_SKY130_FD_SC_HVL__DECAP_8%VPB N_VPB_M1000_b VPB N_VPB_c_15_p VPB
+ PM_SKY130_FD_SC_HVL__DECAP_8%VPB
x_PM_SKY130_FD_SC_HVL__DECAP_8%VGND N_VGND_M1001_s N_VGND_M1000_g N_VGND_M1002_g
+ N_VGND_c_31_n N_VGND_c_32_n N_VGND_c_33_n N_VGND_c_34_n VGND N_VGND_c_37_n
+ PM_SKY130_FD_SC_HVL__DECAP_8%VGND
x_PM_SKY130_FD_SC_HVL__DECAP_8%VPWR N_VPWR_M1000_s N_VPWR_c_78_n N_VPWR_M1001_g
+ N_VPWR_c_79_n N_VPWR_M1003_g N_VPWR_c_82_n N_VPWR_c_80_n N_VPWR_c_84_n
+ N_VPWR_c_81_n VPWR N_VPWR_c_86_n N_VPWR_c_89_n
+ PM_SKY130_FD_SC_HVL__DECAP_8%VPWR
cc_1 N_VNB_M1001_b N_VGND_c_31_n 0.0155366f $X=-0.33 $Y=-0.265 $X2=0.9 $Y2=1.86
cc_2 N_VNB_M1001_b N_VGND_c_32_n 0.0255963f $X=-0.33 $Y=-0.265 $X2=0.9 $Y2=1.86
cc_3 N_VNB_M1001_b N_VGND_c_33_n 0.00665656f $X=-0.33 $Y=-0.265 $X2=2.18
+ $Y2=1.86
cc_4 N_VNB_M1001_b N_VGND_c_34_n 0.0190935f $X=-0.33 $Y=-0.265 $X2=2.18 $Y2=1.86
cc_5 N_VNB_M1001_b VGND 0.110591f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0.255
cc_6 N_VNB_c_6_p VGND 0.410558f $X=0.24 $Y=0 $X2=0 $Y2=0.255
cc_7 N_VNB_M1001_b N_VGND_c_37_n 0.167103f $X=-0.33 $Y=-0.265 $X2=3.22 $Y2=0.805
cc_8 N_VNB_c_6_p N_VGND_c_37_n 0.00779523f $X=0.24 $Y=0 $X2=3.22 $Y2=0.805
cc_9 N_VNB_M1001_b N_VPWR_c_78_n 0.106291f $X=-0.33 $Y=-0.265 $X2=0.9 $Y2=2.57
cc_10 N_VNB_M1001_b N_VPWR_c_79_n 0.10885f $X=-0.33 $Y=-0.265 $X2=1.235 $Y2=2.57
cc_11 N_VNB_M1001_b N_VPWR_c_80_n 0.034203f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_12 N_VNB_M1001_b N_VPWR_c_81_n 0.0465726f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_13 N_VPB_M1000_b N_VGND_M1000_g 0.0958805f $X=-0.33 $Y=1.885 $X2=1.235
+ $Y2=3.2
cc_14 VPB N_VGND_M1000_g 0.0192119f $X=0 $Y=3.955 $X2=1.235 $Y2=3.2
cc_15 N_VPB_c_15_p N_VGND_M1000_g 0.0269766f $X=3.6 $Y=4.07 $X2=1.235 $Y2=3.2
cc_16 N_VPB_M1000_b N_VGND_M1002_g 0.0933222f $X=-0.33 $Y=1.885 $X2=2.515
+ $Y2=3.2
cc_17 VPB N_VGND_M1002_g 0.0192119f $X=0 $Y=3.955 $X2=2.515 $Y2=3.2
cc_18 N_VPB_c_15_p N_VGND_M1002_g 0.0269766f $X=3.6 $Y=4.07 $X2=2.515 $Y2=3.2
cc_19 N_VPB_M1000_b N_VGND_c_32_n 0.0777502f $X=-0.33 $Y=1.885 $X2=0.9 $Y2=1.86
cc_20 N_VPB_M1000_b N_VGND_c_34_n 0.0587107f $X=-0.33 $Y=1.885 $X2=2.18 $Y2=1.86
cc_21 N_VPB_M1000_b N_VPWR_c_82_n 0.0164247f $X=-0.33 $Y=1.885 $X2=2.515
+ $Y2=2.57
cc_22 N_VPB_M1000_b N_VPWR_c_80_n 0.0180125f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_23 N_VPB_M1000_b N_VPWR_c_84_n 0.0337872f $X=-0.33 $Y=1.885 $X2=0.9 $Y2=1.86
cc_24 N_VPB_M1000_b N_VPWR_c_81_n 0.022804f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_25 N_VPB_M1000_b N_VPWR_c_86_n 0.083949f $X=-0.33 $Y=1.885 $X2=2.965 $Y2=0.86
cc_26 VPB N_VPWR_c_86_n 0.407291f $X=0 $Y=3.955 $X2=2.965 $Y2=0.86
cc_27 N_VPB_c_15_p N_VPWR_c_86_n 0.0175711f $X=3.6 $Y=4.07 $X2=2.965 $Y2=0.86
cc_28 N_VPB_M1000_b N_VPWR_c_89_n 0.0316826f $X=-0.33 $Y=1.885 $X2=2.965
+ $Y2=0.475
cc_29 VPB N_VPWR_c_89_n 0.0118359f $X=0 $Y=3.955 $X2=2.965 $Y2=0.475
cc_30 N_VPB_c_15_p N_VPWR_c_89_n 0.133172f $X=3.6 $Y=4.07 $X2=2.965 $Y2=0.475
cc_31 N_VGND_c_31_n N_VPWR_c_78_n 0.0131031f $X=0.9 $Y=1.86 $X2=0.24 $Y2=0
cc_32 N_VGND_c_32_n N_VPWR_c_78_n 0.0159311f $X=0.9 $Y=1.86 $X2=0.24 $Y2=0
cc_33 N_VGND_c_33_n N_VPWR_c_78_n 0.0112448f $X=2.18 $Y=1.86 $X2=0.24 $Y2=0
cc_34 N_VGND_c_37_n N_VPWR_c_78_n 0.13774f $X=3.22 $Y=0.805 $X2=0.24 $Y2=0
cc_35 N_VGND_c_33_n N_VPWR_c_79_n 0.0119641f $X=2.18 $Y=1.86 $X2=0 $Y2=0
cc_36 N_VGND_c_34_n N_VPWR_c_79_n 0.0159311f $X=2.18 $Y=1.86 $X2=0 $Y2=0
cc_37 N_VGND_c_37_n N_VPWR_c_79_n 0.13774f $X=3.22 $Y=0.805 $X2=0 $Y2=0
cc_38 N_VGND_M1000_g N_VPWR_c_82_n 0.0143594f $X=1.235 $Y=3.2 $X2=0 $Y2=0
cc_39 N_VGND_c_31_n N_VPWR_c_82_n 0.0122996f $X=0.9 $Y=1.86 $X2=0 $Y2=0
cc_40 N_VGND_c_32_n N_VPWR_c_82_n 0.0185587f $X=0.9 $Y=1.86 $X2=0 $Y2=0
cc_41 N_VGND_c_33_n N_VPWR_c_82_n 0.0205243f $X=2.18 $Y=1.86 $X2=0 $Y2=0
cc_42 N_VGND_c_34_n N_VPWR_c_82_n 0.0247305f $X=2.18 $Y=1.86 $X2=0 $Y2=0
cc_43 N_VGND_c_37_n N_VPWR_c_82_n 0.0160102f $X=3.22 $Y=0.805 $X2=0 $Y2=0
cc_44 N_VGND_M1000_g N_VPWR_c_80_n 0.00443554f $X=1.235 $Y=3.2 $X2=0 $Y2=0
cc_45 N_VGND_c_31_n N_VPWR_c_80_n 0.00847063f $X=0.9 $Y=1.86 $X2=0 $Y2=0
cc_46 N_VGND_c_32_n N_VPWR_c_80_n 0.00901239f $X=0.9 $Y=1.86 $X2=0 $Y2=0
cc_47 N_VGND_c_33_n N_VPWR_c_80_n 0.00116124f $X=2.18 $Y=1.86 $X2=0 $Y2=0
cc_48 N_VGND_c_34_n N_VPWR_c_80_n 0.0195426f $X=2.18 $Y=1.86 $X2=0 $Y2=0
cc_49 N_VGND_M1002_g N_VPWR_c_84_n 0.0154983f $X=2.515 $Y=3.2 $X2=1.92 $Y2=0.057
cc_50 N_VGND_c_33_n N_VPWR_c_84_n 0.0122996f $X=2.18 $Y=1.86 $X2=1.92 $Y2=0.057
cc_51 N_VGND_c_34_n N_VPWR_c_84_n 0.0185587f $X=2.18 $Y=1.86 $X2=1.92 $Y2=0.057
cc_52 N_VGND_c_37_n N_VPWR_c_84_n 0.0160102f $X=3.22 $Y=0.805 $X2=1.92 $Y2=0.057
cc_53 N_VGND_M1002_g N_VPWR_c_81_n 0.00443554f $X=2.515 $Y=3.2 $X2=1.92
+ $Y2=0.058
cc_54 N_VGND_c_33_n N_VPWR_c_81_n 0.00847063f $X=2.18 $Y=1.86 $X2=1.92 $Y2=0.058
cc_55 N_VGND_c_34_n N_VPWR_c_81_n 0.00901239f $X=2.18 $Y=1.86 $X2=1.92 $Y2=0.058
cc_56 N_VGND_M1000_g N_VPWR_c_86_n 0.00379351f $X=1.235 $Y=3.2 $X2=0 $Y2=0
cc_57 N_VGND_M1002_g N_VPWR_c_86_n 0.00379351f $X=2.515 $Y=3.2 $X2=0 $Y2=0
cc_58 N_VGND_M1000_g N_VPWR_c_89_n 0.135664f $X=1.235 $Y=3.2 $X2=0 $Y2=0
cc_59 N_VGND_M1002_g N_VPWR_c_89_n 0.135652f $X=2.515 $Y=3.2 $X2=0 $Y2=0
cc_60 N_VGND_c_31_n N_VPWR_c_89_n 0.00892742f $X=0.9 $Y=1.86 $X2=0 $Y2=0
cc_61 N_VGND_c_33_n N_VPWR_c_89_n 0.00892742f $X=2.18 $Y=1.86 $X2=0 $Y2=0
