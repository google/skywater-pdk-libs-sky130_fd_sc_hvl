* File: sky130_fd_sc_hvl__xor2_1.spice
* Created: Wed Sep  2 09:11:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__xor2_1.pex.spice"
.subckt sky130_fd_sc_hvl__xor2_1  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1005 N_A_30_443#_M1005_d N_B_M1005_g N_VGND_M1005_s N_VNB_M1005_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.21375 PD=1.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250004 A=0.375 P=2.5 MULT=1
MM1008 N_VGND_M1008_d N_A_M1008_g N_A_30_443#_M1005_d N_VNB_M1005_b NHV L=0.5
+ W=0.75 AD=0.32625 AS=0.105 PD=1.62 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250001
+ SB=250003 A=0.375 P=2.5 MULT=1
MM1003 A_617_107# N_A_M1003_g N_VGND_M1008_d N_VNB_M1005_b NHV L=0.5 W=0.75
+ AD=0.07875 AS=0.32625 PD=0.96 PS=1.62 NRD=7.5924 NRS=89.6724 M=1 R=1.5
+ SA=250002 SB=250002 A=0.375 P=2.5 MULT=1
MM1004 N_X_M1004_d N_B_M1004_g A_617_107# N_VNB_M1005_b NHV L=0.5 W=0.75
+ AD=0.105 AS=0.07875 PD=1.03 PS=0.96 NRD=0 NRS=7.5924 M=1 R=1.5 SA=250003
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1002 N_VGND_M1002_d N_A_30_443#_M1002_g N_X_M1004_d N_VNB_M1005_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.105 PD=2.07 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250004
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1009 A_187_443# N_B_M1009_g N_A_30_443#_M1009_s N_VPB_M1009_b PHV L=0.5 W=1.5
+ AD=0.1575 AS=0.4275 PD=1.71 PS=3.57 NRD=6.3603 NRS=0 M=1 R=3 SA=250000
+ SB=250003 A=0.75 P=4 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_187_443# N_VPB_M1009_b PHV L=0.5 W=1.5
+ AD=0.3825 AS=0.1575 PD=2.01 PS=1.71 NRD=0 NRS=6.3603 M=1 R=3 SA=250001
+ SB=250002 A=0.75 P=4 MULT=1
MM1006 N_A_531_443#_M1006_d N_A_M1006_g N_VPWR_M1007_d N_VPB_M1009_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.3825 PD=1.78 PS=2.01 NRD=0 NRS=29.2803 M=1 R=3 SA=250002
+ SB=250001 A=0.75 P=4 MULT=1
MM1001 N_VPWR_M1001_d N_B_M1001_g N_A_531_443#_M1006_d N_VPB_M1009_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.21 PD=3.57 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250003
+ SB=250000 A=0.75 P=4 MULT=1
MM1000 N_A_531_443#_M1000_d N_A_30_443#_M1000_g N_X_M1000_s N_VPB_M1009_b PHV
+ L=0.5 W=1.5 AD=0.4275 AS=0.4275 PD=3.57 PS=3.57 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
DX10_noxref N_VNB_M1005_b N_VPB_M1009_b NWDIODE A=15.444 P=17.08
*
.include "sky130_fd_sc_hvl__xor2_1.pxi.spice"
*
.ends
*
*
