# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__o21a_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__o21a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.505000 4.195000 1.835000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.550000 2.785000 3.260000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.805000 2.000000 2.120000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.525000 0.380000 1.975000 ;
        RECT 0.125000 1.975000 0.595000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.550000 0.365000 1.315000 1.275000 ;
        RECT 2.785000 0.365000 3.675000 0.925000 ;
      LAYER mcon ;
        RECT 0.600000 0.395000 0.770000 0.565000 ;
        RECT 1.105000 0.395000 1.275000 0.565000 ;
        RECT 2.785000 0.395000 2.955000 0.565000 ;
        RECT 3.145000 0.395000 3.315000 0.565000 ;
        RECT 3.505000 0.395000 3.675000 0.565000 ;
      LAYER met1 ;
        RECT 0.000000 0.255000 4.320000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.320000 0.085000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.115000 4.320000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 4.320000 4.155000 ;
      LAYER mcon ;
        RECT 0.155000 3.985000 0.325000 4.155000 ;
        RECT 0.635000 3.985000 0.805000 4.155000 ;
        RECT 1.115000 3.985000 1.285000 4.155000 ;
        RECT 1.595000 3.985000 1.765000 4.155000 ;
        RECT 2.075000 3.985000 2.245000 4.155000 ;
        RECT 2.555000 3.985000 2.725000 4.155000 ;
        RECT 3.035000 3.985000 3.205000 4.155000 ;
        RECT 3.515000 3.985000 3.685000 4.155000 ;
        RECT 3.995000 3.985000 4.165000 4.155000 ;
      LAYER met1 ;
        RECT 0.000000 3.955000 4.320000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.775000 2.300000 2.025000 3.755000 ;
        RECT 2.965000 2.175000 4.230000 3.755000 ;
      LAYER mcon ;
        RECT 0.775000 3.505000 0.945000 3.675000 ;
        RECT 1.135000 3.505000 1.305000 3.675000 ;
        RECT 1.495000 3.505000 1.665000 3.675000 ;
        RECT 1.855000 3.505000 2.025000 3.675000 ;
        RECT 2.970000 3.505000 3.140000 3.675000 ;
        RECT 3.330000 3.505000 3.500000 3.675000 ;
        RECT 3.690000 3.505000 3.860000 3.675000 ;
        RECT 4.050000 3.505000 4.220000 3.675000 ;
      LAYER met1 ;
        RECT 0.000000 3.445000 4.320000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.550000 1.455000 2.375000 1.625000 ;
      RECT 0.550000 1.625000 0.835000 1.795000 ;
      RECT 1.495000 0.495000 1.825000 1.455000 ;
      RECT 2.205000 1.625000 2.375000 3.755000 ;
      RECT 2.275000 0.495000 2.605000 1.105000 ;
      RECT 2.275000 1.105000 4.185000 1.275000 ;
      RECT 3.855000 0.495000 4.185000 1.105000 ;
      RECT 3.855000 1.275000 4.185000 1.325000 ;
  END
END sky130_fd_sc_hvl__o21a_1
