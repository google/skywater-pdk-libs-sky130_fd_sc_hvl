* File: sky130_fd_sc_hvl__dfsbp_1.pxi.spice
* Created: Fri Aug 28 09:34:21 2020
* 
x_PM_SKY130_FD_SC_HVL__DFSBP_1%VNB N_VNB_M1023_b VNB N_VNB_c_2_p
+ PM_SKY130_FD_SC_HVL__DFSBP_1%VNB
x_PM_SKY130_FD_SC_HVL__DFSBP_1%VPB N_VPB_M1017_b VPB N_VPB_c_132_p
+ PM_SKY130_FD_SC_HVL__DFSBP_1%VPB
x_PM_SKY130_FD_SC_HVL__DFSBP_1%CLK N_CLK_M1023_g N_CLK_M1017_g CLK CLK CLK
+ N_CLK_c_280_n PM_SKY130_FD_SC_HVL__DFSBP_1%CLK
x_PM_SKY130_FD_SC_HVL__DFSBP_1%A_30_112# N_A_30_112#_M1023_s N_A_30_112#_M1017_s
+ N_A_30_112#_M1005_g N_A_30_112#_M1030_g N_A_30_112#_M1014_g
+ N_A_30_112#_c_325_n N_A_30_112#_M1031_g N_A_30_112#_M1028_g
+ N_A_30_112#_c_311_n N_A_30_112#_c_312_n N_A_30_112#_c_314_n
+ N_A_30_112#_c_315_n N_A_30_112#_c_420_p N_A_30_112#_c_382_n
+ N_A_30_112#_c_329_n N_A_30_112#_c_330_n N_A_30_112#_c_333_n
+ N_A_30_112#_c_336_n N_A_30_112#_c_337_n N_A_30_112#_c_338_n
+ N_A_30_112#_c_339_n N_A_30_112#_c_340_n N_A_30_112#_c_343_n
+ N_A_30_112#_c_316_n N_A_30_112#_c_317_n N_A_30_112#_c_347_n
+ N_A_30_112#_c_348_n N_A_30_112#_c_349_n N_A_30_112#_c_350_n
+ N_A_30_112#_c_353_n N_A_30_112#_c_354_n N_A_30_112#_c_451_p
+ N_A_30_112#_c_355_n N_A_30_112#_c_356_n N_A_30_112#_c_359_n
+ N_A_30_112#_c_362_n N_A_30_112#_c_363_n N_A_30_112#_c_364_n
+ N_A_30_112#_c_430_p N_A_30_112#_c_318_n N_A_30_112#_c_319_n
+ N_A_30_112#_c_320_n N_A_30_112#_c_369_n N_A_30_112#_M1000_g
+ N_A_30_112#_c_321_n PM_SKY130_FD_SC_HVL__DFSBP_1%A_30_112#
x_PM_SKY130_FD_SC_HVL__DFSBP_1%D N_D_M1022_g N_D_c_577_n D D N_D_M1001_g
+ PM_SKY130_FD_SC_HVL__DFSBP_1%D
x_PM_SKY130_FD_SC_HVL__DFSBP_1%A_339_112# N_A_339_112#_M1005_d
+ N_A_339_112#_M1030_d N_A_339_112#_c_616_n N_A_339_112#_M1012_g
+ N_A_339_112#_M1021_g N_A_339_112#_M1010_g N_A_339_112#_c_618_n
+ N_A_339_112#_c_619_n N_A_339_112#_c_620_n N_A_339_112#_c_663_n
+ N_A_339_112#_c_621_n N_A_339_112#_c_623_n N_A_339_112#_c_625_n
+ N_A_339_112#_c_711_p N_A_339_112#_c_626_n N_A_339_112#_c_638_n
+ N_A_339_112#_c_627_n N_A_339_112#_c_629_n N_A_339_112#_c_700_p
+ N_A_339_112#_c_677_n N_A_339_112#_c_678_n N_A_339_112#_c_630_n
+ N_A_339_112#_M1007_g N_A_339_112#_c_633_n
+ PM_SKY130_FD_SC_HVL__DFSBP_1%A_339_112#
x_PM_SKY130_FD_SC_HVL__DFSBP_1%A_959_83# N_A_959_83#_M1025_s N_A_959_83#_M1006_d
+ N_A_959_83#_c_796_n N_A_959_83#_M1008_g N_A_959_83#_M1009_g
+ N_A_959_83#_c_797_n N_A_959_83#_c_798_n N_A_959_83#_c_805_n
+ N_A_959_83#_c_799_n N_A_959_83#_c_806_n N_A_959_83#_c_801_n
+ N_A_959_83#_c_802_n PM_SKY130_FD_SC_HVL__DFSBP_1%A_959_83#
x_PM_SKY130_FD_SC_HVL__DFSBP_1%A_761_109# N_A_761_109#_M1014_d
+ N_A_761_109#_M1012_d N_A_761_109#_M1025_g N_A_761_109#_M1006_g
+ N_A_761_109#_M1029_g N_A_761_109#_M1033_g N_A_761_109#_c_879_n
+ N_A_761_109#_c_880_n N_A_761_109#_c_881_n N_A_761_109#_c_892_n
+ N_A_761_109#_c_893_n N_A_761_109#_c_882_n N_A_761_109#_c_883_n
+ N_A_761_109#_c_946_n N_A_761_109#_c_923_n N_A_761_109#_c_924_n
+ N_A_761_109#_c_895_n N_A_761_109#_c_884_n N_A_761_109#_c_885_n
+ PM_SKY130_FD_SC_HVL__DFSBP_1%A_761_109#
x_PM_SKY130_FD_SC_HVL__DFSBP_1%SET_B N_SET_B_c_1013_n N_SET_B_M1027_g
+ N_SET_B_c_1014_n N_SET_B_c_1015_n N_SET_B_M1032_g N_SET_B_M1004_g
+ N_SET_B_c_1016_n N_SET_B_c_1026_n N_SET_B_c_1017_n N_SET_B_c_1036_n
+ N_SET_B_c_1018_n N_SET_B_c_1042_n N_SET_B_c_1019_n N_SET_B_c_1020_n SET_B
+ SET_B N_SET_B_M1020_g N_SET_B_c_1023_n PM_SKY130_FD_SC_HVL__DFSBP_1%SET_B
x_PM_SKY130_FD_SC_HVL__DFSBP_1%A_2156_417# N_A_2156_417#_M1003_s
+ N_A_2156_417#_M1026_s N_A_2156_417#_M1011_g N_A_2156_417#_c_1127_n
+ N_A_2156_417#_M1019_g N_A_2156_417#_c_1130_n N_A_2156_417#_c_1131_n
+ N_A_2156_417#_c_1132_n N_A_2156_417#_c_1139_n N_A_2156_417#_c_1133_n
+ N_A_2156_417#_c_1140_n N_A_2156_417#_c_1141_n N_A_2156_417#_c_1134_n
+ N_A_2156_417#_c_1135_n N_A_2156_417#_c_1161_n N_A_2156_417#_c_1136_n
+ PM_SKY130_FD_SC_HVL__DFSBP_1%A_2156_417#
x_PM_SKY130_FD_SC_HVL__DFSBP_1%A_1874_543# N_A_1874_543#_M1028_d
+ N_A_1874_543#_M1000_d N_A_1874_543#_M1004_d N_A_1874_543#_M1026_g
+ N_A_1874_543#_M1003_g N_A_1874_543#_M1018_g N_A_1874_543#_M1016_g
+ N_A_1874_543#_c_1228_n N_A_1874_543#_c_1229_n N_A_1874_543#_M1024_g
+ N_A_1874_543#_M1013_g N_A_1874_543#_c_1231_n N_A_1874_543#_c_1247_n
+ N_A_1874_543#_c_1232_n N_A_1874_543#_c_1248_n N_A_1874_543#_c_1251_n
+ N_A_1874_543#_c_1233_n N_A_1874_543#_c_1234_n N_A_1874_543#_c_1278_n
+ N_A_1874_543#_c_1254_n N_A_1874_543#_c_1255_n N_A_1874_543#_c_1256_n
+ N_A_1874_543#_c_1235_n N_A_1874_543#_c_1236_n N_A_1874_543#_c_1237_n
+ N_A_1874_543#_c_1283_n N_A_1874_543#_c_1238_n
+ PM_SKY130_FD_SC_HVL__DFSBP_1%A_1874_543#
x_PM_SKY130_FD_SC_HVL__DFSBP_1%A_3129_479# N_A_3129_479#_M1013_s
+ N_A_3129_479#_M1024_s N_A_3129_479#_c_1389_n N_A_3129_479#_c_1393_n
+ N_A_3129_479#_c_1390_n N_A_3129_479#_c_1406_n N_A_3129_479#_c_1408_n
+ N_A_3129_479#_M1002_g N_A_3129_479#_M1015_g
+ PM_SKY130_FD_SC_HVL__DFSBP_1%A_3129_479#
x_PM_SKY130_FD_SC_HVL__DFSBP_1%VPWR N_VPWR_M1017_d N_VPWR_M1022_s N_VPWR_M1009_d
+ N_VPWR_M1032_d N_VPWR_M1011_d N_VPWR_M1026_d N_VPWR_M1024_d VPWR
+ N_VPWR_c_1430_n N_VPWR_c_1433_n N_VPWR_c_1436_n N_VPWR_c_1439_n
+ N_VPWR_c_1442_n N_VPWR_c_1445_n N_VPWR_c_1448_n N_VPWR_c_1451_n
+ PM_SKY130_FD_SC_HVL__DFSBP_1%VPWR
x_PM_SKY130_FD_SC_HVL__DFSBP_1%A_605_109# N_A_605_109#_M1001_d
+ N_A_605_109#_M1022_d N_A_605_109#_c_1543_n N_A_605_109#_c_1544_n
+ N_A_605_109#_c_1546_n PM_SKY130_FD_SC_HVL__DFSBP_1%A_605_109#
x_PM_SKY130_FD_SC_HVL__DFSBP_1%Q_N N_Q_N_M1016_d N_Q_N_M1018_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_1581_n PM_SKY130_FD_SC_HVL__DFSBP_1%Q_N
x_PM_SKY130_FD_SC_HVL__DFSBP_1%Q N_Q_M1002_d N_Q_M1015_d Q Q Q Q Q Q Q
+ N_Q_c_1604_n Q Q PM_SKY130_FD_SC_HVL__DFSBP_1%Q
x_PM_SKY130_FD_SC_HVL__DFSBP_1%VGND N_VGND_M1023_d N_VGND_M1001_s N_VGND_M1008_d
+ N_VGND_M1027_d N_VGND_M1020_d N_VGND_M1003_d N_VGND_M1013_d VGND
+ N_VGND_c_1619_n N_VGND_c_1621_n N_VGND_c_1623_n N_VGND_c_1625_n
+ N_VGND_c_1627_n N_VGND_c_1629_n N_VGND_c_1631_n N_VGND_c_1633_n
+ PM_SKY130_FD_SC_HVL__DFSBP_1%VGND
x_PM_SKY130_FD_SC_HVL__DFSBP_1%A_1642_107# N_A_1642_107#_M1029_d
+ N_A_1642_107#_M1010_d N_A_1642_107#_c_1740_n N_A_1642_107#_c_1741_n
+ N_A_1642_107#_c_1743_n N_A_1642_107#_c_1745_n
+ PM_SKY130_FD_SC_HVL__DFSBP_1%A_1642_107#
x_PM_SKY130_FD_SC_HVL__DFSBP_1%A_1755_153# N_A_1755_153#_M1028_s
+ N_A_1755_153#_M1019_s N_A_1755_153#_c_1774_n N_A_1755_153#_c_1782_n
+ N_A_1755_153#_c_1775_n N_A_1755_153#_c_1783_n N_A_1755_153#_c_1776_n
+ N_A_1755_153#_c_1777_n PM_SKY130_FD_SC_HVL__DFSBP_1%A_1755_153#
cc_1 N_VNB_M1023_b N_CLK_M1023_g 0.0927158f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=0.77
cc_2 N_VNB_c_2_p N_CLK_M1023_g 5.69641e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=0.77
cc_3 N_VNB_M1023_b N_CLK_c_280_n 0.0275535f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=1.795
cc_4 N_VNB_M1023_b N_A_30_112#_M1005_g 0.0461688f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.58
cc_5 N_VNB_c_2_p N_A_30_112#_M1005_g 9.31318e-19 $X=0.24 $Y=0 $X2=0.635 $Y2=1.58
cc_6 N_VNB_M1023_b N_A_30_112#_M1028_g 0.039899f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=1.795
cc_7 N_VNB_M1023_b N_A_30_112#_c_311_n 0.0749484f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_8 N_VNB_M1023_b N_A_30_112#_c_312_n 0.0337007f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_c_2_p N_A_30_112#_c_312_n 5.45461e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_10 N_VNB_M1023_b N_A_30_112#_c_314_n 0.0265337f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1023_b N_A_30_112#_c_315_n 0.013354f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_12 N_VNB_M1023_b N_A_30_112#_c_316_n 0.00139758f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1023_b N_A_30_112#_c_317_n 0.0769718f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_M1023_b N_A_30_112#_c_318_n 0.0514141f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_15 N_VNB_M1023_b N_A_30_112#_c_319_n 0.00811074f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_16 N_VNB_M1023_b N_A_30_112#_c_320_n 0.0760268f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_17 N_VNB_M1023_b N_A_30_112#_c_321_n 0.0370517f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1023_b N_D_M1001_g 0.129313f $X=-0.33 $Y=-0.265 $X2=0.675 $Y2=1.795
cc_19 N_VNB_c_2_p N_D_M1001_g 5.91139e-19 $X=0.24 $Y=0 $X2=0.675 $Y2=1.795
cc_20 N_VNB_M1023_b N_A_339_112#_c_616_n 0.0410683f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=3.035
cc_21 N_VNB_M1023_b N_A_339_112#_M1010_g 0.0869047f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=1.795
cc_22 N_VNB_M1023_b N_A_339_112#_c_618_n 0.00401943f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=1.795
cc_23 N_VNB_M1023_b N_A_339_112#_c_619_n 0.0135409f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=2.405
cc_24 N_VNB_M1023_b N_A_339_112#_c_620_n 0.0268394f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_25 N_VNB_M1023_b N_A_339_112#_c_621_n 0.117501f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_26 N_VNB_c_2_p N_A_339_112#_c_621_n 0.00552846f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_27 N_VNB_M1023_b N_A_339_112#_c_623_n 0.0135851f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_28 N_VNB_c_2_p N_A_339_112#_c_623_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_29 N_VNB_M1023_b N_A_339_112#_c_625_n 0.0528285f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_30 N_VNB_M1023_b N_A_339_112#_c_626_n 0.00421272f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_31 N_VNB_M1023_b N_A_339_112#_c_627_n 0.016759f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_32 N_VNB_c_2_p N_A_339_112#_c_627_n 7.70095e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_33 N_VNB_M1023_b N_A_339_112#_c_629_n 0.00501964f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_M1023_b N_A_339_112#_c_630_n 0.00540057f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_35 N_VNB_M1023_b N_A_339_112#_M1007_g 0.0737786f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_36 N_VNB_c_2_p N_A_339_112#_M1007_g 5.91139e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_37 N_VNB_M1023_b N_A_339_112#_c_633_n 0.0453773f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_38 N_VNB_M1023_b N_A_959_83#_c_796_n 0.0397264f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=3.035
cc_39 N_VNB_M1023_b N_A_959_83#_c_797_n 0.0101666f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=1.795
cc_40 N_VNB_M1023_b N_A_959_83#_c_798_n 0.00711312f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_41 N_VNB_M1023_b N_A_959_83#_c_799_n 0.0172883f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_42 N_VNB_c_2_p N_A_959_83#_c_799_n 7.98897e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_43 N_VNB_M1023_b N_A_959_83#_c_801_n 0.0777768f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_44 N_VNB_M1023_b N_A_959_83#_c_802_n 0.0318405f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_45 N_VNB_M1023_b N_A_761_109#_M1025_g 0.116093f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.58
cc_46 N_VNB_c_2_p N_A_761_109#_M1025_g 0.0023273f $X=0.24 $Y=0 $X2=0.635
+ $Y2=1.58
cc_47 N_VNB_M1023_b N_A_761_109#_M1006_g 0.01101f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_48 N_VNB_M1023_b N_A_761_109#_M1029_g 0.086077f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=1.795
cc_49 N_VNB_c_2_p N_A_761_109#_M1029_g 0.00209457f $X=0.24 $Y=0 $X2=0.725
+ $Y2=1.795
cc_50 N_VNB_M1023_b N_A_761_109#_c_879_n 0.00999022f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=2.035
cc_51 N_VNB_M1023_b N_A_761_109#_c_880_n 0.00331258f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_52 N_VNB_M1023_b N_A_761_109#_c_881_n 2.87267e-19 $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=2.405
cc_53 N_VNB_M1023_b N_A_761_109#_c_882_n 0.0152943f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_54 N_VNB_M1023_b N_A_761_109#_c_883_n 0.0559052f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_55 N_VNB_M1023_b N_A_761_109#_c_884_n 7.27306e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_56 N_VNB_M1023_b N_A_761_109#_c_885_n 0.0951441f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_57 N_VNB_M1023_b N_SET_B_c_1013_n 0.0369441f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=1.61
cc_58 N_VNB_M1023_b N_SET_B_c_1014_n 0.0777311f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_59 N_VNB_M1023_b N_SET_B_c_1015_n 0.042977f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.32
cc_60 N_VNB_M1023_b N_SET_B_c_1016_n 0.0056812f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_61 N_VNB_M1023_b N_SET_B_c_1017_n 0.0172719f $X=-0.33 $Y=-0.265 $X2=0.675
+ $Y2=2.32
cc_62 N_VNB_M1023_b N_SET_B_c_1018_n 0.00807836f $X=-0.33 $Y=-0.265 $X2=0.725
+ $Y2=2.405
cc_63 N_VNB_M1023_b N_SET_B_c_1019_n 0.00448299f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_64 N_VNB_M1023_b N_SET_B_c_1020_n 0.00165963f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_65 N_VNB_M1023_b SET_B 0.0060955f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_66 N_VNB_M1023_b N_SET_B_M1020_g 0.12198f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_67 N_VNB_M1023_b N_SET_B_c_1023_n 0.0067165f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_68 N_VNB_M1023_b N_A_2156_417#_c_1127_n 0.14188f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_69 N_VNB_M1023_b N_A_2156_417#_M1019_g 0.0532257f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=1.795
cc_70 N_VNB_c_2_p N_A_2156_417#_M1019_g 0.0023273f $X=0.24 $Y=0 $X2=0.675
+ $Y2=1.795
cc_71 N_VNB_M1023_b N_A_2156_417#_c_1130_n 0.0220118f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=1.795
cc_72 N_VNB_M1023_b N_A_2156_417#_c_1131_n 0.0370745f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=1.61
cc_73 N_VNB_M1023_b N_A_2156_417#_c_1132_n 0.023055f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_74 N_VNB_M1023_b N_A_2156_417#_c_1133_n 0.00897068f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_75 N_VNB_M1023_b N_A_2156_417#_c_1134_n 0.00127411f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_76 N_VNB_M1023_b N_A_2156_417#_c_1135_n 7.28287e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_77 N_VNB_M1023_b N_A_2156_417#_c_1136_n 0.00326895f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_78 N_VNB_M1023_b N_A_1874_543#_M1003_g 0.0477088f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=1.795
cc_79 N_VNB_M1023_b N_A_1874_543#_M1016_g 0.0497756f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=2.035
cc_80 N_VNB_c_2_p N_A_1874_543#_M1016_g 0.00109849f $X=0.24 $Y=0 $X2=0.725
+ $Y2=2.035
cc_81 N_VNB_M1023_b N_A_1874_543#_c_1228_n 0.0690121f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=2.405
cc_82 N_VNB_M1023_b N_A_1874_543#_c_1229_n 0.0943203f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_83 N_VNB_M1023_b N_A_1874_543#_M1013_g 0.0474107f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_84 N_VNB_M1023_b N_A_1874_543#_c_1231_n 0.0358334f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_85 N_VNB_M1023_b N_A_1874_543#_c_1232_n 0.0084621f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_86 N_VNB_M1023_b N_A_1874_543#_c_1233_n 0.00144875f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_87 N_VNB_M1023_b N_A_1874_543#_c_1234_n 0.0022139f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_88 N_VNB_M1023_b N_A_1874_543#_c_1235_n 0.00396823f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_89 N_VNB_M1023_b N_A_1874_543#_c_1236_n 0.00374841f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_90 N_VNB_M1023_b N_A_1874_543#_c_1237_n 0.0154172f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_91 N_VNB_M1023_b N_A_1874_543#_c_1238_n 0.00390273f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_92 N_VNB_M1023_b N_A_3129_479#_c_1389_n 0.0101045f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=1.58
cc_93 N_VNB_M1023_b N_A_3129_479#_c_1390_n 0.016614f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=1.795
cc_94 N_VNB_M1023_b N_A_3129_479#_M1002_g 0.0972056f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=2.035
cc_95 N_VNB_c_2_p N_A_3129_479#_M1002_g 0.00102867f $X=0.24 $Y=0 $X2=0.725
+ $Y2=2.035
cc_96 N_VNB_M1023_b N_A_605_109#_c_1543_n 0.00795734f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_97 N_VNB_M1023_b N_A_605_109#_c_1544_n 0.00685123f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=1.95
cc_98 N_VNB_M1023_b N_Q_N_c_1581_n 0.0248645f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_99 N_VNB_c_2_p N_Q_N_c_1581_n 9.54498e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_100 N_VNB_M1023_b Q 0.0377143f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_101 N_VNB_M1023_b N_Q_c_1604_n 0.033699f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_102 N_VNB_c_2_p N_Q_c_1604_n 8.31735e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_103 N_VNB_M1023_b N_VGND_c_1619_n 0.0502765f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_104 N_VNB_c_2_p N_VGND_c_1619_n 0.00269208f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_105 N_VNB_M1023_b N_VGND_c_1621_n 0.0230498f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_106 N_VNB_c_2_p N_VGND_c_1621_n 7.04867e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_107 N_VNB_M1023_b N_VGND_c_1623_n 0.0527428f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_108 N_VNB_c_2_p N_VGND_c_1623_n 0.00270208f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_109 N_VNB_M1023_b N_VGND_c_1625_n 0.0501296f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_110 N_VNB_c_2_p N_VGND_c_1625_n 0.00269683f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_111 N_VNB_M1023_b N_VGND_c_1627_n 0.0648402f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_112 N_VNB_c_2_p N_VGND_c_1627_n 0.00269683f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_113 N_VNB_M1023_b N_VGND_c_1629_n 0.0569658f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_114 N_VNB_c_2_p N_VGND_c_1629_n 0.00264916f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_115 N_VNB_M1023_b N_VGND_c_1631_n 0.0614531f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_116 N_VNB_c_2_p N_VGND_c_1631_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_117 N_VNB_M1023_b N_VGND_c_1633_n 0.266309f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_118 N_VNB_c_2_p N_VGND_c_1633_n 1.89891f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_119 N_VNB_M1023_b N_A_1642_107#_c_1740_n 0.00575656f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=1.58
cc_120 N_VNB_M1023_b N_A_1642_107#_c_1741_n 0.148929f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=2.32
cc_121 N_VNB_c_2_p N_A_1642_107#_c_1741_n 0.00739546f $X=0.24 $Y=0 $X2=0.635
+ $Y2=2.32
cc_122 N_VNB_M1023_b N_A_1642_107#_c_1743_n 0.0164759f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_123 N_VNB_c_2_p N_A_1642_107#_c_1743_n 9.24302e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_124 N_VNB_M1023_b N_A_1642_107#_c_1745_n 0.00909231f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=1.795
cc_125 N_VNB_M1023_b N_A_1755_153#_c_1774_n 0.0100837f $X=-0.33 $Y=-0.265
+ $X2=0.685 $Y2=3.035
cc_126 N_VNB_M1023_b N_A_1755_153#_c_1775_n 0.002506f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_127 N_VNB_M1023_b N_A_1755_153#_c_1776_n 0.0021201f $X=-0.33 $Y=-0.265
+ $X2=0.725 $Y2=1.795
cc_128 N_VNB_M1023_b N_A_1755_153#_c_1777_n 0.0188401f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=1.61
cc_129 N_VNB_c_2_p N_A_1755_153#_c_1777_n 8.88297e-19 $X=0.24 $Y=0 $X2=0.675
+ $Y2=1.61
cc_130 N_VPB_M1017_b N_CLK_M1017_g 0.0609627f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=3.035
cc_131 VPB N_CLK_M1017_g 8.73544e-19 $X=0 $Y=3.955 $X2=0.685 $Y2=3.035
cc_132 N_VPB_c_132_p N_CLK_M1017_g 0.00506885f $X=17.52 $Y=4.07 $X2=0.685
+ $Y2=3.035
cc_133 N_VPB_M1017_b N_CLK_c_280_n 0.0441981f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=1.795
cc_134 N_VPB_M1017_b N_A_30_112#_M1030_g 0.103052f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_135 VPB N_A_30_112#_M1030_g 7.38286e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_136 N_VPB_c_132_p N_A_30_112#_M1030_g 0.00413723f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_137 N_VPB_M1017_b N_A_30_112#_c_325_n 0.078472f $X=-0.33 $Y=1.885 $X2=0.675
+ $Y2=1.61
cc_138 N_VPB_M1017_b N_A_30_112#_c_314_n 0.0735243f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_139 VPB N_A_30_112#_c_314_n 5.28399e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_140 N_VPB_c_132_p N_A_30_112#_c_314_n 0.00522679f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_141 N_VPB_M1017_b N_A_30_112#_c_329_n 0.00104405f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_142 N_VPB_M1017_b N_A_30_112#_c_330_n 0.0130406f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_143 VPB N_A_30_112#_c_330_n 0.00234164f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_144 N_VPB_c_132_p N_A_30_112#_c_330_n 0.0450224f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_145 N_VPB_M1017_b N_A_30_112#_c_333_n 0.00262294f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_146 VPB N_A_30_112#_c_333_n 5.66512e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_147 N_VPB_c_132_p N_A_30_112#_c_333_n 0.0111824f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_148 N_VPB_M1017_b N_A_30_112#_c_336_n 0.0234826f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_149 N_VPB_M1017_b N_A_30_112#_c_337_n 0.0150627f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_150 N_VPB_M1017_b N_A_30_112#_c_338_n 0.00919848f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_151 N_VPB_M1017_b N_A_30_112#_c_339_n 0.00389099f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_152 N_VPB_M1017_b N_A_30_112#_c_340_n 0.0158523f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_153 VPB N_A_30_112#_c_340_n 0.00156736f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_154 N_VPB_c_132_p N_A_30_112#_c_340_n 0.0164773f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_155 N_VPB_M1017_b N_A_30_112#_c_343_n 0.00293407f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_156 VPB N_A_30_112#_c_343_n 3.71311e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_157 N_VPB_c_132_p N_A_30_112#_c_343_n 0.00411424f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_158 N_VPB_M1017_b N_A_30_112#_c_316_n 0.0032117f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_159 N_VPB_M1017_b N_A_30_112#_c_347_n 0.00611493f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_160 N_VPB_M1017_b N_A_30_112#_c_348_n 0.00711056f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_161 N_VPB_M1017_b N_A_30_112#_c_349_n 0.00269328f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_162 N_VPB_M1017_b N_A_30_112#_c_350_n 0.0327428f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_163 VPB N_A_30_112#_c_350_n 0.00358573f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_164 N_VPB_c_132_p N_A_30_112#_c_350_n 0.0379188f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_165 N_VPB_M1017_b N_A_30_112#_c_353_n 0.00389099f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_166 N_VPB_M1017_b N_A_30_112#_c_354_n 0.00584769f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_167 N_VPB_M1017_b N_A_30_112#_c_355_n 0.00389099f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_168 N_VPB_M1017_b N_A_30_112#_c_356_n 0.024836f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_169 VPB N_A_30_112#_c_356_n 0.00240926f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_170 N_VPB_c_132_p N_A_30_112#_c_356_n 0.0255422f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_171 N_VPB_M1017_b N_A_30_112#_c_359_n 0.00293407f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_172 VPB N_A_30_112#_c_359_n 3.71311e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_173 N_VPB_c_132_p N_A_30_112#_c_359_n 0.00411424f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_174 N_VPB_M1017_b N_A_30_112#_c_362_n 0.00713783f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_175 N_VPB_M1017_b N_A_30_112#_c_363_n 0.0202867f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_176 N_VPB_M1017_b N_A_30_112#_c_364_n 0.00419077f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_177 N_VPB_M1017_b N_A_30_112#_c_318_n 0.0551103f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_178 VPB N_A_30_112#_c_318_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_179 N_VPB_c_132_p N_A_30_112#_c_318_n 0.0193768f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_180 N_VPB_M1017_b N_A_30_112#_c_320_n 0.0015968f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_181 N_VPB_M1017_b N_A_30_112#_c_369_n 0.00178428f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_182 VPB N_A_30_112#_c_369_n 3.71311e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_183 N_VPB_c_132_p N_A_30_112#_c_369_n 0.00411424f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_184 N_VPB_M1017_b N_D_M1022_g 0.0384518f $X=-0.33 $Y=1.885 $X2=0.665 $Y2=0.77
cc_185 N_VPB_M1017_b N_D_c_577_n 0.0893846f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_186 N_VPB_M1017_b N_D_M1001_g 0.0226059f $X=-0.33 $Y=1.885 $X2=0.675
+ $Y2=1.795
cc_187 N_VPB_M1017_b N_A_339_112#_c_616_n 0.0586512f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=3.035
cc_188 N_VPB_M1017_b N_A_339_112#_M1012_g 0.0713962f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_189 N_VPB_M1017_b N_A_339_112#_M1021_g 0.0413018f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_190 N_VPB_M1017_b N_A_339_112#_c_619_n 0.0190435f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=2.405
cc_191 N_VPB_M1017_b N_A_339_112#_c_638_n 9.92399e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_192 N_VPB_M1017_b N_A_339_112#_c_630_n 0.00521088f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_193 N_VPB_M1017_b N_A_339_112#_c_633_n 0.0363617f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_194 N_VPB_M1017_b N_A_959_83#_M1009_g 0.0380299f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_195 N_VPB_M1017_b N_A_959_83#_c_798_n 0.00632536f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_196 N_VPB_M1017_b N_A_959_83#_c_805_n 0.0557302f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=2.035
cc_197 N_VPB_M1017_b N_A_959_83#_c_806_n 0.00467826f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_198 N_VPB_M1017_b N_A_959_83#_c_802_n 0.0199255f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_199 N_VPB_M1017_b N_A_761_109#_M1006_g 0.059858f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_200 N_VPB_M1017_b N_A_761_109#_M1033_g 0.0374725f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_201 VPB N_A_761_109#_M1033_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_202 N_VPB_c_132_p N_A_761_109#_M1033_g 0.013947f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_203 N_VPB_M1017_b N_A_761_109#_c_880_n 0.008452f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_204 N_VPB_M1017_b N_A_761_109#_c_881_n 0.00105331f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=2.405
cc_205 N_VPB_M1017_b N_A_761_109#_c_892_n 0.00168283f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_206 N_VPB_M1017_b N_A_761_109#_c_893_n 0.00643858f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_207 N_VPB_M1017_b N_A_761_109#_c_882_n 0.00433335f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_208 N_VPB_M1017_b N_A_761_109#_c_895_n 0.00472876f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_209 N_VPB_M1017_b N_A_761_109#_c_885_n 0.0392669f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_210 N_VPB_M1017_b N_SET_B_M1004_g 0.0457752f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=2.32
cc_211 N_VPB_M1017_b N_SET_B_c_1016_n 0.0576609f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_212 N_VPB_M1017_b N_SET_B_c_1026_n 0.124208f $X=-0.33 $Y=1.885 $X2=0.725
+ $Y2=1.795
cc_213 N_VPB_M1017_b SET_B 0.00367657f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_214 N_VPB_M1017_b N_SET_B_M1020_g 0.0212474f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_215 N_VPB_M1017_b N_SET_B_c_1023_n 0.00564436f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_216 N_VPB_M1017_b N_A_2156_417#_M1011_g 0.0377709f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=1.58
cc_217 N_VPB_M1017_b N_A_2156_417#_c_1131_n 0.0191259f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=1.61
cc_218 N_VPB_M1017_b N_A_2156_417#_c_1139_n 0.0181205f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_219 N_VPB_M1017_b N_A_2156_417#_c_1140_n 0.00375909f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_220 N_VPB_M1017_b N_A_2156_417#_c_1141_n 0.00498311f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_221 N_VPB_M1017_b N_A_1874_543#_M1026_g 0.0630298f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_222 N_VPB_M1017_b N_A_1874_543#_M1018_g 0.0600755f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=1.665
cc_223 VPB N_A_1874_543#_M1018_g 0.00970178f $X=0 $Y=3.955 $X2=0.725 $Y2=1.665
cc_224 N_VPB_c_132_p N_A_1874_543#_M1018_g 0.0160603f $X=17.52 $Y=4.07 $X2=0.725
+ $Y2=1.665
cc_225 N_VPB_M1017_b N_A_1874_543#_c_1228_n 0.0286609f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=2.405
cc_226 N_VPB_M1017_b N_A_1874_543#_c_1229_n 0.0115386f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_227 N_VPB_M1017_b N_A_1874_543#_M1024_g 0.0429403f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_228 N_VPB_M1017_b N_A_1874_543#_c_1231_n 0.0403284f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_229 N_VPB_M1017_b N_A_1874_543#_c_1247_n 0.0137115f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_230 N_VPB_M1017_b N_A_1874_543#_c_1248_n 0.0190473f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_231 VPB N_A_1874_543#_c_1248_n 0.00268541f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_232 N_VPB_c_132_p N_A_1874_543#_c_1248_n 0.044426f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_233 N_VPB_M1017_b N_A_1874_543#_c_1251_n 0.0016386f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_234 VPB N_A_1874_543#_c_1251_n 0.00106066f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_235 N_VPB_c_132_p N_A_1874_543#_c_1251_n 0.0173392f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_236 N_VPB_M1017_b N_A_1874_543#_c_1254_n 0.0173313f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_237 N_VPB_M1017_b N_A_1874_543#_c_1255_n 0.0511099f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_238 N_VPB_M1017_b N_A_1874_543#_c_1256_n 0.00770453f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_239 N_VPB_M1017_b N_A_1874_543#_c_1235_n 0.00921842f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_240 N_VPB_M1017_b N_A_1874_543#_c_1238_n 0.00801338f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_241 N_VPB_M1017_b N_A_3129_479#_c_1393_n 0.0172582f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_242 N_VPB_M1017_b N_A_3129_479#_M1002_g 0.0832267f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=2.035
cc_243 VPB N_A_3129_479#_M1002_g 9.59033e-19 $X=0 $Y=3.955 $X2=0.725 $Y2=2.035
cc_244 N_VPB_c_132_p N_A_3129_479#_M1002_g 0.00514877f $X=17.52 $Y=4.07
+ $X2=0.725 $Y2=2.035
cc_245 N_VPB_M1017_b N_VPWR_c_1430_n 0.00581737f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1430_n 0.00166879f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_247 N_VPB_c_132_p N_VPWR_c_1430_n 0.0254284f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_248 N_VPB_M1017_b N_VPWR_c_1433_n 0.016594f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1433_n 5.76128e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_250 N_VPB_c_132_p N_VPWR_c_1433_n 0.00877885f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_251 N_VPB_M1017_b N_VPWR_c_1436_n 0.0219438f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1436_n 0.00159783f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_253 N_VPB_c_132_p N_VPWR_c_1436_n 0.0243473f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_254 N_VPB_M1017_b N_VPWR_c_1439_n 0.00666465f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1439_n 0.00364355f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_256 N_VPB_c_132_p N_VPWR_c_1439_n 0.0372768f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_257 N_VPB_M1017_b N_VPWR_c_1442_n 0.0317448f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1442_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_259 N_VPB_c_132_p N_VPWR_c_1442_n 0.0409968f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_260 N_VPB_M1017_b N_VPWR_c_1445_n 0.0470438f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1445_n 0.00335473f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_262 N_VPB_c_132_p N_VPWR_c_1445_n 0.0490696f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_263 N_VPB_M1017_b N_VPWR_c_1448_n 0.037926f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1448_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_265 N_VPB_c_132_p N_VPWR_c_1448_n 0.0409968f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_266 N_VPB_M1017_b N_VPWR_c_1451_n 0.27012f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1451_n 1.89708f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_268 N_VPB_c_132_p N_VPWR_c_1451_n 0.0903761f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_269 N_VPB_M1017_b N_A_605_109#_c_1543_n 0.00723995f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_270 N_VPB_M1017_b N_A_605_109#_c_1546_n 0.00926588f $X=-0.33 $Y=1.885
+ $X2=0.725 $Y2=1.795
cc_271 N_VPB_M1017_b N_Q_N_c_1581_n 0.0263058f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_272 VPB N_Q_N_c_1581_n 0.00117356f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_273 N_VPB_c_132_p N_Q_N_c_1581_n 0.0187434f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_274 N_VPB_M1017_b Q 0.0233716f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_275 N_VPB_M1017_b Q 0.038437f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_276 N_VPB_c_132_p Q 0.00532177f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_277 N_VPB_M1017_b Q 0.00979711f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_278 N_CLK_M1023_g N_A_30_112#_M1005_g 0.0403941f $X=0.665 $Y=0.77 $X2=0 $Y2=0
cc_279 CLK N_A_30_112#_M1030_g 0.0026784f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_280 N_CLK_c_280_n N_A_30_112#_M1030_g 0.0492733f $X=0.725 $Y=1.795 $X2=0
+ $Y2=0
cc_281 N_CLK_M1023_g N_A_30_112#_c_312_n 0.0106989f $X=0.665 $Y=0.77 $X2=0 $Y2=0
cc_282 N_CLK_M1023_g N_A_30_112#_c_314_n 0.0312393f $X=0.665 $Y=0.77 $X2=0 $Y2=0
cc_283 N_CLK_M1017_g N_A_30_112#_c_314_n 0.0161658f $X=0.685 $Y=3.035 $X2=0
+ $Y2=0
cc_284 CLK N_A_30_112#_c_314_n 0.0722943f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_285 N_CLK_M1023_g N_A_30_112#_c_315_n 0.0337391f $X=0.665 $Y=0.77 $X2=0 $Y2=0
cc_286 CLK N_A_30_112#_c_315_n 0.0238596f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_287 N_CLK_c_280_n N_A_30_112#_c_315_n 7.69999e-19 $X=0.725 $Y=1.795 $X2=0
+ $Y2=0
cc_288 N_CLK_M1023_g N_A_30_112#_c_382_n 0.00134648f $X=0.665 $Y=0.77 $X2=0
+ $Y2=0
cc_289 CLK N_A_30_112#_c_382_n 0.0128147f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_290 N_CLK_c_280_n N_A_30_112#_c_382_n 9.90963e-19 $X=0.725 $Y=1.795 $X2=0
+ $Y2=0
cc_291 N_CLK_M1017_g N_A_30_112#_c_329_n 3.20227e-19 $X=0.685 $Y=3.035 $X2=0
+ $Y2=0
cc_292 CLK N_A_30_112#_c_329_n 0.0182465f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_293 N_CLK_c_280_n N_A_30_112#_c_329_n 0.00281056f $X=0.725 $Y=1.795 $X2=0
+ $Y2=0
cc_294 CLK N_A_30_112#_c_320_n 0.00136943f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_295 N_CLK_c_280_n N_A_30_112#_c_320_n 0.0144734f $X=0.725 $Y=1.795 $X2=0
+ $Y2=0
cc_296 N_CLK_M1017_g N_VPWR_c_1430_n 0.04785f $X=0.685 $Y=3.035 $X2=0 $Y2=0
cc_297 CLK N_VPWR_c_1430_n 0.0192337f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_298 N_CLK_M1017_g N_VPWR_c_1451_n 0.0139367f $X=0.685 $Y=3.035 $X2=0 $Y2=0
cc_299 N_CLK_M1023_g N_VGND_c_1619_n 0.0404474f $X=0.665 $Y=0.77 $X2=0 $Y2=0
cc_300 N_CLK_M1023_g N_VGND_c_1633_n 0.00530347f $X=0.665 $Y=0.77 $X2=0 $Y2=0
cc_301 N_A_30_112#_c_336_n N_D_M1022_g 0.00236488f $X=2.205 $Y=3.63 $X2=0 $Y2=0
cc_302 N_A_30_112#_c_339_n N_D_M1022_g 0.0286535f $X=2.94 $Y=3.355 $X2=0 $Y2=0
cc_303 N_A_30_112#_c_340_n N_D_M1022_g 0.011476f $X=3.725 $Y=3.44 $X2=0 $Y2=0
cc_304 N_A_30_112#_c_347_n N_D_M1022_g 7.07982e-19 $X=3.81 $Y=3.355 $X2=0 $Y2=0
cc_305 N_A_30_112#_c_336_n N_D_c_577_n 0.00252115f $X=2.205 $Y=3.63 $X2=0 $Y2=0
cc_306 N_A_30_112#_c_337_n N_D_c_577_n 0.0348789f $X=2.855 $Y=2.41 $X2=0 $Y2=0
cc_307 N_A_30_112#_c_339_n N_D_c_577_n 0.00457028f $X=2.94 $Y=3.355 $X2=0 $Y2=0
cc_308 N_A_30_112#_c_316_n N_D_c_577_n 3.87639e-19 $X=3.64 $Y=1.27 $X2=0 $Y2=0
cc_309 N_A_30_112#_c_317_n N_D_c_577_n 6.28282e-19 $X=3.64 $Y=1.27 $X2=0 $Y2=0
cc_310 N_A_30_112#_c_347_n N_D_c_577_n 2.78048e-19 $X=3.81 $Y=3.355 $X2=0 $Y2=0
cc_311 N_A_30_112#_c_349_n N_D_c_577_n 5.98758e-19 $X=3.895 $Y=2.31 $X2=0 $Y2=0
cc_312 N_A_30_112#_c_337_n D 0.0252735f $X=2.855 $Y=2.41 $X2=0.24 $Y2=0
cc_313 N_A_30_112#_c_317_n D 2.42417e-19 $X=3.64 $Y=1.27 $X2=0.24 $Y2=0
cc_314 N_A_30_112#_c_321_n N_D_M1001_g 0.0447945f $X=3.565 $Y=1.085 $X2=0 $Y2=0
cc_315 N_A_30_112#_c_325_n N_A_339_112#_c_616_n 0.00837546f $X=4.63 $Y=2.655
+ $X2=0 $Y2=0
cc_316 N_A_30_112#_c_316_n N_A_339_112#_c_616_n 0.0137611f $X=3.64 $Y=1.27 $X2=0
+ $Y2=0
cc_317 N_A_30_112#_c_317_n N_A_339_112#_c_616_n 0.0366018f $X=3.64 $Y=1.27 $X2=0
+ $Y2=0
cc_318 N_A_30_112#_c_348_n N_A_339_112#_c_616_n 0.00732677f $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_319 N_A_30_112#_c_325_n N_A_339_112#_M1012_g 0.0299606f $X=4.63 $Y=2.655
+ $X2=0 $Y2=0
cc_320 N_A_30_112#_c_339_n N_A_339_112#_M1012_g 5.17767e-19 $X=2.94 $Y=3.355
+ $X2=0 $Y2=0
cc_321 N_A_30_112#_c_340_n N_A_339_112#_M1012_g 0.00564101f $X=3.725 $Y=3.44
+ $X2=0 $Y2=0
cc_322 N_A_30_112#_c_316_n N_A_339_112#_M1012_g 0.00203814f $X=3.64 $Y=1.27
+ $X2=0 $Y2=0
cc_323 N_A_30_112#_c_347_n N_A_339_112#_M1012_g 0.0395784f $X=3.81 $Y=3.355
+ $X2=0 $Y2=0
cc_324 N_A_30_112#_c_348_n N_A_339_112#_M1012_g 0.0184101f $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_325 N_A_30_112#_c_349_n N_A_339_112#_M1012_g 0.0161527f $X=3.895 $Y=2.31
+ $X2=0 $Y2=0
cc_326 N_A_30_112#_c_350_n N_A_339_112#_M1012_g 0.00887434f $X=5.33 $Y=3.44
+ $X2=0 $Y2=0
cc_327 N_A_30_112#_M1028_g N_A_339_112#_M1010_g 0.0282023f $X=9.31 $Y=0.975
+ $X2=17.52 $Y2=0
cc_328 N_A_30_112#_c_318_n N_A_339_112#_M1010_g 0.00262917f $X=9.035 $Y=2.05
+ $X2=17.52 $Y2=0
cc_329 N_A_30_112#_M1005_g N_A_339_112#_c_618_n 0.00462856f $X=1.445 $Y=0.77
+ $X2=8.88 $Y2=0.057
cc_330 N_A_30_112#_c_320_n N_A_339_112#_c_618_n 0.00253702f $X=1.425 $Y=1.365
+ $X2=8.88 $Y2=0.057
cc_331 N_A_30_112#_c_420_p N_A_339_112#_c_619_n 0.00264134f $X=1.425 $Y=1.37
+ $X2=0 $Y2=0
cc_332 N_A_30_112#_c_382_n N_A_339_112#_c_619_n 0.116895f $X=1.425 $Y=1.705
+ $X2=0 $Y2=0
cc_333 N_A_30_112#_c_330_n N_A_339_112#_c_619_n 0.0115077f $X=2.12 $Y=3.715
+ $X2=0 $Y2=0
cc_334 N_A_30_112#_c_336_n N_A_339_112#_c_619_n 0.0679877f $X=2.205 $Y=3.63
+ $X2=0 $Y2=0
cc_335 N_A_30_112#_c_338_n N_A_339_112#_c_619_n 0.0137874f $X=2.29 $Y=2.41 $X2=0
+ $Y2=0
cc_336 N_A_30_112#_c_320_n N_A_339_112#_c_619_n 0.0412383f $X=1.425 $Y=1.365
+ $X2=0 $Y2=0
cc_337 N_A_30_112#_c_321_n N_A_339_112#_c_663_n 0.00135947f $X=3.565 $Y=1.085
+ $X2=0 $Y2=0
cc_338 N_A_30_112#_c_316_n N_A_339_112#_c_621_n 0.00178274f $X=3.64 $Y=1.27
+ $X2=0 $Y2=0
cc_339 N_A_30_112#_c_321_n N_A_339_112#_c_621_n 0.0198924f $X=3.565 $Y=1.085
+ $X2=0 $Y2=0
cc_340 N_A_30_112#_c_311_n N_A_339_112#_c_625_n 0.0345876f $X=9.215 $Y=1.815
+ $X2=0 $Y2=0
cc_341 N_A_30_112#_c_430_p N_A_339_112#_c_625_n 0.0159387f $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_342 N_A_30_112#_c_311_n N_A_339_112#_c_626_n 0.0100213f $X=9.215 $Y=1.815
+ $X2=0 $Y2=0
cc_343 N_A_30_112#_c_430_p N_A_339_112#_c_626_n 0.0279901f $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_344 N_A_30_112#_c_318_n N_A_339_112#_c_626_n 0.0155429f $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_345 N_A_30_112#_c_430_p N_A_339_112#_c_638_n 0.0127038f $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_346 N_A_30_112#_c_318_n N_A_339_112#_c_638_n 0.00892932f $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_347 N_A_30_112#_M1005_g N_A_339_112#_c_627_n 0.00986844f $X=1.445 $Y=0.77
+ $X2=0 $Y2=0
cc_348 N_A_30_112#_c_320_n N_A_339_112#_c_627_n 9.82694e-19 $X=1.425 $Y=1.365
+ $X2=0 $Y2=0
cc_349 N_A_30_112#_c_420_p N_A_339_112#_c_629_n 0.011522f $X=1.425 $Y=1.37 $X2=0
+ $Y2=0
cc_350 N_A_30_112#_c_320_n N_A_339_112#_c_629_n 0.00583517f $X=1.425 $Y=1.365
+ $X2=0 $Y2=0
cc_351 N_A_30_112#_c_321_n N_A_339_112#_c_677_n 0.00110836f $X=3.565 $Y=1.085
+ $X2=0 $Y2=0
cc_352 N_A_30_112#_c_318_n N_A_339_112#_c_678_n 4.52465e-19 $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_353 N_A_30_112#_c_311_n N_A_339_112#_c_630_n 0.00265748f $X=9.215 $Y=1.815
+ $X2=0 $Y2=0
cc_354 N_A_30_112#_c_317_n N_A_339_112#_M1007_g 0.0177345f $X=3.64 $Y=1.27 $X2=0
+ $Y2=0
cc_355 N_A_30_112#_c_321_n N_A_339_112#_M1007_g 0.013253f $X=3.565 $Y=1.085
+ $X2=0 $Y2=0
cc_356 N_A_30_112#_c_363_n N_A_339_112#_c_633_n 5.82642e-19 $X=8.87 $Y=2.63
+ $X2=0 $Y2=0
cc_357 N_A_30_112#_c_430_p N_A_339_112#_c_633_n 4.43783e-19 $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_358 N_A_30_112#_c_318_n N_A_339_112#_c_633_n 0.0267816f $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_359 N_A_30_112#_c_350_n N_A_959_83#_M1009_g 0.00987559f $X=5.33 $Y=3.44 $X2=0
+ $Y2=0
cc_360 N_A_30_112#_c_353_n N_A_959_83#_M1009_g 0.0287332f $X=5.415 $Y=3.355
+ $X2=0 $Y2=0
cc_361 N_A_30_112#_c_354_n N_A_959_83#_M1009_g 0.00768126f $X=6.425 $Y=2.64
+ $X2=0 $Y2=0
cc_362 N_A_30_112#_c_451_p N_A_959_83#_M1009_g 0.00418231f $X=5.5 $Y=2.64 $X2=0
+ $Y2=0
cc_363 N_A_30_112#_c_354_n N_A_959_83#_c_798_n 0.0762842f $X=6.425 $Y=2.64
+ $X2=8.88 $Y2=0
cc_364 N_A_30_112#_c_451_p N_A_959_83#_c_798_n 0.0123662f $X=5.5 $Y=2.64
+ $X2=8.88 $Y2=0
cc_365 N_A_30_112#_c_325_n N_A_959_83#_c_805_n 0.0687138f $X=4.63 $Y=2.655 $X2=0
+ $Y2=0
cc_366 N_A_30_112#_c_348_n N_A_959_83#_c_805_n 2.94613e-19 $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_367 N_A_30_112#_c_354_n N_A_959_83#_c_805_n 0.00509682f $X=6.425 $Y=2.64
+ $X2=0 $Y2=0
cc_368 N_A_30_112#_c_451_p N_A_959_83#_c_805_n 0.00344114f $X=5.5 $Y=2.64 $X2=0
+ $Y2=0
cc_369 N_A_30_112#_c_354_n N_A_959_83#_c_806_n 0.0129543f $X=6.425 $Y=2.64 $X2=0
+ $Y2=0
cc_370 N_A_30_112#_c_355_n N_A_959_83#_c_806_n 0.0160292f $X=6.51 $Y=3.355 $X2=0
+ $Y2=0
cc_371 N_A_30_112#_c_356_n N_A_959_83#_c_806_n 0.0181935f $X=7.505 $Y=3.44 $X2=0
+ $Y2=0
cc_372 N_A_30_112#_c_362_n N_A_959_83#_c_806_n 0.00782114f $X=7.59 $Y=3.355
+ $X2=0 $Y2=0
cc_373 N_A_30_112#_c_364_n N_A_959_83#_c_806_n 0.00641676f $X=7.675 $Y=2.63
+ $X2=0 $Y2=0
cc_374 N_A_30_112#_c_325_n N_A_959_83#_c_801_n 0.00108151f $X=4.63 $Y=2.655
+ $X2=0 $Y2=0
cc_375 N_A_30_112#_c_354_n N_A_761_109#_M1006_g 0.0239883f $X=6.425 $Y=2.64
+ $X2=0 $Y2=0
cc_376 N_A_30_112#_c_355_n N_A_761_109#_M1006_g 0.0288719f $X=6.51 $Y=3.355
+ $X2=0 $Y2=0
cc_377 N_A_30_112#_c_356_n N_A_761_109#_M1006_g 0.00564101f $X=7.505 $Y=3.44
+ $X2=0 $Y2=0
cc_378 N_A_30_112#_c_311_n N_A_761_109#_M1029_g 0.00940124f $X=9.215 $Y=1.815
+ $X2=17.52 $Y2=0
cc_379 N_A_30_112#_c_356_n N_A_761_109#_M1033_g 6.33268e-19 $X=7.505 $Y=3.44
+ $X2=8.88 $Y2=0
cc_380 N_A_30_112#_c_362_n N_A_761_109#_M1033_g 0.00353252f $X=7.59 $Y=3.355
+ $X2=8.88 $Y2=0
cc_381 N_A_30_112#_c_363_n N_A_761_109#_M1033_g 0.0167882f $X=8.87 $Y=2.63
+ $X2=8.88 $Y2=0
cc_382 N_A_30_112#_c_318_n N_A_761_109#_M1033_g 0.0735751f $X=9.035 $Y=2.05
+ $X2=8.88 $Y2=0
cc_383 N_A_30_112#_c_316_n N_A_761_109#_c_879_n 0.0516123f $X=3.64 $Y=1.27 $X2=0
+ $Y2=0
cc_384 N_A_30_112#_c_317_n N_A_761_109#_c_879_n 0.00523f $X=3.64 $Y=1.27 $X2=0
+ $Y2=0
cc_385 N_A_30_112#_c_321_n N_A_761_109#_c_879_n 0.00167751f $X=3.565 $Y=1.085
+ $X2=0 $Y2=0
cc_386 N_A_30_112#_c_325_n N_A_761_109#_c_880_n 0.0082024f $X=4.63 $Y=2.655
+ $X2=0 $Y2=0
cc_387 N_A_30_112#_c_348_n N_A_761_109#_c_880_n 0.0472026f $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_388 N_A_30_112#_c_316_n N_A_761_109#_c_881_n 0.0135362f $X=3.64 $Y=1.27 $X2=0
+ $Y2=0
cc_389 N_A_30_112#_c_348_n N_A_761_109#_c_881_n 0.0113249f $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_390 N_A_30_112#_c_325_n N_A_761_109#_c_892_n 0.0264704f $X=4.63 $Y=2.655
+ $X2=0 $Y2=0
cc_391 N_A_30_112#_c_348_n N_A_761_109#_c_892_n 0.0115248f $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_392 N_A_30_112#_c_350_n N_A_761_109#_c_892_n 0.0488664f $X=5.33 $Y=3.44 $X2=0
+ $Y2=0
cc_393 N_A_30_112#_c_353_n N_A_761_109#_c_892_n 0.0123662f $X=5.415 $Y=3.355
+ $X2=0 $Y2=0
cc_394 N_A_30_112#_c_325_n N_A_761_109#_c_893_n 0.00893547f $X=4.63 $Y=2.655
+ $X2=0 $Y2=0
cc_395 N_A_30_112#_c_348_n N_A_761_109#_c_893_n 0.0230013f $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_396 N_A_30_112#_c_353_n N_A_761_109#_c_893_n 0.0180635f $X=5.415 $Y=3.355
+ $X2=0 $Y2=0
cc_397 N_A_30_112#_c_451_p N_A_761_109#_c_893_n 0.0122935f $X=5.5 $Y=2.64 $X2=0
+ $Y2=0
cc_398 N_A_30_112#_c_363_n N_A_761_109#_c_882_n 0.00172781f $X=8.87 $Y=2.63
+ $X2=0 $Y2=0
cc_399 N_A_30_112#_c_364_n N_A_761_109#_c_882_n 0.00660241f $X=7.675 $Y=2.63
+ $X2=0 $Y2=0
cc_400 N_A_30_112#_c_354_n N_A_761_109#_c_883_n 4.87086e-19 $X=6.425 $Y=2.64
+ $X2=0 $Y2=0
cc_401 N_A_30_112#_c_363_n N_A_761_109#_c_923_n 0.0232944f $X=8.87 $Y=2.63 $X2=0
+ $Y2=0
cc_402 N_A_30_112#_c_321_n N_A_761_109#_c_924_n 0.00891464f $X=3.565 $Y=1.085
+ $X2=0 $Y2=0
cc_403 N_A_30_112#_c_325_n N_A_761_109#_c_895_n 0.0108751f $X=4.63 $Y=2.655
+ $X2=0 $Y2=0
cc_404 N_A_30_112#_c_347_n N_A_761_109#_c_895_n 0.0341066f $X=3.81 $Y=3.355
+ $X2=0 $Y2=0
cc_405 N_A_30_112#_c_348_n N_A_761_109#_c_895_n 0.0187562f $X=4.585 $Y=2.31
+ $X2=0 $Y2=0
cc_406 N_A_30_112#_c_350_n N_A_761_109#_c_895_n 0.0234526f $X=5.33 $Y=3.44 $X2=0
+ $Y2=0
cc_407 N_A_30_112#_c_311_n N_A_761_109#_c_885_n 0.0735751f $X=9.215 $Y=1.815
+ $X2=0 $Y2=0
cc_408 N_A_30_112#_c_363_n N_A_761_109#_c_885_n 0.0434208f $X=8.87 $Y=2.63 $X2=0
+ $Y2=0
cc_409 N_A_30_112#_c_430_p N_A_761_109#_c_885_n 0.00509103f $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_410 N_A_30_112#_c_355_n N_SET_B_c_1016_n 6.67141e-19 $X=6.51 $Y=3.355 $X2=0
+ $Y2=0
cc_411 N_A_30_112#_c_356_n N_SET_B_c_1016_n 0.0222507f $X=7.505 $Y=3.44 $X2=0
+ $Y2=0
cc_412 N_A_30_112#_c_362_n N_SET_B_c_1016_n 0.00892546f $X=7.59 $Y=3.355 $X2=0
+ $Y2=0
cc_413 N_A_30_112#_c_364_n N_SET_B_c_1016_n 0.0035729f $X=7.675 $Y=2.63 $X2=0
+ $Y2=0
cc_414 N_A_30_112#_M1028_g N_SET_B_c_1017_n 0.0212488f $X=9.31 $Y=0.975 $X2=0
+ $Y2=0
cc_415 N_A_30_112#_c_311_n N_SET_B_c_1017_n 0.0164459f $X=9.215 $Y=1.815 $X2=0
+ $Y2=0
cc_416 N_A_30_112#_c_311_n N_SET_B_c_1036_n 0.00104792f $X=9.215 $Y=1.815 $X2=0
+ $Y2=0
cc_417 N_A_30_112#_c_363_n N_A_1874_543#_c_1247_n 0.00254904f $X=8.87 $Y=2.63
+ $X2=0 $Y2=0
cc_418 N_A_30_112#_c_318_n N_A_1874_543#_c_1247_n 0.0219828f $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_419 N_A_30_112#_c_311_n N_A_1874_543#_c_1232_n 0.00383527f $X=9.215 $Y=1.815
+ $X2=0 $Y2=0
cc_420 N_A_30_112#_c_318_n N_A_1874_543#_c_1232_n 4.94323e-19 $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_421 N_A_30_112#_c_318_n N_A_1874_543#_c_1251_n 0.00473136f $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_422 N_A_30_112#_c_318_n N_A_1874_543#_c_1234_n 6.55769e-19 $X=9.035 $Y=2.05
+ $X2=0 $Y2=0
cc_423 N_A_30_112#_c_354_n N_VPWR_M1009_d 0.00663512f $X=6.425 $Y=2.64 $X2=0
+ $Y2=0
cc_424 N_A_30_112#_c_362_n N_VPWR_M1032_d 0.00743038f $X=7.59 $Y=3.355 $X2=0
+ $Y2=0
cc_425 N_A_30_112#_M1030_g N_VPWR_c_1430_n 0.0181469f $X=1.465 $Y=3.035 $X2=0
+ $Y2=0
cc_426 N_A_30_112#_c_314_n N_VPWR_c_1430_n 0.0223146f $X=0.295 $Y=2.785 $X2=0
+ $Y2=0
cc_427 N_A_30_112#_c_329_n N_VPWR_c_1430_n 0.0651976f $X=1.505 $Y=3.63 $X2=0
+ $Y2=0
cc_428 N_A_30_112#_c_333_n N_VPWR_c_1430_n 0.00523754f $X=1.59 $Y=3.715 $X2=0
+ $Y2=0
cc_429 N_A_30_112#_c_330_n N_VPWR_c_1433_n 0.00515224f $X=2.12 $Y=3.715 $X2=0
+ $Y2=0
cc_430 N_A_30_112#_c_336_n N_VPWR_c_1433_n 0.0682337f $X=2.205 $Y=3.63 $X2=0
+ $Y2=0
cc_431 N_A_30_112#_c_337_n N_VPWR_c_1433_n 0.0158625f $X=2.855 $Y=2.41 $X2=0
+ $Y2=0
cc_432 N_A_30_112#_c_339_n N_VPWR_c_1433_n 0.0470219f $X=2.94 $Y=3.355 $X2=0
+ $Y2=0
cc_433 N_A_30_112#_c_343_n N_VPWR_c_1433_n 0.0128895f $X=3.025 $Y=3.44 $X2=0
+ $Y2=0
cc_434 N_A_30_112#_c_350_n N_VPWR_c_1436_n 0.013534f $X=5.33 $Y=3.44 $X2=0 $Y2=0
cc_435 N_A_30_112#_c_353_n N_VPWR_c_1436_n 0.0339881f $X=5.415 $Y=3.355 $X2=0
+ $Y2=0
cc_436 N_A_30_112#_c_354_n N_VPWR_c_1436_n 0.0393194f $X=6.425 $Y=2.64 $X2=0
+ $Y2=0
cc_437 N_A_30_112#_c_355_n N_VPWR_c_1436_n 0.0327847f $X=6.51 $Y=3.355 $X2=0
+ $Y2=0
cc_438 N_A_30_112#_c_359_n N_VPWR_c_1436_n 0.013534f $X=6.595 $Y=3.44 $X2=0
+ $Y2=0
cc_439 N_A_30_112#_c_356_n N_VPWR_c_1439_n 0.0136632f $X=7.505 $Y=3.44 $X2=0
+ $Y2=0
cc_440 N_A_30_112#_c_362_n N_VPWR_c_1439_n 0.036368f $X=7.59 $Y=3.355 $X2=0
+ $Y2=0
cc_441 N_A_30_112#_c_363_n N_VPWR_c_1439_n 0.0669591f $X=8.87 $Y=2.63 $X2=0
+ $Y2=0
cc_442 N_A_30_112#_c_318_n N_VPWR_c_1439_n 0.0106898f $X=9.035 $Y=2.05 $X2=0
+ $Y2=0
cc_443 N_A_30_112#_M1030_g N_VPWR_c_1451_n 0.0191627f $X=1.465 $Y=3.035 $X2=0
+ $Y2=0
cc_444 N_A_30_112#_c_314_n N_VPWR_c_1451_n 0.0212012f $X=0.295 $Y=2.785 $X2=0
+ $Y2=0
cc_445 N_A_30_112#_c_329_n N_VPWR_c_1451_n 0.0190406f $X=1.505 $Y=3.63 $X2=0
+ $Y2=0
cc_446 N_A_30_112#_c_330_n N_VPWR_c_1451_n 0.0305282f $X=2.12 $Y=3.715 $X2=0
+ $Y2=0
cc_447 N_A_30_112#_c_333_n N_VPWR_c_1451_n 0.00770899f $X=1.59 $Y=3.715 $X2=0
+ $Y2=0
cc_448 N_A_30_112#_c_336_n N_VPWR_c_1451_n 0.0192692f $X=2.205 $Y=3.63 $X2=0
+ $Y2=0
cc_449 N_A_30_112#_c_340_n N_VPWR_c_1451_n 0.0323939f $X=3.725 $Y=3.44 $X2=0
+ $Y2=0
cc_450 N_A_30_112#_c_343_n N_VPWR_c_1451_n 0.0101279f $X=3.025 $Y=3.44 $X2=0
+ $Y2=0
cc_451 N_A_30_112#_c_350_n N_VPWR_c_1451_n 0.0702119f $X=5.33 $Y=3.44 $X2=0
+ $Y2=0
cc_452 N_A_30_112#_c_356_n N_VPWR_c_1451_n 0.0587115f $X=7.505 $Y=3.44 $X2=0
+ $Y2=0
cc_453 N_A_30_112#_c_359_n N_VPWR_c_1451_n 0.0101279f $X=6.595 $Y=3.44 $X2=0
+ $Y2=0
cc_454 N_A_30_112#_c_318_n N_VPWR_c_1451_n 0.0310979f $X=9.035 $Y=2.05 $X2=0
+ $Y2=0
cc_455 N_A_30_112#_c_369_n N_VPWR_c_1451_n 0.00928606f $X=3.81 $Y=3.44 $X2=0
+ $Y2=0
cc_456 N_A_30_112#_c_337_n N_A_605_109#_c_1543_n 0.0123662f $X=2.855 $Y=2.41
+ $X2=0 $Y2=0
cc_457 N_A_30_112#_c_339_n N_A_605_109#_c_1543_n 0.0115568f $X=2.94 $Y=3.355
+ $X2=0 $Y2=0
cc_458 N_A_30_112#_c_316_n N_A_605_109#_c_1543_n 0.0758454f $X=3.64 $Y=1.27
+ $X2=0 $Y2=0
cc_459 N_A_30_112#_c_317_n N_A_605_109#_c_1543_n 0.0202672f $X=3.64 $Y=1.27
+ $X2=0 $Y2=0
cc_460 N_A_30_112#_c_347_n N_A_605_109#_c_1543_n 0.0117018f $X=3.81 $Y=3.355
+ $X2=0 $Y2=0
cc_461 N_A_30_112#_c_349_n N_A_605_109#_c_1543_n 0.0136213f $X=3.895 $Y=2.31
+ $X2=0 $Y2=0
cc_462 N_A_30_112#_c_321_n N_A_605_109#_c_1543_n 0.00273793f $X=3.565 $Y=1.085
+ $X2=0 $Y2=0
cc_463 N_A_30_112#_c_321_n N_A_605_109#_c_1544_n 0.0123147f $X=3.565 $Y=1.085
+ $X2=0.24 $Y2=0
cc_464 N_A_30_112#_c_339_n N_A_605_109#_c_1546_n 0.0342204f $X=2.94 $Y=3.355
+ $X2=17.52 $Y2=0
cc_465 N_A_30_112#_c_340_n N_A_605_109#_c_1546_n 0.0239177f $X=3.725 $Y=3.44
+ $X2=17.52 $Y2=0
cc_466 N_A_30_112#_c_347_n N_A_605_109#_c_1546_n 0.0192587f $X=3.81 $Y=3.355
+ $X2=17.52 $Y2=0
cc_467 N_A_30_112#_M1005_g N_VGND_c_1619_n 0.036391f $X=1.445 $Y=0.77 $X2=0
+ $Y2=0
cc_468 N_A_30_112#_c_312_n N_VGND_c_1619_n 0.0216845f $X=0.275 $Y=0.77 $X2=0
+ $Y2=0
cc_469 N_A_30_112#_c_315_n N_VGND_c_1619_n 0.0529258f $X=1.26 $Y=1.285 $X2=0
+ $Y2=0
cc_470 N_A_30_112#_c_420_p N_VGND_c_1619_n 0.0178729f $X=1.425 $Y=1.37 $X2=0
+ $Y2=0
cc_471 N_A_30_112#_M1005_g N_VGND_c_1621_n 0.00253062f $X=1.445 $Y=0.77 $X2=0
+ $Y2=0
cc_472 N_A_30_112#_M1023_s N_VGND_c_1633_n 7.41599e-19 $X=0.15 $Y=0.56 $X2=0
+ $Y2=0
cc_473 N_A_30_112#_M1005_g N_VGND_c_1633_n 0.00935568f $X=1.445 $Y=0.77 $X2=0
+ $Y2=0
cc_474 N_A_30_112#_M1028_g N_VGND_c_1633_n 0.0173305f $X=9.31 $Y=0.975 $X2=0
+ $Y2=0
cc_475 N_A_30_112#_c_312_n N_VGND_c_1633_n 0.0238999f $X=0.275 $Y=0.77 $X2=0
+ $Y2=0
cc_476 N_A_30_112#_c_315_n N_VGND_c_1633_n 0.00686642f $X=1.26 $Y=1.285 $X2=0
+ $Y2=0
cc_477 N_A_30_112#_c_420_p N_VGND_c_1633_n 0.00398203f $X=1.425 $Y=1.37 $X2=0
+ $Y2=0
cc_478 N_A_30_112#_c_316_n N_VGND_c_1633_n 0.00376901f $X=3.64 $Y=1.27 $X2=0
+ $Y2=0
cc_479 N_A_30_112#_c_319_n N_VGND_c_1633_n 7.63525e-19 $X=0.245 $Y=1.285 $X2=0
+ $Y2=0
cc_480 N_A_30_112#_c_321_n N_VGND_c_1633_n 0.0157659f $X=3.565 $Y=1.085 $X2=0
+ $Y2=0
cc_481 N_A_30_112#_M1028_g N_A_1642_107#_c_1740_n 0.00313088f $X=9.31 $Y=0.975
+ $X2=0 $Y2=0
cc_482 N_A_30_112#_M1028_g N_A_1642_107#_c_1741_n 0.0143115f $X=9.31 $Y=0.975
+ $X2=0.24 $Y2=0
cc_483 N_A_30_112#_M1028_g N_A_1755_153#_c_1774_n 0.0277836f $X=9.31 $Y=0.975
+ $X2=0 $Y2=0
cc_484 N_A_30_112#_c_311_n N_A_1755_153#_c_1774_n 8.20966e-19 $X=9.215 $Y=1.815
+ $X2=0 $Y2=0
cc_485 N_D_c_577_n N_A_339_112#_c_616_n 0.0180507f $X=3.07 $Y=2.335 $X2=0 $Y2=0
cc_486 N_D_M1001_g N_A_339_112#_c_616_n 0.00131588f $X=2.775 $Y=0.755 $X2=0
+ $Y2=0
cc_487 N_D_M1022_g N_A_339_112#_M1012_g 0.0180507f $X=3.07 $Y=2.925 $X2=0 $Y2=0
cc_488 N_D_c_577_n N_A_339_112#_c_619_n 6.22594e-19 $X=3.07 $Y=2.335 $X2=0 $Y2=0
cc_489 D N_A_339_112#_c_619_n 0.0186335f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_490 N_D_M1001_g N_A_339_112#_c_619_n 0.0206336f $X=2.775 $Y=0.755 $X2=0 $Y2=0
cc_491 D N_A_339_112#_c_620_n 0.0225889f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_492 N_D_M1001_g N_A_339_112#_c_620_n 0.0184443f $X=2.775 $Y=0.755 $X2=0 $Y2=0
cc_493 N_D_M1001_g N_A_339_112#_c_663_n 0.0302836f $X=2.775 $Y=0.755 $X2=0 $Y2=0
cc_494 N_D_M1001_g N_A_339_112#_c_621_n 0.00864871f $X=2.775 $Y=0.755 $X2=0
+ $Y2=0
cc_495 N_D_M1001_g N_A_339_112#_c_623_n 0.0033683f $X=2.775 $Y=0.755 $X2=0 $Y2=0
cc_496 N_D_M1001_g N_A_339_112#_c_627_n 0.00418102f $X=2.775 $Y=0.755 $X2=0
+ $Y2=0
cc_497 N_D_M1022_g N_VPWR_c_1433_n 0.0149779f $X=3.07 $Y=2.925 $X2=0 $Y2=0
cc_498 N_D_c_577_n N_VPWR_c_1433_n 0.00449573f $X=3.07 $Y=2.335 $X2=0 $Y2=0
cc_499 N_D_M1022_g N_VPWR_c_1451_n 0.00113143f $X=3.07 $Y=2.925 $X2=0 $Y2=0
cc_500 N_D_M1022_g N_A_605_109#_c_1543_n 0.00333266f $X=3.07 $Y=2.925 $X2=0
+ $Y2=0
cc_501 N_D_c_577_n N_A_605_109#_c_1543_n 0.0231863f $X=3.07 $Y=2.335 $X2=0 $Y2=0
cc_502 D N_A_605_109#_c_1543_n 0.0287249f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_503 N_D_M1001_g N_A_605_109#_c_1543_n 0.0154712f $X=2.775 $Y=0.755 $X2=0
+ $Y2=0
cc_504 N_D_M1001_g N_A_605_109#_c_1544_n 0.0082888f $X=2.775 $Y=0.755 $X2=0.24
+ $Y2=0
cc_505 N_D_M1022_g N_A_605_109#_c_1546_n 0.0147803f $X=3.07 $Y=2.925 $X2=17.52
+ $Y2=0
cc_506 N_D_M1001_g N_VGND_c_1621_n 0.00415578f $X=2.775 $Y=0.755 $X2=0 $Y2=0
cc_507 N_D_M1001_g N_VGND_c_1633_n 0.01471f $X=2.775 $Y=0.755 $X2=0 $Y2=0
cc_508 N_A_339_112#_c_677_n N_A_959_83#_c_796_n 0.00155215f $X=4.42 $Y=1.105
+ $X2=0 $Y2=0
cc_509 N_A_339_112#_M1007_g N_A_959_83#_c_796_n 0.0399147f $X=4.335 $Y=0.755
+ $X2=0 $Y2=0
cc_510 N_A_339_112#_c_625_n N_A_959_83#_c_797_n 0.0864964f $X=9.3 $Y=1.59
+ $X2=17.52 $Y2=0
cc_511 N_A_339_112#_c_700_p N_A_959_83#_c_797_n 0.00952671f $X=4.42 $Y=1.24
+ $X2=17.52 $Y2=0
cc_512 N_A_339_112#_c_677_n N_A_959_83#_c_797_n 6.00174e-19 $X=4.42 $Y=1.105
+ $X2=17.52 $Y2=0
cc_513 N_A_339_112#_M1007_g N_A_959_83#_c_797_n 7.15069e-19 $X=4.335 $Y=0.755
+ $X2=17.52 $Y2=0
cc_514 N_A_339_112#_c_616_n N_A_959_83#_c_801_n 0.0399147f $X=3.85 $Y=2.195
+ $X2=0 $Y2=0
cc_515 N_A_339_112#_c_625_n N_A_959_83#_c_801_n 0.0246987f $X=9.3 $Y=1.59 $X2=0
+ $Y2=0
cc_516 N_A_339_112#_c_700_p N_A_959_83#_c_801_n 0.00235183f $X=4.42 $Y=1.24
+ $X2=0 $Y2=0
cc_517 N_A_339_112#_c_616_n N_A_959_83#_c_802_n 0.0110515f $X=3.85 $Y=2.195
+ $X2=0 $Y2=0
cc_518 N_A_339_112#_c_625_n N_A_959_83#_c_802_n 0.0152482f $X=9.3 $Y=1.59 $X2=0
+ $Y2=0
cc_519 N_A_339_112#_c_625_n N_A_761_109#_M1025_g 0.0414448f $X=9.3 $Y=1.59 $X2=0
+ $Y2=0
cc_520 N_A_339_112#_c_625_n N_A_761_109#_M1029_g 0.0316742f $X=9.3 $Y=1.59
+ $X2=17.52 $Y2=0
cc_521 N_A_339_112#_c_616_n N_A_761_109#_c_879_n 0.0156608f $X=3.85 $Y=2.195
+ $X2=0 $Y2=0
cc_522 N_A_339_112#_c_711_p N_A_761_109#_c_879_n 0.0123662f $X=4.585 $Y=1.59
+ $X2=0 $Y2=0
cc_523 N_A_339_112#_c_700_p N_A_761_109#_c_879_n 0.0285319f $X=4.42 $Y=1.24
+ $X2=0 $Y2=0
cc_524 N_A_339_112#_c_677_n N_A_761_109#_c_879_n 0.00946202f $X=4.42 $Y=1.105
+ $X2=0 $Y2=0
cc_525 N_A_339_112#_M1007_g N_A_761_109#_c_879_n 0.00457816f $X=4.335 $Y=0.755
+ $X2=0 $Y2=0
cc_526 N_A_339_112#_c_616_n N_A_761_109#_c_880_n 0.0276042f $X=3.85 $Y=2.195
+ $X2=0 $Y2=0
cc_527 N_A_339_112#_c_625_n N_A_761_109#_c_880_n 0.0284956f $X=9.3 $Y=1.59 $X2=0
+ $Y2=0
cc_528 N_A_339_112#_c_711_p N_A_761_109#_c_880_n 0.0237237f $X=4.585 $Y=1.59
+ $X2=0 $Y2=0
cc_529 N_A_339_112#_c_616_n N_A_761_109#_c_881_n 0.00976143f $X=3.85 $Y=2.195
+ $X2=0 $Y2=0
cc_530 N_A_339_112#_c_616_n N_A_761_109#_c_893_n 0.00414834f $X=3.85 $Y=2.195
+ $X2=0 $Y2=0
cc_531 N_A_339_112#_c_625_n N_A_761_109#_c_882_n 0.174574f $X=9.3 $Y=1.59 $X2=0
+ $Y2=0
cc_532 N_A_339_112#_c_625_n N_A_761_109#_c_883_n 0.00279601f $X=9.3 $Y=1.59
+ $X2=0 $Y2=0
cc_533 N_A_339_112#_c_625_n N_A_761_109#_c_946_n 0.0234399f $X=9.3 $Y=1.59 $X2=0
+ $Y2=0
cc_534 N_A_339_112#_c_621_n N_A_761_109#_c_924_n 0.0198719f $X=4.29 $Y=0.35
+ $X2=0 $Y2=0
cc_535 N_A_339_112#_c_677_n N_A_761_109#_c_924_n 0.0210746f $X=4.42 $Y=1.105
+ $X2=0 $Y2=0
cc_536 N_A_339_112#_M1007_g N_A_761_109#_c_924_n 0.00627368f $X=4.335 $Y=0.755
+ $X2=0 $Y2=0
cc_537 N_A_339_112#_M1012_g N_A_761_109#_c_895_n 0.0102472f $X=3.85 $Y=2.925
+ $X2=0 $Y2=0
cc_538 N_A_339_112#_c_625_n N_A_761_109#_c_884_n 0.0132851f $X=9.3 $Y=1.59 $X2=0
+ $Y2=0
cc_539 N_A_339_112#_c_625_n N_A_761_109#_c_885_n 0.0206002f $X=9.3 $Y=1.59 $X2=0
+ $Y2=0
cc_540 N_A_339_112#_c_626_n N_A_761_109#_c_885_n 5.16297e-19 $X=9.385 $Y=2.305
+ $X2=0 $Y2=0
cc_541 N_A_339_112#_c_625_n N_SET_B_c_1014_n 0.0334358f $X=9.3 $Y=1.59 $X2=0
+ $Y2=0
cc_542 N_A_339_112#_M1010_g N_SET_B_c_1017_n 0.0159643f $X=10.32 $Y=1.14 $X2=0
+ $Y2=0
cc_543 N_A_339_112#_c_625_n N_SET_B_c_1017_n 0.169797f $X=9.3 $Y=1.59 $X2=0
+ $Y2=0
cc_544 N_A_339_112#_M1010_g N_SET_B_c_1036_n 0.0167094f $X=10.32 $Y=1.14 $X2=0
+ $Y2=0
cc_545 N_A_339_112#_M1010_g N_SET_B_c_1018_n 0.016065f $X=10.32 $Y=1.14 $X2=0
+ $Y2=0
cc_546 N_A_339_112#_M1010_g N_SET_B_c_1042_n 0.0065245f $X=10.32 $Y=1.14 $X2=0
+ $Y2=0
cc_547 N_A_339_112#_M1010_g N_SET_B_c_1019_n 0.00493001f $X=10.32 $Y=1.14 $X2=0
+ $Y2=0
cc_548 N_A_339_112#_M1010_g N_SET_B_c_1020_n 0.0017297f $X=10.32 $Y=1.14 $X2=0
+ $Y2=0
cc_549 N_A_339_112#_M1021_g N_A_2156_417#_M1011_g 0.0118851f $X=10.015 $Y=2.925
+ $X2=0 $Y2=0
cc_550 N_A_339_112#_M1010_g N_A_2156_417#_c_1127_n 0.0183088f $X=10.32 $Y=1.14
+ $X2=0 $Y2=0
cc_551 N_A_339_112#_c_633_n N_A_2156_417#_c_1131_n 0.0354412f $X=10.32 $Y=2.335
+ $X2=0 $Y2=0
cc_552 N_A_339_112#_M1021_g N_A_1874_543#_c_1247_n 0.0170954f $X=10.015 $Y=2.925
+ $X2=0 $Y2=0
cc_553 N_A_339_112#_c_638_n N_A_1874_543#_c_1247_n 0.0101295f $X=9.47 $Y=2.39
+ $X2=0 $Y2=0
cc_554 N_A_339_112#_c_630_n N_A_1874_543#_c_1247_n 0.0153283f $X=9.855 $Y=2.43
+ $X2=0 $Y2=0
cc_555 N_A_339_112#_M1010_g N_A_1874_543#_c_1232_n 0.00897765f $X=10.32 $Y=1.14
+ $X2=0 $Y2=0
cc_556 N_A_339_112#_c_625_n N_A_1874_543#_c_1232_n 0.0136587f $X=9.3 $Y=1.59
+ $X2=0 $Y2=0
cc_557 N_A_339_112#_c_626_n N_A_1874_543#_c_1232_n 0.0207149f $X=9.385 $Y=2.305
+ $X2=0 $Y2=0
cc_558 N_A_339_112#_M1021_g N_A_1874_543#_c_1248_n 0.0155348f $X=10.015 $Y=2.925
+ $X2=0 $Y2=0
cc_559 N_A_339_112#_M1010_g N_A_1874_543#_c_1233_n 0.0166551f $X=10.32 $Y=1.14
+ $X2=0 $Y2=0
cc_560 N_A_339_112#_c_678_n N_A_1874_543#_c_1233_n 0.0136453f $X=10.02 $Y=2.39
+ $X2=0 $Y2=0
cc_561 N_A_339_112#_c_633_n N_A_1874_543#_c_1233_n 0.0142894f $X=10.32 $Y=2.335
+ $X2=0 $Y2=0
cc_562 N_A_339_112#_c_626_n N_A_1874_543#_c_1234_n 0.013786f $X=9.385 $Y=2.305
+ $X2=0 $Y2=0
cc_563 N_A_339_112#_c_630_n N_A_1874_543#_c_1234_n 0.0249918f $X=9.855 $Y=2.43
+ $X2=0 $Y2=0
cc_564 N_A_339_112#_c_633_n N_A_1874_543#_c_1234_n 0.00930087f $X=10.32 $Y=2.335
+ $X2=0 $Y2=0
cc_565 N_A_339_112#_c_678_n N_A_1874_543#_c_1278_n 0.00134959f $X=10.02 $Y=2.39
+ $X2=0 $Y2=0
cc_566 N_A_339_112#_c_633_n N_A_1874_543#_c_1278_n 0.0133813f $X=10.32 $Y=2.335
+ $X2=0 $Y2=0
cc_567 N_A_339_112#_M1021_g N_A_1874_543#_c_1254_n 0.0184676f $X=10.015 $Y=2.925
+ $X2=0 $Y2=0
cc_568 N_A_339_112#_c_678_n N_A_1874_543#_c_1254_n 0.00401203f $X=10.02 $Y=2.39
+ $X2=0 $Y2=0
cc_569 N_A_339_112#_c_633_n N_A_1874_543#_c_1254_n 0.00888017f $X=10.32 $Y=2.335
+ $X2=0 $Y2=0
cc_570 N_A_339_112#_c_678_n N_A_1874_543#_c_1283_n 0.0136541f $X=10.02 $Y=2.39
+ $X2=0 $Y2=0
cc_571 N_A_339_112#_c_633_n N_A_1874_543#_c_1283_n 0.00525246f $X=10.32 $Y=2.335
+ $X2=0 $Y2=0
cc_572 N_A_339_112#_c_633_n N_A_1874_543#_c_1238_n 0.00424666f $X=10.32 $Y=2.335
+ $X2=0 $Y2=0
cc_573 N_A_339_112#_M1021_g N_VPWR_c_1451_n 0.0156697f $X=10.015 $Y=2.925 $X2=0
+ $Y2=0
cc_574 N_A_339_112#_c_619_n N_VPWR_c_1451_n 0.0116583f $X=1.855 $Y=2.785 $X2=0
+ $Y2=0
cc_575 N_A_339_112#_c_616_n N_A_605_109#_c_1543_n 7.09853e-19 $X=3.85 $Y=2.195
+ $X2=0 $Y2=0
cc_576 N_A_339_112#_M1012_g N_A_605_109#_c_1543_n 0.00266015f $X=3.85 $Y=2.925
+ $X2=0 $Y2=0
cc_577 N_A_339_112#_c_620_n N_A_605_109#_c_1543_n 0.00733277f $X=2.65 $Y=1.25
+ $X2=0 $Y2=0
cc_578 N_A_339_112#_c_663_n N_A_605_109#_c_1543_n 0.00618285f $X=2.735 $Y=1.165
+ $X2=0 $Y2=0
cc_579 N_A_339_112#_c_663_n N_A_605_109#_c_1544_n 0.0268011f $X=2.735 $Y=1.165
+ $X2=0.24 $Y2=0
cc_580 N_A_339_112#_c_621_n N_A_605_109#_c_1544_n 0.0226433f $X=4.29 $Y=0.35
+ $X2=0.24 $Y2=0
cc_581 N_A_339_112#_M1012_g N_A_605_109#_c_1546_n 8.59971e-19 $X=3.85 $Y=2.925
+ $X2=17.52 $Y2=0
cc_582 N_A_339_112#_c_618_n N_VGND_c_1619_n 0.00109122f $X=1.885 $Y=1.165 $X2=0
+ $Y2=0
cc_583 N_A_339_112#_c_627_n N_VGND_c_1619_n 0.0336784f $X=1.835 $Y=0.77 $X2=0
+ $Y2=0
cc_584 N_A_339_112#_c_620_n N_VGND_c_1621_n 0.0193283f $X=2.65 $Y=1.25 $X2=0
+ $Y2=0
cc_585 N_A_339_112#_c_663_n N_VGND_c_1621_n 0.0231783f $X=2.735 $Y=1.165 $X2=0
+ $Y2=0
cc_586 N_A_339_112#_c_623_n N_VGND_c_1621_n 0.00474345f $X=2.82 $Y=0.35 $X2=0
+ $Y2=0
cc_587 N_A_339_112#_c_627_n N_VGND_c_1621_n 0.0292464f $X=1.835 $Y=0.77 $X2=0
+ $Y2=0
cc_588 N_A_339_112#_c_621_n N_VGND_c_1623_n 0.00452123f $X=4.29 $Y=0.35 $X2=0
+ $Y2=0
cc_589 N_A_339_112#_c_625_n N_VGND_c_1623_n 0.00768125f $X=9.3 $Y=1.59 $X2=0
+ $Y2=0
cc_590 N_A_339_112#_c_677_n N_VGND_c_1623_n 0.0318399f $X=4.42 $Y=1.105 $X2=0
+ $Y2=0
cc_591 N_A_339_112#_M1007_g N_VGND_c_1623_n 0.00364101f $X=4.335 $Y=0.755 $X2=0
+ $Y2=0
cc_592 N_A_339_112#_c_625_n N_VGND_c_1625_n 0.00633648f $X=9.3 $Y=1.59 $X2=0
+ $Y2=0
cc_593 N_A_339_112#_M1010_g N_VGND_c_1633_n 0.0173305f $X=10.32 $Y=1.14 $X2=0
+ $Y2=0
cc_594 N_A_339_112#_c_620_n N_VGND_c_1633_n 0.0140541f $X=2.65 $Y=1.25 $X2=0
+ $Y2=0
cc_595 N_A_339_112#_c_663_n N_VGND_c_1633_n 0.0199629f $X=2.735 $Y=1.165 $X2=0
+ $Y2=0
cc_596 N_A_339_112#_c_621_n N_VGND_c_1633_n 0.0586403f $X=4.29 $Y=0.35 $X2=0
+ $Y2=0
cc_597 N_A_339_112#_c_623_n N_VGND_c_1633_n 0.007754f $X=2.82 $Y=0.35 $X2=0
+ $Y2=0
cc_598 N_A_339_112#_c_627_n N_VGND_c_1633_n 0.0284415f $X=1.835 $Y=0.77 $X2=0
+ $Y2=0
cc_599 N_A_339_112#_c_700_p N_VGND_c_1633_n 0.00498399f $X=4.42 $Y=1.24 $X2=0
+ $Y2=0
cc_600 N_A_339_112#_c_677_n N_VGND_c_1633_n 0.0200485f $X=4.42 $Y=1.105 $X2=0
+ $Y2=0
cc_601 N_A_339_112#_M1007_g N_VGND_c_1633_n 0.0121419f $X=4.335 $Y=0.755 $X2=0
+ $Y2=0
cc_602 N_A_339_112#_M1010_g N_A_1642_107#_c_1741_n 0.0143108f $X=10.32 $Y=1.14
+ $X2=0.24 $Y2=0
cc_603 N_A_339_112#_M1010_g N_A_1642_107#_c_1745_n 0.00517879f $X=10.32 $Y=1.14
+ $X2=0 $Y2=0
cc_604 N_A_339_112#_M1010_g N_A_1755_153#_c_1774_n 0.0327995f $X=10.32 $Y=1.14
+ $X2=0 $Y2=0
cc_605 N_A_339_112#_M1010_g N_A_1755_153#_c_1782_n 0.0140611f $X=10.32 $Y=1.14
+ $X2=0 $Y2=0
cc_606 N_A_339_112#_M1010_g N_A_1755_153#_c_1783_n 0.00765891f $X=10.32 $Y=1.14
+ $X2=0 $Y2=0
cc_607 N_A_959_83#_c_797_n N_A_761_109#_M1025_g 0.0111481f $X=5.82 $Y=1.205
+ $X2=0 $Y2=0
cc_608 N_A_959_83#_c_799_n N_A_761_109#_M1025_g 0.0176628f $X=5.985 $Y=0.745
+ $X2=0 $Y2=0
cc_609 N_A_959_83#_c_801_n N_A_761_109#_M1025_g 0.0123115f $X=5.34 $Y=1.325
+ $X2=0 $Y2=0
cc_610 N_A_959_83#_M1009_g N_A_761_109#_M1006_g 0.0112862f $X=5.34 $Y=2.925
+ $X2=0 $Y2=0
cc_611 N_A_959_83#_c_798_n N_A_761_109#_M1006_g 0.0196459f $X=6.775 $Y=2.29
+ $X2=0 $Y2=0
cc_612 N_A_959_83#_c_805_n N_A_761_109#_M1006_g 0.00865651f $X=5.495 $Y=2.29
+ $X2=0 $Y2=0
cc_613 N_A_959_83#_c_806_n N_A_761_109#_M1006_g 0.00645782f $X=6.86 $Y=2.925
+ $X2=0 $Y2=0
cc_614 N_A_959_83#_c_801_n N_A_761_109#_c_880_n 7.99782e-19 $X=5.34 $Y=1.325
+ $X2=0 $Y2=0
cc_615 N_A_959_83#_M1009_g N_A_761_109#_c_892_n 0.00549672f $X=5.34 $Y=2.925
+ $X2=0 $Y2=0
cc_616 N_A_959_83#_M1009_g N_A_761_109#_c_893_n 0.0101163f $X=5.34 $Y=2.925
+ $X2=0 $Y2=0
cc_617 N_A_959_83#_c_798_n N_A_761_109#_c_893_n 0.0122207f $X=6.775 $Y=2.29
+ $X2=0 $Y2=0
cc_618 N_A_959_83#_c_805_n N_A_761_109#_c_893_n 0.0219443f $X=5.495 $Y=2.29
+ $X2=0 $Y2=0
cc_619 N_A_959_83#_c_802_n N_A_761_109#_c_893_n 0.00367211f $X=5.385 $Y=2.085
+ $X2=0 $Y2=0
cc_620 N_A_959_83#_c_798_n N_A_761_109#_c_882_n 0.117131f $X=6.775 $Y=2.29 $X2=0
+ $Y2=0
cc_621 N_A_959_83#_c_805_n N_A_761_109#_c_882_n 0.0025171f $X=5.495 $Y=2.29
+ $X2=0 $Y2=0
cc_622 N_A_959_83#_c_802_n N_A_761_109#_c_882_n 0.0278397f $X=5.385 $Y=2.085
+ $X2=0 $Y2=0
cc_623 N_A_959_83#_c_798_n N_A_761_109#_c_883_n 0.0139875f $X=6.775 $Y=2.29
+ $X2=0 $Y2=0
cc_624 N_A_959_83#_c_805_n N_A_761_109#_c_883_n 0.00613239f $X=5.495 $Y=2.29
+ $X2=0 $Y2=0
cc_625 N_A_959_83#_c_802_n N_A_761_109#_c_883_n 0.0123115f $X=5.385 $Y=2.085
+ $X2=0 $Y2=0
cc_626 N_A_959_83#_M1009_g N_A_761_109#_c_895_n 2.36902e-19 $X=5.34 $Y=2.925
+ $X2=0 $Y2=0
cc_627 N_A_959_83#_c_801_n N_A_761_109#_c_884_n 6.70336e-19 $X=5.34 $Y=1.325
+ $X2=0 $Y2=0
cc_628 N_A_959_83#_c_802_n N_A_761_109#_c_884_n 0.00512555f $X=5.385 $Y=2.085
+ $X2=0 $Y2=0
cc_629 N_A_959_83#_c_798_n N_A_761_109#_c_885_n 5.32359e-19 $X=6.775 $Y=2.29
+ $X2=0 $Y2=0
cc_630 N_A_959_83#_c_806_n N_A_761_109#_c_885_n 5.62441e-19 $X=6.86 $Y=2.925
+ $X2=0 $Y2=0
cc_631 N_A_959_83#_c_799_n N_SET_B_c_1013_n 7.02088e-19 $X=5.985 $Y=0.745 $X2=0
+ $Y2=0
cc_632 N_A_959_83#_c_797_n N_SET_B_c_1014_n 7.30599e-19 $X=5.82 $Y=1.205 $X2=0
+ $Y2=0
cc_633 N_A_959_83#_c_798_n N_SET_B_c_1015_n 0.00621075f $X=6.775 $Y=2.29
+ $X2=-0.33 $Y2=-0.265
cc_634 N_A_959_83#_c_798_n N_SET_B_c_1016_n 0.00231202f $X=6.775 $Y=2.29 $X2=0
+ $Y2=0
cc_635 N_A_959_83#_c_806_n N_SET_B_c_1016_n 0.0253759f $X=6.86 $Y=2.925 $X2=0
+ $Y2=0
cc_636 N_A_959_83#_M1009_g N_VPWR_c_1436_n 0.0049218f $X=5.34 $Y=2.925 $X2=0
+ $Y2=0
cc_637 N_A_959_83#_M1009_g N_VPWR_c_1451_n 0.0028551f $X=5.34 $Y=2.925 $X2=0
+ $Y2=0
cc_638 N_A_959_83#_c_806_n N_VPWR_c_1451_n 0.0016537f $X=6.86 $Y=2.925 $X2=0
+ $Y2=0
cc_639 N_A_959_83#_c_796_n N_VGND_c_1623_n 0.0456206f $X=5.045 $Y=1.075 $X2=0
+ $Y2=0
cc_640 N_A_959_83#_c_797_n N_VGND_c_1623_n 0.0441116f $X=5.82 $Y=1.205 $X2=0
+ $Y2=0
cc_641 N_A_959_83#_c_799_n N_VGND_c_1623_n 0.0268355f $X=5.985 $Y=0.745 $X2=0
+ $Y2=0
cc_642 N_A_959_83#_c_801_n N_VGND_c_1623_n 0.00784689f $X=5.34 $Y=1.325 $X2=0
+ $Y2=0
cc_643 N_A_959_83#_c_799_n N_VGND_c_1625_n 0.00576706f $X=5.985 $Y=0.745 $X2=0
+ $Y2=0
cc_644 N_A_959_83#_c_797_n N_VGND_c_1633_n 0.0111097f $X=5.82 $Y=1.205 $X2=0
+ $Y2=0
cc_645 N_A_959_83#_c_799_n N_VGND_c_1633_n 0.032098f $X=5.985 $Y=0.745 $X2=0
+ $Y2=0
cc_646 N_A_761_109#_M1025_g N_SET_B_c_1013_n 0.0806932f $X=6.375 $Y=0.745 $X2=0
+ $Y2=0
cc_647 N_A_761_109#_M1029_g N_SET_B_c_1013_n 0.0157048f $X=7.96 $Y=0.91 $X2=0
+ $Y2=0
cc_648 N_A_761_109#_M1025_g N_SET_B_c_1014_n 0.0098594f $X=6.375 $Y=0.745 $X2=0
+ $Y2=0
cc_649 N_A_761_109#_M1029_g N_SET_B_c_1014_n 0.0594811f $X=7.96 $Y=0.91 $X2=0
+ $Y2=0
cc_650 N_A_761_109#_c_882_n N_SET_B_c_1014_n 4.76725e-19 $X=7.73 $Y=1.94 $X2=0
+ $Y2=0
cc_651 N_A_761_109#_c_883_n N_SET_B_c_1014_n 0.0297409f $X=6.31 $Y=1.94 $X2=0
+ $Y2=0
cc_652 N_A_761_109#_M1006_g N_SET_B_c_1015_n 0.0297409f $X=6.47 $Y=2.925
+ $X2=-0.33 $Y2=-0.265
cc_653 N_A_761_109#_c_882_n N_SET_B_c_1015_n 0.0424697f $X=7.73 $Y=1.94
+ $X2=-0.33 $Y2=-0.265
cc_654 N_A_761_109#_c_923_n N_SET_B_c_1015_n 0.00242501f $X=7.895 $Y=2.28
+ $X2=-0.33 $Y2=-0.265
cc_655 N_A_761_109#_c_885_n N_SET_B_c_1015_n 0.0381309f $X=8.41 $Y=2.17
+ $X2=-0.33 $Y2=-0.265
cc_656 N_A_761_109#_M1006_g N_SET_B_c_1016_n 0.0127783f $X=6.47 $Y=2.925 $X2=0
+ $Y2=0
cc_657 N_A_761_109#_M1033_g N_SET_B_c_1016_n 0.00538985f $X=8.41 $Y=3.215 $X2=0
+ $Y2=0
cc_658 N_A_761_109#_M1025_g N_SET_B_c_1017_n 8.88573e-19 $X=6.375 $Y=0.745 $X2=0
+ $Y2=0
cc_659 N_A_761_109#_M1029_g N_SET_B_c_1017_n 0.032351f $X=7.96 $Y=0.91 $X2=0
+ $Y2=0
cc_660 N_A_761_109#_M1033_g N_A_1874_543#_c_1247_n 0.00104583f $X=8.41 $Y=3.215
+ $X2=0 $Y2=0
cc_661 N_A_761_109#_M1033_g N_A_1874_543#_c_1251_n 3.82301e-19 $X=8.41 $Y=3.215
+ $X2=0 $Y2=0
cc_662 N_A_761_109#_M1006_g N_VPWR_c_1436_n 0.0138587f $X=6.47 $Y=2.925 $X2=0
+ $Y2=0
cc_663 N_A_761_109#_M1033_g N_VPWR_c_1439_n 0.0636386f $X=8.41 $Y=3.215 $X2=0
+ $Y2=0
cc_664 N_A_761_109#_c_885_n N_VPWR_c_1439_n 0.00159688f $X=8.41 $Y=2.17 $X2=0
+ $Y2=0
cc_665 N_A_761_109#_M1006_g N_VPWR_c_1451_n 0.005707f $X=6.47 $Y=2.925 $X2=0
+ $Y2=0
cc_666 N_A_761_109#_M1033_g N_VPWR_c_1451_n 0.00376027f $X=8.41 $Y=3.215 $X2=0
+ $Y2=0
cc_667 N_A_761_109#_c_892_n N_VPWR_c_1451_n 0.00429716f $X=4.98 $Y=3.09 $X2=0
+ $Y2=0
cc_668 N_A_761_109#_c_895_n N_VPWR_c_1451_n 0.00211585f $X=4.24 $Y=2.925 $X2=0
+ $Y2=0
cc_669 N_A_761_109#_c_879_n N_A_605_109#_c_1544_n 0.00549275f $X=3.99 $Y=1.855
+ $X2=0.24 $Y2=0
cc_670 N_A_761_109#_c_924_n N_A_605_109#_c_1544_n 0.0115154f $X=3.945 $Y=0.77
+ $X2=0.24 $Y2=0
cc_671 N_A_761_109#_c_892_n A_976_543# 0.00160253f $X=4.98 $Y=3.09 $X2=0 $Y2=0
cc_672 N_A_761_109#_c_893_n A_976_543# 0.00367563f $X=5.065 $Y=3.005 $X2=0 $Y2=0
cc_673 N_A_761_109#_M1025_g N_VGND_c_1623_n 0.00263805f $X=6.375 $Y=0.745 $X2=0
+ $Y2=0
cc_674 N_A_761_109#_M1025_g N_VGND_c_1625_n 0.00417633f $X=6.375 $Y=0.745 $X2=0
+ $Y2=0
cc_675 N_A_761_109#_M1029_g N_VGND_c_1625_n 0.017108f $X=7.96 $Y=0.91 $X2=0
+ $Y2=0
cc_676 N_A_761_109#_M1025_g N_VGND_c_1633_n 0.033371f $X=6.375 $Y=0.745 $X2=0
+ $Y2=0
cc_677 N_A_761_109#_M1029_g N_VGND_c_1633_n 0.0139995f $X=7.96 $Y=0.91 $X2=0
+ $Y2=0
cc_678 N_A_761_109#_c_924_n N_VGND_c_1633_n 0.0212222f $X=3.945 $Y=0.77 $X2=0
+ $Y2=0
cc_679 N_A_761_109#_M1029_g N_A_1642_107#_c_1740_n 0.0118714f $X=7.96 $Y=0.91
+ $X2=0 $Y2=0
cc_680 N_A_761_109#_M1029_g N_A_1642_107#_c_1743_n 0.00649391f $X=7.96 $Y=0.91
+ $X2=0 $Y2=0
cc_681 N_SET_B_M1004_g N_A_2156_417#_M1011_g 0.01454f $X=11.81 $Y=2.925 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_1026_n N_A_2156_417#_c_1127_n 0.0296515f $X=12.595 $Y=2.335
+ $X2=0 $Y2=0
cc_683 N_SET_B_c_1018_n N_A_2156_417#_c_1127_n 0.00500535f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_684 N_SET_B_c_1019_n N_A_2156_417#_c_1127_n 0.00433478f $X=10.8 $Y=1.975
+ $X2=0 $Y2=0
cc_685 SET_B N_A_2156_417#_c_1127_n 0.00342636f $X=12.635 $Y=1.58 $X2=0 $Y2=0
cc_686 N_SET_B_c_1023_n N_A_2156_417#_c_1127_n 0.0137361f $X=12.15 $Y=1.85 $X2=0
+ $Y2=0
cc_687 N_SET_B_M1020_g N_A_2156_417#_M1019_g 0.0984514f $X=12.595 $Y=0.745 $X2=0
+ $Y2=0
cc_688 N_SET_B_c_1023_n N_A_2156_417#_c_1130_n 0.0119157f $X=12.15 $Y=1.85
+ $X2=17.52 $Y2=0
cc_689 N_SET_B_c_1026_n N_A_2156_417#_c_1131_n 0.037059f $X=12.595 $Y=2.335
+ $X2=0 $Y2=0
cc_690 N_SET_B_c_1020_n N_A_2156_417#_c_1131_n 0.00468944f $X=10.885 $Y=2.06
+ $X2=0 $Y2=0
cc_691 N_SET_B_c_1023_n N_A_2156_417#_c_1131_n 0.0139195f $X=12.15 $Y=1.85 $X2=0
+ $Y2=0
cc_692 SET_B N_A_2156_417#_c_1132_n 0.0502636f $X=12.635 $Y=1.58 $X2=8.88 $Y2=0
cc_693 N_SET_B_M1020_g N_A_2156_417#_c_1132_n 0.0291215f $X=12.595 $Y=0.745
+ $X2=8.88 $Y2=0
cc_694 N_SET_B_c_1023_n N_A_2156_417#_c_1132_n 0.00496312f $X=12.15 $Y=1.85
+ $X2=8.88 $Y2=0
cc_695 N_SET_B_c_1026_n N_A_2156_417#_c_1139_n 0.00130613f $X=12.595 $Y=2.335
+ $X2=0 $Y2=0
cc_696 N_SET_B_M1020_g N_A_2156_417#_c_1133_n 0.00694832f $X=12.595 $Y=0.745
+ $X2=0 $Y2=0
cc_697 N_SET_B_c_1026_n N_A_2156_417#_c_1161_n 3.18668e-19 $X=12.595 $Y=2.335
+ $X2=0 $Y2=0
cc_698 SET_B N_A_2156_417#_c_1161_n 0.0193025f $X=12.635 $Y=1.58 $X2=0 $Y2=0
cc_699 N_SET_B_M1020_g N_A_2156_417#_c_1161_n 0.00135957f $X=12.595 $Y=0.745
+ $X2=0 $Y2=0
cc_700 N_SET_B_c_1023_n N_A_2156_417#_c_1161_n 0.0249746f $X=12.15 $Y=1.85 $X2=0
+ $Y2=0
cc_701 N_SET_B_c_1017_n N_A_1874_543#_M1028_d 0.00966945f $X=10.16 $Y=1.24 $X2=0
+ $Y2=0
cc_702 N_SET_B_c_1017_n N_A_1874_543#_c_1232_n 0.0254361f $X=10.16 $Y=1.24 $X2=0
+ $Y2=0
cc_703 N_SET_B_c_1036_n N_A_1874_543#_c_1232_n 0.00718574f $X=10.245 $Y=1.605
+ $X2=0 $Y2=0
cc_704 N_SET_B_c_1042_n N_A_1874_543#_c_1232_n 0.0136587f $X=10.33 $Y=1.69 $X2=0
+ $Y2=0
cc_705 N_SET_B_c_1017_n N_A_1874_543#_c_1233_n 0.0038374f $X=10.16 $Y=1.24 $X2=0
+ $Y2=0
cc_706 N_SET_B_c_1018_n N_A_1874_543#_c_1233_n 0.0145675f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_707 N_SET_B_c_1042_n N_A_1874_543#_c_1233_n 0.0122708f $X=10.33 $Y=1.69 $X2=0
+ $Y2=0
cc_708 N_SET_B_c_1019_n N_A_1874_543#_c_1233_n 0.00149394f $X=10.8 $Y=1.975
+ $X2=0 $Y2=0
cc_709 N_SET_B_c_1020_n N_A_1874_543#_c_1233_n 0.0127633f $X=10.885 $Y=2.06
+ $X2=0 $Y2=0
cc_710 N_SET_B_c_1020_n N_A_1874_543#_c_1278_n 0.0015133f $X=10.885 $Y=2.06
+ $X2=0 $Y2=0
cc_711 N_SET_B_c_1026_n N_A_1874_543#_c_1255_n 0.0299257f $X=12.595 $Y=2.335
+ $X2=0 $Y2=0
cc_712 N_SET_B_M1004_g N_A_1874_543#_c_1256_n 0.0221442f $X=11.81 $Y=2.925 $X2=0
+ $Y2=0
cc_713 N_SET_B_c_1026_n N_A_1874_543#_c_1256_n 0.0280914f $X=12.595 $Y=2.335
+ $X2=0 $Y2=0
cc_714 SET_B N_A_1874_543#_c_1256_n 0.0690533f $X=12.635 $Y=1.58 $X2=0 $Y2=0
cc_715 SET_B N_A_1874_543#_c_1235_n 0.0319827f $X=12.635 $Y=1.58 $X2=0 $Y2=0
cc_716 N_SET_B_M1020_g N_A_1874_543#_c_1235_n 0.0179674f $X=12.595 $Y=0.745
+ $X2=0 $Y2=0
cc_717 SET_B N_A_1874_543#_c_1236_n 0.014426f $X=12.635 $Y=1.58 $X2=0 $Y2=0
cc_718 N_SET_B_M1020_g N_A_1874_543#_c_1236_n 0.00437494f $X=12.595 $Y=0.745
+ $X2=0 $Y2=0
cc_719 N_SET_B_c_1026_n N_A_1874_543#_c_1238_n 0.0332227f $X=12.595 $Y=2.335
+ $X2=0 $Y2=0
cc_720 N_SET_B_c_1018_n N_A_1874_543#_c_1238_n 0.00571288f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_721 N_SET_B_c_1020_n N_A_1874_543#_c_1238_n 0.012665f $X=10.885 $Y=2.06 $X2=0
+ $Y2=0
cc_722 N_SET_B_c_1023_n N_A_1874_543#_c_1238_n 0.0690533f $X=12.15 $Y=1.85 $X2=0
+ $Y2=0
cc_723 N_SET_B_M1004_g N_VPWR_c_1442_n 0.0274222f $X=11.81 $Y=2.925 $X2=0 $Y2=0
cc_724 N_SET_B_M1004_g N_VPWR_c_1451_n 0.0124104f $X=11.81 $Y=2.925 $X2=0 $Y2=0
cc_725 N_SET_B_c_1017_n N_VGND_M1027_d 0.00222494f $X=10.16 $Y=1.24 $X2=0 $Y2=0
cc_726 N_SET_B_c_1013_n N_VGND_c_1625_n 0.0535393f $X=7.085 $Y=1.065 $X2=0 $Y2=0
cc_727 N_SET_B_c_1014_n N_VGND_c_1625_n 0.00105041f $X=7.215 $Y=1.83 $X2=0 $Y2=0
cc_728 N_SET_B_c_1017_n N_VGND_c_1625_n 0.0498214f $X=10.16 $Y=1.24 $X2=0 $Y2=0
cc_729 N_SET_B_M1020_g N_VGND_c_1627_n 0.0493878f $X=12.595 $Y=0.745 $X2=0 $Y2=0
cc_730 N_SET_B_c_1017_n N_VGND_c_1633_n 0.0245081f $X=10.16 $Y=1.24 $X2=0 $Y2=0
cc_731 N_SET_B_c_1017_n N_A_1642_107#_M1029_d 0.00282677f $X=10.16 $Y=1.24 $X2=0
+ $Y2=0
cc_732 N_SET_B_c_1017_n N_A_1642_107#_c_1740_n 0.0201798f $X=10.16 $Y=1.24 $X2=0
+ $Y2=0
cc_733 N_SET_B_c_1017_n N_A_1642_107#_c_1741_n 0.00400487f $X=10.16 $Y=1.24
+ $X2=0.24 $Y2=0
cc_734 N_SET_B_c_1017_n N_A_1755_153#_M1028_s 0.00243888f $X=10.16 $Y=1.24 $X2=0
+ $Y2=0
cc_735 N_SET_B_c_1017_n N_A_1755_153#_c_1774_n 0.0945695f $X=10.16 $Y=1.24 $X2=0
+ $Y2=0
cc_736 N_SET_B_c_1018_n N_A_1755_153#_c_1774_n 0.00421096f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_737 N_SET_B_c_1017_n N_A_1755_153#_c_1782_n 0.00724174f $X=10.16 $Y=1.24
+ $X2=0 $Y2=0
cc_738 N_SET_B_c_1018_n N_A_1755_153#_c_1775_n 0.0157109f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_739 N_SET_B_c_1023_n N_A_1755_153#_c_1775_n 0.0173967f $X=12.15 $Y=1.85 $X2=0
+ $Y2=0
cc_740 N_SET_B_c_1017_n N_A_1755_153#_c_1783_n 0.00565696f $X=10.16 $Y=1.24
+ $X2=0 $Y2=0
cc_741 N_SET_B_c_1036_n N_A_1755_153#_c_1783_n 0.00724174f $X=10.245 $Y=1.605
+ $X2=0 $Y2=0
cc_742 N_SET_B_c_1018_n N_A_1755_153#_c_1783_n 0.0106579f $X=10.715 $Y=1.69
+ $X2=0 $Y2=0
cc_743 N_SET_B_M1020_g N_A_1755_153#_c_1777_n 3.2976e-19 $X=12.595 $Y=0.745
+ $X2=0 $Y2=0
cc_744 N_A_2156_417#_c_1139_n N_A_1874_543#_M1026_g 0.020712f $X=13.525 $Y=2.425
+ $X2=0 $Y2=0
cc_745 N_A_2156_417#_c_1140_n N_A_1874_543#_M1026_g 0.0209739f $X=14.225 $Y=1.99
+ $X2=0 $Y2=0
cc_746 N_A_2156_417#_c_1141_n N_A_1874_543#_M1026_g 0.00358665f $X=13.69 $Y=1.99
+ $X2=0 $Y2=0
cc_747 N_A_2156_417#_c_1133_n N_A_1874_543#_M1003_g 0.0132329f $X=13.555
+ $Y=1.075 $X2=17.52 $Y2=0
cc_748 N_A_2156_417#_c_1134_n N_A_1874_543#_M1003_g 0.0257016f $X=14.225 $Y=1.29
+ $X2=17.52 $Y2=0
cc_749 N_A_2156_417#_c_1135_n N_A_1874_543#_M1003_g 0.00108054f $X=14.31
+ $Y=1.905 $X2=17.52 $Y2=0
cc_750 N_A_2156_417#_c_1136_n N_A_1874_543#_M1003_g 0.00336264f $X=13.555
+ $Y=1.29 $X2=17.52 $Y2=0
cc_751 N_A_2156_417#_c_1140_n N_A_1874_543#_M1018_g 0.00246575f $X=14.225
+ $Y=1.99 $X2=0 $Y2=0
cc_752 N_A_2156_417#_c_1134_n N_A_1874_543#_M1016_g 0.002534f $X=14.225 $Y=1.29
+ $X2=0 $Y2=0
cc_753 N_A_2156_417#_c_1135_n N_A_1874_543#_M1016_g 4.78632e-19 $X=14.31
+ $Y=1.905 $X2=0 $Y2=0
cc_754 N_A_2156_417#_c_1140_n N_A_1874_543#_c_1229_n 0.0127443f $X=14.225
+ $Y=1.99 $X2=0 $Y2=0
cc_755 N_A_2156_417#_c_1141_n N_A_1874_543#_c_1229_n 5.98882e-19 $X=13.69
+ $Y=1.99 $X2=0 $Y2=0
cc_756 N_A_2156_417#_c_1135_n N_A_1874_543#_c_1229_n 0.0392431f $X=14.31
+ $Y=1.905 $X2=0 $Y2=0
cc_757 N_A_2156_417#_c_1136_n N_A_1874_543#_c_1229_n 9.54986e-19 $X=13.555
+ $Y=1.29 $X2=0 $Y2=0
cc_758 N_A_2156_417#_c_1131_n N_A_1874_543#_c_1278_n 0.00127092f $X=11.065
+ $Y=2.585 $X2=0 $Y2=0
cc_759 N_A_2156_417#_M1011_g N_A_1874_543#_c_1254_n 0.00390604f $X=11.03
+ $Y=2.925 $X2=0 $Y2=0
cc_760 N_A_2156_417#_c_1131_n N_A_1874_543#_c_1254_n 6.23343e-19 $X=11.065
+ $Y=2.585 $X2=0 $Y2=0
cc_761 N_A_2156_417#_c_1139_n N_A_1874_543#_c_1255_n 0.0297311f $X=13.525
+ $Y=2.425 $X2=0 $Y2=0
cc_762 N_A_2156_417#_c_1131_n N_A_1874_543#_c_1256_n 2.7579e-19 $X=11.065
+ $Y=2.585 $X2=0 $Y2=0
cc_763 N_A_2156_417#_c_1139_n N_A_1874_543#_c_1235_n 0.0189622f $X=13.525
+ $Y=2.425 $X2=0 $Y2=0
cc_764 N_A_2156_417#_c_1141_n N_A_1874_543#_c_1235_n 0.0137876f $X=13.69 $Y=1.99
+ $X2=0 $Y2=0
cc_765 N_A_2156_417#_c_1132_n N_A_1874_543#_c_1236_n 0.0137879f $X=13.39 $Y=1.29
+ $X2=0 $Y2=0
cc_766 N_A_2156_417#_c_1132_n N_A_1874_543#_c_1237_n 0.0151165f $X=13.39 $Y=1.29
+ $X2=0 $Y2=0
cc_767 N_A_2156_417#_c_1140_n N_A_1874_543#_c_1237_n 0.0229516f $X=14.225
+ $Y=1.99 $X2=0 $Y2=0
cc_768 N_A_2156_417#_c_1141_n N_A_1874_543#_c_1237_n 0.0265557f $X=13.69 $Y=1.99
+ $X2=0 $Y2=0
cc_769 N_A_2156_417#_c_1134_n N_A_1874_543#_c_1237_n 0.0210093f $X=14.225
+ $Y=1.29 $X2=0 $Y2=0
cc_770 N_A_2156_417#_c_1135_n N_A_1874_543#_c_1237_n 0.0122207f $X=14.31
+ $Y=1.905 $X2=0 $Y2=0
cc_771 N_A_2156_417#_c_1136_n N_A_1874_543#_c_1237_n 0.0259826f $X=13.555
+ $Y=1.29 $X2=0 $Y2=0
cc_772 N_A_2156_417#_c_1131_n N_A_1874_543#_c_1238_n 0.0276943f $X=11.065
+ $Y=2.585 $X2=0 $Y2=0
cc_773 N_A_2156_417#_M1011_g N_VPWR_c_1442_n 0.0541085f $X=11.03 $Y=2.925 $X2=0
+ $Y2=0
cc_774 N_A_2156_417#_c_1131_n N_VPWR_c_1442_n 0.00211209f $X=11.065 $Y=2.585
+ $X2=0 $Y2=0
cc_775 N_A_2156_417#_c_1139_n N_VPWR_c_1445_n 0.031873f $X=13.525 $Y=2.425 $X2=0
+ $Y2=0
cc_776 N_A_2156_417#_c_1140_n N_VPWR_c_1445_n 0.0386444f $X=14.225 $Y=1.99 $X2=0
+ $Y2=0
cc_777 N_A_2156_417#_c_1140_n N_Q_N_c_1581_n 0.00532565f $X=14.225 $Y=1.99 $X2=0
+ $Y2=0
cc_778 N_A_2156_417#_c_1134_n N_Q_N_c_1581_n 0.00523966f $X=14.225 $Y=1.29 $X2=0
+ $Y2=0
cc_779 N_A_2156_417#_c_1135_n N_Q_N_c_1581_n 0.0131306f $X=14.31 $Y=1.905 $X2=0
+ $Y2=0
cc_780 N_A_2156_417#_c_1134_n N_VGND_M1003_d 0.00283596f $X=14.225 $Y=1.29 $X2=0
+ $Y2=0
cc_781 N_A_2156_417#_M1019_g N_VGND_c_1627_n 0.00872065f $X=11.885 $Y=0.745
+ $X2=0 $Y2=0
cc_782 N_A_2156_417#_c_1132_n N_VGND_c_1627_n 0.05681f $X=13.39 $Y=1.29 $X2=0
+ $Y2=0
cc_783 N_A_2156_417#_c_1133_n N_VGND_c_1627_n 0.0103492f $X=13.555 $Y=1.075
+ $X2=0 $Y2=0
cc_784 N_A_2156_417#_c_1133_n N_VGND_c_1629_n 0.0151776f $X=13.555 $Y=1.075
+ $X2=0 $Y2=0
cc_785 N_A_2156_417#_c_1134_n N_VGND_c_1629_n 0.0327012f $X=14.225 $Y=1.29 $X2=0
+ $Y2=0
cc_786 N_A_2156_417#_c_1127_n N_VGND_c_1633_n 0.003897f $X=11.885 $Y=1.085 $X2=0
+ $Y2=0
cc_787 N_A_2156_417#_M1019_g N_VGND_c_1633_n 0.0189029f $X=11.885 $Y=0.745 $X2=0
+ $Y2=0
cc_788 N_A_2156_417#_c_1132_n N_VGND_c_1633_n 0.0181744f $X=13.39 $Y=1.29 $X2=0
+ $Y2=0
cc_789 N_A_2156_417#_c_1133_n N_VGND_c_1633_n 0.0177601f $X=13.555 $Y=1.075
+ $X2=0 $Y2=0
cc_790 N_A_2156_417#_c_1134_n N_VGND_c_1633_n 0.00718403f $X=14.225 $Y=1.29
+ $X2=0 $Y2=0
cc_791 N_A_2156_417#_c_1161_n N_VGND_c_1633_n 0.0102612f $X=11.805 $Y=1.305
+ $X2=0 $Y2=0
cc_792 N_A_2156_417#_M1019_g N_A_1642_107#_c_1741_n 0.00197299f $X=11.885
+ $Y=0.745 $X2=0.24 $Y2=0
cc_793 N_A_2156_417#_M1019_g N_A_1642_107#_c_1745_n 6.08683e-19 $X=11.885
+ $Y=0.745 $X2=0 $Y2=0
cc_794 N_A_2156_417#_c_1127_n N_A_1755_153#_c_1782_n 0.00156149f $X=11.885
+ $Y=1.085 $X2=0 $Y2=0
cc_795 N_A_2156_417#_c_1127_n N_A_1755_153#_c_1775_n 0.0242011f $X=11.885
+ $Y=1.085 $X2=0 $Y2=0
cc_796 N_A_2156_417#_c_1131_n N_A_1755_153#_c_1775_n 0.0014335f $X=11.065
+ $Y=2.585 $X2=0 $Y2=0
cc_797 N_A_2156_417#_c_1161_n N_A_1755_153#_c_1775_n 0.013473f $X=11.805
+ $Y=1.305 $X2=0 $Y2=0
cc_798 N_A_2156_417#_c_1127_n N_A_1755_153#_c_1776_n 0.0142338f $X=11.885
+ $Y=1.085 $X2=17.52 $Y2=0
cc_799 N_A_2156_417#_M1019_g N_A_1755_153#_c_1776_n 0.00429069f $X=11.885
+ $Y=0.745 $X2=17.52 $Y2=0
cc_800 N_A_2156_417#_c_1161_n N_A_1755_153#_c_1776_n 0.00703219f $X=11.805
+ $Y=1.305 $X2=17.52 $Y2=0
cc_801 N_A_2156_417#_c_1127_n N_A_1755_153#_c_1777_n 0.00859857f $X=11.885
+ $Y=1.085 $X2=0 $Y2=0
cc_802 N_A_2156_417#_M1019_g N_A_1755_153#_c_1777_n 0.0127971f $X=11.885
+ $Y=0.745 $X2=0 $Y2=0
cc_803 N_A_2156_417#_c_1161_n N_A_1755_153#_c_1777_n 0.00142968f $X=11.805
+ $Y=1.305 $X2=0 $Y2=0
cc_804 N_A_1874_543#_M1016_g N_A_3129_479#_c_1389_n 0.00157514f $X=14.82 $Y=0.91
+ $X2=0 $Y2=0
cc_805 N_A_1874_543#_c_1228_n N_A_3129_479#_c_1389_n 0.00951467f $X=15.93
+ $Y=1.665 $X2=0 $Y2=0
cc_806 N_A_1874_543#_M1013_g N_A_3129_479#_c_1389_n 0.0176553f $X=16.2 $Y=1.075
+ $X2=0 $Y2=0
cc_807 N_A_1874_543#_c_1231_n N_A_3129_479#_c_1389_n 0.00438153f $X=16.19
+ $Y=1.665 $X2=0 $Y2=0
cc_808 N_A_1874_543#_M1018_g N_A_3129_479#_c_1393_n 0.00297992f $X=14.81
+ $Y=2.965 $X2=0 $Y2=0
cc_809 N_A_1874_543#_c_1228_n N_A_3129_479#_c_1393_n 0.0162842f $X=15.93
+ $Y=1.665 $X2=0 $Y2=0
cc_810 N_A_1874_543#_M1024_g N_A_3129_479#_c_1393_n 0.024051f $X=16.18 $Y=2.77
+ $X2=0 $Y2=0
cc_811 N_A_1874_543#_c_1231_n N_A_3129_479#_c_1393_n 0.0348705f $X=16.19
+ $Y=1.665 $X2=0 $Y2=0
cc_812 N_A_1874_543#_c_1231_n N_A_3129_479#_c_1390_n 0.0432777f $X=16.19
+ $Y=1.665 $X2=0 $Y2=0
cc_813 N_A_1874_543#_c_1228_n N_A_3129_479#_c_1406_n 0.0078988f $X=15.93
+ $Y=1.665 $X2=0 $Y2=0
cc_814 N_A_1874_543#_c_1231_n N_A_3129_479#_c_1406_n 0.00170675f $X=16.19
+ $Y=1.665 $X2=0 $Y2=0
cc_815 N_A_1874_543#_c_1231_n N_A_3129_479#_c_1408_n 0.00335075f $X=16.19
+ $Y=1.665 $X2=8.88 $Y2=0
cc_816 N_A_1874_543#_M1024_g N_A_3129_479#_M1002_g 0.0176917f $X=16.18 $Y=2.77
+ $X2=0 $Y2=0
cc_817 N_A_1874_543#_M1013_g N_A_3129_479#_M1002_g 0.0491409f $X=16.2 $Y=1.075
+ $X2=0 $Y2=0
cc_818 N_A_1874_543#_c_1247_n N_VPWR_c_1439_n 0.0205261f $X=9.51 $Y=2.84 $X2=0
+ $Y2=0
cc_819 N_A_1874_543#_c_1251_n N_VPWR_c_1439_n 0.00188358f $X=9.675 $Y=3.67 $X2=0
+ $Y2=0
cc_820 N_A_1874_543#_c_1248_n N_VPWR_c_1442_n 0.00839908f $X=10.365 $Y=3.67
+ $X2=0 $Y2=0
cc_821 N_A_1874_543#_c_1254_n N_VPWR_c_1442_n 0.0703823f $X=10.45 $Y=3.585 $X2=0
+ $Y2=0
cc_822 N_A_1874_543#_c_1256_n N_VPWR_c_1442_n 0.0224501f $X=12.46 $Y=2.75 $X2=0
+ $Y2=0
cc_823 N_A_1874_543#_c_1238_n N_VPWR_c_1442_n 0.0715692f $X=12.035 $Y=2.75 $X2=0
+ $Y2=0
cc_824 N_A_1874_543#_M1026_g N_VPWR_c_1445_n 0.04426f $X=13.915 $Y=2.425 $X2=0
+ $Y2=0
cc_825 N_A_1874_543#_M1018_g N_VPWR_c_1445_n 0.0749039f $X=14.81 $Y=2.965 $X2=0
+ $Y2=0
cc_826 N_A_1874_543#_c_1229_n N_VPWR_c_1445_n 0.00366047f $X=15.07 $Y=1.665
+ $X2=0 $Y2=0
cc_827 N_A_1874_543#_M1024_g N_VPWR_c_1448_n 0.0779387f $X=16.18 $Y=2.77 $X2=0
+ $Y2=0
cc_828 N_A_1874_543#_c_1231_n N_VPWR_c_1448_n 0.0010557f $X=16.19 $Y=1.665 $X2=0
+ $Y2=0
cc_829 N_A_1874_543#_M1018_g N_VPWR_c_1451_n 0.0120329f $X=14.81 $Y=2.965 $X2=0
+ $Y2=0
cc_830 N_A_1874_543#_M1024_g N_VPWR_c_1451_n 0.00649418f $X=16.18 $Y=2.77 $X2=0
+ $Y2=0
cc_831 N_A_1874_543#_c_1247_n N_VPWR_c_1451_n 0.0318324f $X=9.51 $Y=2.84 $X2=0
+ $Y2=0
cc_832 N_A_1874_543#_c_1248_n N_VPWR_c_1451_n 0.0415875f $X=10.365 $Y=3.67 $X2=0
+ $Y2=0
cc_833 N_A_1874_543#_c_1251_n N_VPWR_c_1451_n 0.0119407f $X=9.675 $Y=3.67 $X2=0
+ $Y2=0
cc_834 N_A_1874_543#_c_1254_n N_VPWR_c_1451_n 0.0185161f $X=10.45 $Y=3.585 $X2=0
+ $Y2=0
cc_835 N_A_1874_543#_c_1255_n N_VPWR_c_1451_n 0.00877051f $X=13.01 $Y=2.75 $X2=0
+ $Y2=0
cc_836 N_A_1874_543#_c_1256_n N_VPWR_c_1451_n 0.0504106f $X=12.46 $Y=2.75 $X2=0
+ $Y2=0
cc_837 N_A_1874_543#_c_1254_n A_2053_543# 0.0118196f $X=10.45 $Y=3.585 $X2=0
+ $Y2=0
cc_838 N_A_1874_543#_M1018_g N_Q_N_c_1581_n 0.0489451f $X=14.81 $Y=2.965 $X2=0
+ $Y2=0
cc_839 N_A_1874_543#_M1016_g N_Q_N_c_1581_n 0.0306998f $X=14.82 $Y=0.91 $X2=0
+ $Y2=0
cc_840 N_A_1874_543#_c_1228_n N_Q_N_c_1581_n 0.0338552f $X=15.93 $Y=1.665 $X2=0
+ $Y2=0
cc_841 N_A_1874_543#_c_1229_n N_Q_N_c_1581_n 0.0169156f $X=15.07 $Y=1.665 $X2=0
+ $Y2=0
cc_842 N_A_1874_543#_M1024_g N_Q_N_c_1581_n 0.00258088f $X=16.18 $Y=2.77 $X2=0
+ $Y2=0
cc_843 N_A_1874_543#_M1013_g N_Q_N_c_1581_n 0.00398099f $X=16.2 $Y=1.075 $X2=0
+ $Y2=0
cc_844 N_A_1874_543#_c_1231_n N_Q_N_c_1581_n 0.00364019f $X=16.19 $Y=1.665 $X2=0
+ $Y2=0
cc_845 N_A_1874_543#_M1003_g N_VGND_c_1627_n 0.00325727f $X=13.945 $Y=1.075
+ $X2=0 $Y2=0
cc_846 N_A_1874_543#_M1003_g N_VGND_c_1629_n 0.0301013f $X=13.945 $Y=1.075 $X2=0
+ $Y2=0
cc_847 N_A_1874_543#_M1016_g N_VGND_c_1629_n 0.04711f $X=14.82 $Y=0.91 $X2=0
+ $Y2=0
cc_848 N_A_1874_543#_c_1229_n N_VGND_c_1629_n 0.00365804f $X=15.07 $Y=1.665
+ $X2=0 $Y2=0
cc_849 N_A_1874_543#_M1013_g N_VGND_c_1631_n 0.0464513f $X=16.2 $Y=1.075 $X2=0
+ $Y2=0
cc_850 N_A_1874_543#_M1003_g N_VGND_c_1633_n 0.00672879f $X=13.945 $Y=1.075
+ $X2=0 $Y2=0
cc_851 N_A_1874_543#_M1016_g N_VGND_c_1633_n 0.0121699f $X=14.82 $Y=0.91 $X2=0
+ $Y2=0
cc_852 N_A_1874_543#_M1013_g N_VGND_c_1633_n 0.00672879f $X=16.2 $Y=1.075 $X2=0
+ $Y2=0
cc_853 N_A_1874_543#_M1028_d N_A_1755_153#_c_1774_n 0.00610903f $X=9.56 $Y=0.765
+ $X2=0 $Y2=0
cc_854 N_A_3129_479#_c_1393_n N_VPWR_c_1448_n 0.0629871f $X=15.79 $Y=2.52 $X2=0
+ $Y2=0
cc_855 N_A_3129_479#_c_1408_n N_VPWR_c_1448_n 0.019212f $X=17.01 $Y=1.67 $X2=0
+ $Y2=0
cc_856 N_A_3129_479#_M1002_g N_VPWR_c_1448_n 0.0613135f $X=17.075 $Y=0.91 $X2=0
+ $Y2=0
cc_857 N_A_3129_479#_c_1393_n N_VPWR_c_1451_n 0.0170977f $X=15.79 $Y=2.52 $X2=0
+ $Y2=0
cc_858 N_A_3129_479#_M1002_g N_VPWR_c_1451_n 0.0145323f $X=17.075 $Y=0.91 $X2=0
+ $Y2=0
cc_859 N_A_3129_479#_c_1389_n N_Q_N_c_1581_n 0.0429608f $X=15.81 $Y=1.075 $X2=0
+ $Y2=0
cc_860 N_A_3129_479#_c_1393_n N_Q_N_c_1581_n 0.0946662f $X=15.79 $Y=2.52 $X2=0
+ $Y2=0
cc_861 N_A_3129_479#_c_1406_n N_Q_N_c_1581_n 0.0100196f $X=15.8 $Y=1.59 $X2=0
+ $Y2=0
cc_862 N_A_3129_479#_c_1408_n Q 0.0416943f $X=17.01 $Y=1.67 $X2=0 $Y2=0
cc_863 N_A_3129_479#_M1002_g Q 0.0361542f $X=17.075 $Y=0.91 $X2=0 $Y2=0
cc_864 N_A_3129_479#_M1002_g Q 0.0176721f $X=17.075 $Y=0.91 $X2=0 $Y2=0
cc_865 N_A_3129_479#_M1002_g N_Q_c_1604_n 0.0138385f $X=17.075 $Y=0.91 $X2=0
+ $Y2=0
cc_866 N_A_3129_479#_M1002_g Q 0.00506627f $X=17.075 $Y=0.91 $X2=0 $Y2=0
cc_867 N_A_3129_479#_c_1389_n N_VGND_c_1631_n 0.0365819f $X=15.81 $Y=1.075 $X2=0
+ $Y2=0
cc_868 N_A_3129_479#_c_1390_n N_VGND_c_1631_n 0.049195f $X=16.845 $Y=1.59 $X2=0
+ $Y2=0
cc_869 N_A_3129_479#_c_1408_n N_VGND_c_1631_n 0.0192002f $X=17.01 $Y=1.67 $X2=0
+ $Y2=0
cc_870 N_A_3129_479#_M1002_g N_VGND_c_1631_n 0.0500842f $X=17.075 $Y=0.91 $X2=0
+ $Y2=0
cc_871 N_A_3129_479#_c_1389_n N_VGND_c_1633_n 0.0192623f $X=15.81 $Y=1.075 $X2=0
+ $Y2=0
cc_872 N_A_3129_479#_M1002_g N_VGND_c_1633_n 0.0124139f $X=17.075 $Y=0.91 $X2=0
+ $Y2=0
cc_873 N_VPWR_c_1451_n N_A_605_109#_c_1546_n 0.00215844f $X=16.97 $Y=3.59
+ $X2=17.52 $Y2=4.07
cc_874 N_VPWR_c_1439_n A_1732_543# 0.0123114f $X=8.02 $Y=2.995 $X2=0 $Y2=3.985
cc_875 N_VPWR_c_1451_n A_1732_543# 0.00275248f $X=16.97 $Y=3.59 $X2=0 $Y2=3.985
cc_876 N_VPWR_c_1442_n A_2053_543# 0.00417521f $X=11.42 $Y=2.925 $X2=0 $Y2=3.985
cc_877 N_VPWR_c_1445_n N_Q_N_c_1581_n 0.102672f $X=14.42 $Y=2.34 $X2=8.88
+ $Y2=4.07
cc_878 N_VPWR_c_1451_n N_Q_N_c_1581_n 0.0489796f $X=16.97 $Y=3.59 $X2=8.88
+ $Y2=4.07
cc_879 N_VPWR_c_1451_n Q 0.015253f $X=16.97 $Y=3.59 $X2=0.24 $Y2=4.07
cc_880 N_VPWR_c_1448_n Q 0.0711583f $X=16.685 $Y=2.52 $X2=0 $Y2=0
cc_881 N_A_605_109#_c_1544_n N_VGND_c_1633_n 0.0246727f $X=3.165 $Y=0.77 $X2=0
+ $Y2=0
cc_882 N_Q_N_c_1581_n N_VGND_c_1629_n 0.0385345f $X=15.21 $Y=0.66 $X2=0 $Y2=0
cc_883 N_Q_N_c_1581_n N_VGND_c_1633_n 0.0370341f $X=15.21 $Y=0.66 $X2=0 $Y2=0
cc_884 N_Q_c_1604_n N_VGND_c_1631_n 0.0557295f $X=17.465 $Y=0.66 $X2=0 $Y2=0
cc_885 N_Q_c_1604_n N_VGND_c_1633_n 0.0337615f $X=17.465 $Y=0.66 $X2=0 $Y2=0
cc_886 N_VGND_c_1623_n A_917_109# 0.00471723f $X=5.485 $Y=0.48 $X2=0 $Y2=0
cc_887 N_VGND_c_1633_n A_917_109# 0.00271077f $X=16.99 $Y=0.48 $X2=0 $Y2=0
cc_888 N_VGND_c_1633_n A_1325_107# 0.00663096f $X=16.99 $Y=0.48 $X2=0 $Y2=0
cc_889 N_VGND_c_1625_n N_A_1642_107#_c_1740_n 0.0141247f $X=7.62 $Y=0.48 $X2=0
+ $Y2=0
cc_890 N_VGND_c_1633_n N_A_1642_107#_c_1740_n 0.0135661f $X=16.99 $Y=0.48 $X2=0
+ $Y2=0
cc_891 N_VGND_c_1633_n N_A_1642_107#_c_1741_n 0.0936031f $X=16.99 $Y=0.48
+ $X2=0.24 $Y2=0
cc_892 N_VGND_c_1625_n N_A_1642_107#_c_1743_n 0.00346782f $X=7.62 $Y=0.48 $X2=0
+ $Y2=0
cc_893 N_VGND_c_1633_n N_A_1642_107#_c_1743_n 0.0126019f $X=16.99 $Y=0.48 $X2=0
+ $Y2=0
cc_894 N_VGND_c_1633_n N_A_1642_107#_c_1745_n 0.0187652f $X=16.99 $Y=0.48 $X2=0
+ $Y2=0
cc_895 N_VGND_c_1633_n N_A_1755_153#_c_1774_n 0.0626285f $X=16.99 $Y=0.48 $X2=0
+ $Y2=0
cc_896 N_VGND_c_1627_n N_A_1755_153#_c_1777_n 0.0135394f $X=13.035 $Y=0.48 $X2=0
+ $Y2=0
cc_897 N_VGND_c_1633_n N_A_1755_153#_c_1777_n 0.0244072f $X=16.99 $Y=0.48 $X2=0
+ $Y2=0
cc_898 N_VGND_c_1627_n A_2427_107# 0.005615f $X=13.035 $Y=0.48 $X2=0 $Y2=0
cc_899 N_VGND_c_1633_n A_2427_107# 9.14588e-19 $X=16.99 $Y=0.48 $X2=0 $Y2=0
cc_900 N_A_1642_107#_M1010_d N_A_1755_153#_c_1774_n 0.00238654f $X=10.57
+ $Y=0.765 $X2=0 $Y2=0
cc_901 N_A_1642_107#_c_1740_n N_A_1755_153#_c_1774_n 0.0172255f $X=8.35 $Y=0.785
+ $X2=0 $Y2=0
cc_902 N_A_1642_107#_c_1741_n N_A_1755_153#_c_1774_n 0.118696f $X=10.86 $Y=0.46
+ $X2=0 $Y2=0
cc_903 N_A_1642_107#_c_1745_n N_A_1755_153#_c_1774_n 0.020138f $X=10.945 $Y=0.91
+ $X2=0 $Y2=0
cc_904 N_A_1642_107#_M1010_d N_A_1755_153#_c_1782_n 0.00387692f $X=10.57
+ $Y=0.765 $X2=0 $Y2=0
cc_905 N_A_1642_107#_c_1745_n N_A_1755_153#_c_1782_n 0.00713326f $X=10.945
+ $Y=0.91 $X2=0 $Y2=0
cc_906 N_A_1642_107#_M1010_d N_A_1755_153#_c_1775_n 0.0163933f $X=10.57 $Y=0.765
+ $X2=0 $Y2=0
cc_907 N_A_1642_107#_c_1745_n N_A_1755_153#_c_1775_n 0.0195017f $X=10.945
+ $Y=0.91 $X2=0 $Y2=0
cc_908 N_A_1642_107#_M1010_d N_A_1755_153#_c_1783_n 6.02853e-19 $X=10.57
+ $Y=0.765 $X2=0 $Y2=0
cc_909 N_A_1642_107#_c_1741_n N_A_1755_153#_c_1777_n 0.00207984f $X=10.86
+ $Y=0.46 $X2=0 $Y2=0
cc_910 N_A_1642_107#_c_1745_n N_A_1755_153#_c_1777_n 0.0404719f $X=10.945
+ $Y=0.91 $X2=0 $Y2=0
