* File: sky130_fd_sc_hvl__sdfxtp_1.pxi.spice
* Created: Wed Sep  2 09:10:32 2020
* 
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%VNB N_VNB_M1011_b VNB N_VNB_c_2_p
+ PM_SKY130_FD_SC_HVL__SDFXTP_1%VNB
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%VPB N_VPB_M1003_b VPB N_VPB_c_119_p
+ PM_SKY130_FD_SC_HVL__SDFXTP_1%VPB
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%SCE N_SCE_M1011_g N_SCE_c_261_n N_SCE_c_262_n
+ N_SCE_M1003_g N_SCE_c_265_n N_SCE_M1014_g N_SCE_c_254_n N_SCE_c_255_n SCE SCE
+ SCE N_SCE_M1015_g N_SCE_c_258_n N_SCE_c_259_n N_SCE_c_260_n
+ PM_SKY130_FD_SC_HVL__SDFXTP_1%SCE
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%D N_D_M1025_g N_D_c_326_n N_D_M1016_g
+ N_D_c_327_n D D D D D N_D_c_333_n PM_SKY130_FD_SC_HVL__SDFXTP_1%D
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%A_30_593# N_A_30_593#_M1011_s
+ N_A_30_593#_M1003_s N_A_30_593#_c_370_n N_A_30_593#_M1027_g
+ N_A_30_593#_M1006_g N_A_30_593#_c_372_n N_A_30_593#_c_374_n
+ N_A_30_593#_c_375_n N_A_30_593#_c_376_n N_A_30_593#_c_394_n
+ N_A_30_593#_c_377_n PM_SKY130_FD_SC_HVL__SDFXTP_1%A_30_593#
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%SCD N_SCD_M1018_g N_SCD_M1007_g N_SCD_c_436_n
+ SCD N_SCD_c_442_n N_SCD_c_437_n PM_SKY130_FD_SC_HVL__SDFXTP_1%SCD
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%CLK N_CLK_M1008_g N_CLK_M1009_g CLK
+ N_CLK_c_477_n N_CLK_c_478_n PM_SKY130_FD_SC_HVL__SDFXTP_1%CLK
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%A_1204_107# N_A_1204_107#_M1019_d
+ N_A_1204_107#_M1020_d N_A_1204_107#_c_525_n N_A_1204_107#_M1030_g
+ N_A_1204_107#_M1029_g N_A_1204_107#_M1023_g N_A_1204_107#_c_513_n
+ N_A_1204_107#_c_527_n N_A_1204_107#_c_514_n N_A_1204_107#_c_516_n
+ N_A_1204_107#_c_528_n N_A_1204_107#_c_531_n N_A_1204_107#_c_534_n
+ N_A_1204_107#_c_518_n N_A_1204_107#_c_546_p N_A_1204_107#_c_520_n
+ N_A_1204_107#_c_565_p N_A_1204_107#_c_577_p N_A_1204_107#_c_535_n
+ N_A_1204_107#_c_536_n N_A_1204_107#_c_521_n N_A_1204_107#_M1021_g
+ N_A_1204_107#_c_524_n PM_SKY130_FD_SC_HVL__SDFXTP_1%A_1204_107#
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%A_938_107# N_A_938_107#_M1008_d
+ N_A_938_107#_M1009_d N_A_938_107#_c_659_n N_A_938_107#_M1020_g
+ N_A_938_107#_c_660_n N_A_938_107#_M1028_g N_A_938_107#_M1024_g
+ N_A_938_107#_c_679_n N_A_938_107#_c_662_n N_A_938_107#_c_663_n
+ N_A_938_107#_c_664_n N_A_938_107#_c_682_n N_A_938_107#_c_683_n
+ N_A_938_107#_c_706_n N_A_938_107#_c_748_p N_A_938_107#_c_764_p
+ N_A_938_107#_c_684_n N_A_938_107#_c_686_n N_A_938_107#_c_725_n
+ N_A_938_107#_c_688_n N_A_938_107#_c_665_n N_A_938_107#_c_666_n
+ N_A_938_107#_c_827_p N_A_938_107#_c_744_p N_A_938_107#_c_692_n
+ N_A_938_107#_c_731_n N_A_938_107#_c_695_n N_A_938_107#_M1019_g
+ N_A_938_107#_M1031_g N_A_938_107#_M1000_g N_A_938_107#_c_672_n
+ PM_SKY130_FD_SC_HVL__SDFXTP_1%A_938_107#
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%A_1688_81# N_A_1688_81#_M1013_d
+ N_A_1688_81#_M1017_d N_A_1688_81#_M1022_g N_A_1688_81#_M1026_g
+ N_A_1688_81#_c_851_n N_A_1688_81#_c_853_n N_A_1688_81#_c_860_n
+ N_A_1688_81#_c_854_n N_A_1688_81#_c_861_n N_A_1688_81#_c_856_n
+ N_A_1688_81#_c_879_n N_A_1688_81#_c_881_n N_A_1688_81#_c_894_n
+ N_A_1688_81#_c_857_n N_A_1688_81#_c_863_n N_A_1688_81#_c_864_n
+ N_A_1688_81#_c_865_n N_A_1688_81#_c_858_n
+ PM_SKY130_FD_SC_HVL__SDFXTP_1%A_1688_81#
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%A_1490_107# N_A_1490_107#_M1028_d
+ N_A_1490_107#_M1030_d N_A_1490_107#_c_937_n N_A_1490_107#_c_942_n
+ N_A_1490_107#_c_943_n N_A_1490_107#_c_938_n N_A_1490_107#_c_939_n
+ N_A_1490_107#_c_961_n N_A_1490_107#_c_944_n N_A_1490_107#_M1013_g
+ N_A_1490_107#_M1017_g PM_SKY130_FD_SC_HVL__SDFXTP_1%A_1490_107#
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%A_2352_81# N_A_2352_81#_M1002_d
+ N_A_2352_81#_M1005_d N_A_2352_81#_M1001_g N_A_2352_81#_M1004_g
+ N_A_2352_81#_M1012_g N_A_2352_81#_M1010_g N_A_2352_81#_c_1016_n
+ N_A_2352_81#_c_1017_n N_A_2352_81#_c_1018_n N_A_2352_81#_c_1019_n
+ N_A_2352_81#_c_1021_n N_A_2352_81#_c_1029_n N_A_2352_81#_c_1044_p
+ N_A_2352_81#_c_1022_n PM_SKY130_FD_SC_HVL__SDFXTP_1%A_2352_81#
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%A_2123_543# N_A_2123_543#_M1029_d
+ N_A_2123_543#_M1031_d N_A_2123_543#_M1002_g N_A_2123_543#_M1005_g
+ N_A_2123_543#_c_1107_n N_A_2123_543#_c_1108_n N_A_2123_543#_c_1110_n
+ N_A_2123_543#_c_1112_n N_A_2123_543#_c_1119_n N_A_2123_543#_c_1120_n
+ N_A_2123_543#_c_1170_n N_A_2123_543#_c_1113_n N_A_2123_543#_c_1122_n
+ PM_SKY130_FD_SC_HVL__SDFXTP_1%A_2123_543#
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%VPWR N_VPWR_M1003_d N_VPWR_M1007_d
+ N_VPWR_M1020_s N_VPWR_M1026_d N_VPWR_M1004_d N_VPWR_M1010_d VPWR
+ N_VPWR_c_1201_n N_VPWR_c_1204_n N_VPWR_c_1207_n N_VPWR_c_1210_n
+ N_VPWR_c_1213_n N_VPWR_c_1216_n N_VPWR_c_1219_n
+ PM_SKY130_FD_SC_HVL__SDFXTP_1%VPWR
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%A_484_107# N_A_484_107#_M1027_d
+ N_A_484_107#_M1028_s N_A_484_107#_M1016_d N_A_484_107#_M1030_s
+ N_A_484_107#_c_1295_n N_A_484_107#_c_1303_n N_A_484_107#_c_1296_n
+ N_A_484_107#_c_1304_n N_A_484_107#_c_1297_n N_A_484_107#_c_1298_n
+ N_A_484_107#_c_1299_n N_A_484_107#_c_1306_n N_A_484_107#_c_1301_n
+ N_A_484_107#_c_1302_n N_A_484_107#_c_1309_n N_A_484_107#_c_1310_n
+ N_A_484_107#_c_1311_n PM_SKY130_FD_SC_HVL__SDFXTP_1%A_484_107#
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%Q N_Q_M1012_s N_Q_M1010_s N_Q_c_1392_n
+ N_Q_c_1396_n N_Q_c_1394_n N_Q_c_1399_n N_Q_c_1400_n Q Q
+ PM_SKY130_FD_SC_HVL__SDFXTP_1%Q
x_PM_SKY130_FD_SC_HVL__SDFXTP_1%VGND N_VGND_M1011_d N_VGND_M1018_d
+ N_VGND_M1019_s N_VGND_M1022_d N_VGND_M1001_d N_VGND_M1012_d VGND
+ N_VGND_c_1430_n N_VGND_c_1432_n N_VGND_c_1434_n N_VGND_c_1436_n
+ N_VGND_c_1438_n N_VGND_c_1440_n N_VGND_c_1442_n
+ PM_SKY130_FD_SC_HVL__SDFXTP_1%VGND
cc_1 N_VNB_M1011_b N_SCE_M1011_g 0.081977f $X=-0.33 $Y=-0.265 $X2=0.68 $Y2=0.745
cc_2 N_VNB_c_2_p N_SCE_M1011_g 0.00221094f $X=0.24 $Y=0 $X2=0.68 $Y2=0.745
cc_3 N_VNB_M1011_b N_SCE_c_254_n 0.0103657f $X=-0.33 $Y=-0.265 $X2=2.72 $Y2=1.94
cc_4 N_VNB_M1011_b N_SCE_c_255_n 0.00141347f $X=-0.33 $Y=-0.265 $X2=2.885
+ $Y2=1.25
cc_5 N_VNB_M1011_b N_SCE_M1015_g 0.113176f $X=-0.33 $Y=-0.265 $X2=2.95 $Y2=0.745
cc_6 N_VNB_c_2_p N_SCE_M1015_g 0.0023273f $X=0.24 $Y=0 $X2=2.95 $Y2=0.745
cc_7 N_VNB_M1011_b N_SCE_c_258_n 0.0491807f $X=-0.33 $Y=-0.265 $X2=0.77
+ $Y2=1.565
cc_8 N_VNB_M1011_b N_SCE_c_259_n 0.00261716f $X=-0.33 $Y=-0.265 $X2=1.505
+ $Y2=1.735
cc_9 N_VNB_M1011_b N_SCE_c_260_n 0.0042798f $X=-0.33 $Y=-0.265 $X2=1.795
+ $Y2=1.735
cc_10 N_VNB_M1011_b N_D_M1025_g 0.0584448f $X=-0.33 $Y=-0.265 $X2=0.68 $Y2=0.745
cc_11 N_VNB_M1011_b N_D_c_326_n 0.0200735f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=2.355
cc_12 N_VNB_M1011_b N_D_c_327_n 0.024524f $X=-0.33 $Y=-0.265 $X2=1.465 $Y2=3.175
cc_13 N_VNB_M1011_b N_A_30_593#_c_370_n 0.0481768f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.855
cc_14 N_VNB_c_2_p N_A_30_593#_c_370_n 0.0023273f $X=0.24 $Y=0 $X2=0.685
+ $Y2=2.855
cc_15 N_VNB_M1011_b N_A_30_593#_c_372_n 0.0310029f $X=-0.33 $Y=-0.265 $X2=2.72
+ $Y2=1.94
cc_16 N_VNB_c_2_p N_A_30_593#_c_372_n 7.98897e-19 $X=0.24 $Y=0 $X2=2.72 $Y2=1.94
cc_17 N_VNB_M1011_b N_A_30_593#_c_374_n 0.0317946f $X=-0.33 $Y=-0.265 $X2=2.885
+ $Y2=1.25
cc_18 N_VNB_M1011_b N_A_30_593#_c_375_n 0.00996101f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_19 N_VNB_M1011_b N_A_30_593#_c_376_n 0.00974601f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_20 N_VNB_M1011_b N_A_30_593#_c_377_n 0.0806777f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_21 N_VNB_M1011_b N_SCD_M1018_g 0.042028f $X=-0.33 $Y=-0.265 $X2=0.68
+ $Y2=0.745
cc_22 N_VNB_c_2_p N_SCD_M1018_g 7.95938e-19 $X=0.24 $Y=0 $X2=0.68 $Y2=0.745
cc_23 N_VNB_M1011_b N_SCD_c_436_n 0.0481725f $X=-0.33 $Y=-0.265 $X2=1.465
+ $Y2=3.175
cc_24 N_VNB_M1011_b N_SCD_c_437_n 0.0277447f $X=-0.33 $Y=-0.265 $X2=2.885
+ $Y2=1.855
cc_25 N_VNB_M1011_b N_CLK_M1009_g 0.0121236f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=2.355
cc_26 N_VNB_M1011_b N_CLK_c_477_n 0.0943646f $X=-0.33 $Y=-0.265 $X2=1.465
+ $Y2=3.175
cc_27 N_VNB_M1011_b N_CLK_c_478_n 0.0456844f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.605
cc_28 N_VNB_c_2_p N_CLK_c_478_n 9.58849e-19 $X=0.24 $Y=0 $X2=0.685 $Y2=2.605
cc_29 N_VNB_M1011_b N_A_1204_107#_M1029_g 0.0837573f $X=-0.33 $Y=-0.265
+ $X2=1.465 $Y2=3.175
cc_30 N_VNB_c_2_p N_A_1204_107#_M1029_g 0.0023273f $X=0.24 $Y=0 $X2=1.465
+ $Y2=3.175
cc_31 N_VNB_M1011_b N_A_1204_107#_c_513_n 0.0129166f $X=-0.33 $Y=-0.265
+ $X2=2.885 $Y2=1.25
cc_32 N_VNB_M1011_b N_A_1204_107#_c_514_n 0.0596738f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_33 N_VNB_c_2_p N_A_1204_107#_c_514_n 0.0025323f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_34 N_VNB_M1011_b N_A_1204_107#_c_516_n 0.0257487f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_35 N_VNB_c_2_p N_A_1204_107#_c_516_n 0.00109373f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_36 N_VNB_M1011_b N_A_1204_107#_c_518_n 0.0699818f $X=-0.33 $Y=-0.265
+ $X2=0.692 $Y2=1.565
cc_37 N_VNB_c_2_p N_A_1204_107#_c_518_n 0.00324159f $X=0.24 $Y=0 $X2=0.692
+ $Y2=1.565
cc_38 N_VNB_M1011_b N_A_1204_107#_c_520_n 0.0175371f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_39 N_VNB_M1011_b N_A_1204_107#_c_521_n 0.0121104f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_c_2_p N_A_1204_107#_c_521_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_41 N_VNB_M1011_b N_A_1204_107#_M1021_g 0.073611f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_42 N_VNB_M1011_b N_A_1204_107#_c_524_n 0.0940497f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_M1011_b N_A_938_107#_c_659_n 0.0717999f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.855
cc_44 N_VNB_M1011_b N_A_938_107#_c_660_n 0.0811053f $X=-0.33 $Y=-0.265 $X2=1.465
+ $Y2=3.175
cc_45 N_VNB_M1011_b N_A_938_107#_M1028_g 0.0601813f $X=-0.33 $Y=-0.265 $X2=1.465
+ $Y2=2.855
cc_46 N_VNB_M1011_b N_A_938_107#_c_662_n 0.0049209f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_47 N_VNB_M1011_b N_A_938_107#_c_663_n 0.0151365f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_M1011_b N_A_938_107#_c_664_n 0.00482705f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_49 N_VNB_M1011_b N_A_938_107#_c_665_n 0.00293898f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_M1011_b N_A_938_107#_c_666_n 0.019659f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_51 N_VNB_c_2_p N_A_938_107#_c_666_n 8.65353e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_52 N_VNB_M1011_b N_A_938_107#_M1019_g 0.0723749f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_53 N_VNB_c_2_p N_A_938_107#_M1019_g 8.8903e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_54 N_VNB_M1011_b N_A_938_107#_M1000_g 0.0839299f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_55 N_VNB_c_2_p N_A_938_107#_M1000_g 0.0023273f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_56 N_VNB_M1011_b N_A_938_107#_c_672_n 0.0790785f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_57 N_VNB_M1011_b N_A_1688_81#_c_851_n 0.0424185f $X=-0.33 $Y=-0.265 $X2=2.72
+ $Y2=1.94
cc_58 N_VNB_c_2_p N_A_1688_81#_c_851_n 0.00112176f $X=0.24 $Y=0 $X2=2.72
+ $Y2=1.94
cc_59 N_VNB_M1011_b N_A_1688_81#_c_853_n 0.0496677f $X=-0.33 $Y=-0.265 $X2=1.795
+ $Y2=1.94
cc_60 N_VNB_M1011_b N_A_1688_81#_c_854_n 0.0119173f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_61 N_VNB_c_2_p N_A_1688_81#_c_854_n 8.20147e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_62 N_VNB_M1011_b N_A_1688_81#_c_856_n 5.9799e-19 $X=-0.33 $Y=-0.265 $X2=2.95
+ $Y2=0.745
cc_63 N_VNB_M1011_b N_A_1688_81#_c_857_n 0.00246408f $X=-0.33 $Y=-0.265 $X2=0.77
+ $Y2=1.565
cc_64 N_VNB_M1011_b N_A_1688_81#_c_858_n 0.0280007f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_65 N_VNB_M1011_b N_A_1490_107#_c_937_n 0.0053143f $X=-0.33 $Y=-0.265
+ $X2=0.685 $Y2=3.175
cc_66 N_VNB_M1011_b N_A_1490_107#_c_938_n 0.0200187f $X=-0.33 $Y=-0.265
+ $X2=1.795 $Y2=1.94
cc_67 N_VNB_M1011_b N_A_1490_107#_c_939_n 6.35731e-19 $X=-0.33 $Y=-0.265
+ $X2=2.885 $Y2=1.25
cc_68 N_VNB_M1011_b N_A_1490_107#_M1013_g 0.086529f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_69 N_VNB_c_2_p N_A_1490_107#_M1013_g 9.58849e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_70 N_VNB_M1011_b N_A_2352_81#_M1001_g 0.0742874f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=3.175
cc_71 N_VNB_c_2_p N_A_2352_81#_M1001_g 0.00102867f $X=0.24 $Y=0 $X2=0.685
+ $Y2=3.175
cc_72 N_VNB_M1011_b N_A_2352_81#_M1012_g 0.0528302f $X=-0.33 $Y=-0.265 $X2=1.795
+ $Y2=1.94
cc_73 N_VNB_c_2_p N_A_2352_81#_M1012_g 9.80755e-19 $X=0.24 $Y=0 $X2=1.795
+ $Y2=1.94
cc_74 N_VNB_M1011_b N_A_2352_81#_c_1016_n 0.0505088f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=1.58
cc_75 N_VNB_M1011_b N_A_2352_81#_c_1017_n 0.0330269f $X=-0.33 $Y=-0.265
+ $X2=1.115 $Y2=1.58
cc_76 N_VNB_M1011_b N_A_2352_81#_c_1018_n 0.0118519f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_77 N_VNB_M1011_b N_A_2352_81#_c_1019_n 0.0203594f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_78 N_VNB_c_2_p N_A_2352_81#_c_1019_n 7.98897e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_79 N_VNB_M1011_b N_A_2352_81#_c_1021_n 2.63736e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_80 N_VNB_M1011_b N_A_2352_81#_c_1022_n 0.0427844f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_81 N_VNB_M1011_b N_A_2123_543#_M1002_g 0.0833452f $X=-0.33 $Y=-0.265
+ $X2=0.685 $Y2=3.175
cc_82 N_VNB_c_2_p N_A_2123_543#_M1002_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.685
+ $Y2=3.175
cc_83 N_VNB_M1011_b N_A_2123_543#_c_1107_n 0.00662538f $X=-0.33 $Y=-0.265
+ $X2=2.885 $Y2=1.855
cc_84 N_VNB_M1011_b N_A_2123_543#_c_1108_n 0.0195854f $X=-0.33 $Y=-0.265
+ $X2=2.885 $Y2=1.25
cc_85 N_VNB_c_2_p N_A_2123_543#_c_1108_n 0.00251265f $X=0.24 $Y=0 $X2=2.885
+ $Y2=1.25
cc_86 N_VNB_M1011_b N_A_2123_543#_c_1110_n 0.00908061f $X=-0.33 $Y=-0.265
+ $X2=2.885 $Y2=1.25
cc_87 N_VNB_c_2_p N_A_2123_543#_c_1110_n 6.39361e-19 $X=0.24 $Y=0 $X2=2.885
+ $Y2=1.25
cc_88 N_VNB_M1011_b N_A_2123_543#_c_1112_n 0.00649691f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_89 N_VNB_M1011_b N_A_2123_543#_c_1113_n 0.00669549f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_90 N_VNB_M1011_b N_A_484_107#_c_1295_n 0.00636292f $X=-0.33 $Y=-0.265
+ $X2=0.685 $Y2=2.605
cc_91 N_VNB_M1011_b N_A_484_107#_c_1296_n 0.0181924f $X=-0.33 $Y=-0.265
+ $X2=2.885 $Y2=1.855
cc_92 N_VNB_M1011_b N_A_484_107#_c_1297_n 0.0231084f $X=-0.33 $Y=-0.265
+ $X2=2.885 $Y2=1.25
cc_93 N_VNB_M1011_b N_A_484_107#_c_1298_n 0.00663763f $X=-0.33 $Y=-0.265
+ $X2=1.115 $Y2=1.58
cc_94 N_VNB_M1011_b N_A_484_107#_c_1299_n 0.0109104f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_95 N_VNB_c_2_p N_A_484_107#_c_1299_n 8.65969e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_96 N_VNB_M1011_b N_A_484_107#_c_1301_n 2.20731e-19 $X=-0.33 $Y=-0.265
+ $X2=0.692 $Y2=1.38
cc_97 N_VNB_M1011_b N_A_484_107#_c_1302_n 0.00648341f $X=-0.33 $Y=-0.265
+ $X2=1.505 $Y2=1.735
cc_98 N_VNB_M1011_b N_Q_c_1392_n 0.0160961f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=3.175
cc_99 N_VNB_c_2_p N_Q_c_1392_n 8.28544e-19 $X=0.24 $Y=0 $X2=0.685 $Y2=3.175
cc_100 N_VNB_M1011_b N_Q_c_1394_n 0.00363283f $X=-0.33 $Y=-0.265 $X2=2.885
+ $Y2=1.855
cc_101 N_VNB_M1011_b Q 0.0188356f $X=-0.33 $Y=-0.265 $X2=0.635 $Y2=1.58
cc_102 N_VNB_M1011_b N_VGND_c_1430_n 0.0482941f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_103 N_VNB_c_2_p N_VGND_c_1430_n 0.00270129f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_104 N_VNB_M1011_b N_VGND_c_1432_n 0.0548945f $X=-0.33 $Y=-0.265 $X2=2.95
+ $Y2=1.25
cc_105 N_VNB_c_2_p N_VGND_c_1432_n 0.00256586f $X=0.24 $Y=0 $X2=2.95 $Y2=1.25
cc_106 N_VNB_M1011_b N_VGND_c_1434_n 0.0380477f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_107 N_VNB_c_2_p N_VGND_c_1434_n 0.00167165f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_108 N_VNB_M1011_b N_VGND_c_1436_n 0.0478162f $X=-0.33 $Y=-0.265 $X2=1.795
+ $Y2=1.735
cc_109 N_VNB_c_2_p N_VGND_c_1436_n 0.00268867f $X=0.24 $Y=0 $X2=1.795 $Y2=1.735
cc_110 N_VNB_M1011_b N_VGND_c_1438_n 0.0503599f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_111 N_VNB_c_2_p N_VGND_c_1438_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_112 N_VNB_M1011_b N_VGND_c_1440_n 0.0662666f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_113 N_VNB_c_2_p N_VGND_c_1440_n 0.00166879f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_114 N_VNB_M1011_b N_VGND_c_1442_n 0.195716f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_115 N_VNB_c_2_p N_VGND_c_1442_n 1.59109f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_116 N_VPB_M1003_b N_SCE_c_261_n 0.120654f $X=-0.33 $Y=1.885 $X2=0.695
+ $Y2=2.355
cc_117 N_VPB_M1003_b N_SCE_c_262_n 0.0799733f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.855
cc_118 VPB N_SCE_c_262_n 0.0102703f $X=0 $Y=3.955 $X2=0.685 $Y2=2.855
cc_119 N_VPB_c_119_p N_SCE_c_262_n 0.0217401f $X=14.64 $Y=4.07 $X2=0.685
+ $Y2=2.855
cc_120 N_VPB_M1003_b N_SCE_c_265_n 0.0746941f $X=-0.33 $Y=1.885 $X2=1.465
+ $Y2=2.855
cc_121 VPB N_SCE_c_265_n 0.0102703f $X=0 $Y=3.955 $X2=1.465 $Y2=2.855
cc_122 N_VPB_c_119_p N_SCE_c_265_n 0.0155394f $X=14.64 $Y=4.07 $X2=1.465
+ $Y2=2.855
cc_123 N_VPB_M1003_b N_SCE_c_254_n 0.00394111f $X=-0.33 $Y=1.885 $X2=2.72
+ $Y2=1.94
cc_124 N_VPB_M1003_b N_SCE_c_258_n 0.0206918f $X=-0.33 $Y=1.885 $X2=0.77
+ $Y2=1.565
cc_125 N_VPB_M1003_b N_SCE_c_259_n 0.00317485f $X=-0.33 $Y=1.885 $X2=1.505
+ $Y2=1.735
cc_126 N_VPB_M1003_b N_D_c_326_n 0.00694143f $X=-0.33 $Y=1.885 $X2=0.695
+ $Y2=2.355
cc_127 N_VPB_M1003_b N_D_M1016_g 0.04872f $X=-0.33 $Y=1.885 $X2=0.685 $Y2=3.175
cc_128 VPB N_D_M1016_g 0.00196852f $X=0 $Y=3.955 $X2=0.685 $Y2=3.175
cc_129 N_VPB_c_119_p N_D_M1016_g 0.00869308f $X=14.64 $Y=4.07 $X2=0.685
+ $Y2=3.175
cc_130 N_VPB_M1003_b D 0.0176132f $X=-0.33 $Y=1.885 $X2=2.72 $Y2=1.94
cc_131 N_VPB_M1003_b N_D_c_333_n 0.105594f $X=-0.33 $Y=1.885 $X2=1.115 $Y2=1.58
cc_132 N_VPB_M1003_b N_A_30_593#_M1006_g 0.0897964f $X=-0.33 $Y=1.885 $X2=1.465
+ $Y2=3.175
cc_133 VPB N_A_30_593#_M1006_g 0.00196852f $X=0 $Y=3.955 $X2=1.465 $Y2=3.175
cc_134 N_VPB_c_119_p N_A_30_593#_M1006_g 0.00869308f $X=14.64 $Y=4.07 $X2=1.465
+ $Y2=3.175
cc_135 N_VPB_M1003_b N_A_30_593#_c_374_n 0.0784522f $X=-0.33 $Y=1.885 $X2=2.885
+ $Y2=1.25
cc_136 N_VPB_c_119_p N_A_30_593#_c_374_n 0.00396086f $X=14.64 $Y=4.07 $X2=2.885
+ $Y2=1.25
cc_137 N_VPB_M1003_b N_A_30_593#_c_377_n 0.0733372f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_138 N_VPB_M1003_b N_SCD_M1007_g 0.0381249f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.855
cc_139 VPB N_SCD_M1007_g 8.70087e-19 $X=0 $Y=3.955 $X2=0.685 $Y2=2.855
cc_140 N_VPB_c_119_p N_SCD_M1007_g 0.00487832f $X=14.64 $Y=4.07 $X2=0.685
+ $Y2=2.855
cc_141 N_VPB_M1003_b SCD 0.0116197f $X=-0.33 $Y=1.885 $X2=0.685 $Y2=2.605
cc_142 N_VPB_M1003_b N_SCD_c_442_n 0.0670622f $X=-0.33 $Y=1.885 $X2=2.72
+ $Y2=1.94
cc_143 N_VPB_M1003_b N_SCD_c_437_n 0.0211142f $X=-0.33 $Y=1.885 $X2=2.885
+ $Y2=1.855
cc_144 N_VPB_M1003_b N_CLK_M1009_g 0.138883f $X=-0.33 $Y=1.885 $X2=0.695
+ $Y2=2.355
cc_145 VPB N_CLK_M1009_g 0.00970178f $X=0 $Y=3.955 $X2=0.695 $Y2=2.355
cc_146 N_VPB_c_119_p N_CLK_M1009_g 0.0159423f $X=14.64 $Y=4.07 $X2=0.695
+ $Y2=2.355
cc_147 N_VPB_M1003_b N_A_1204_107#_c_525_n 0.0991564f $X=-0.33 $Y=1.885
+ $X2=0.685 $Y2=2.855
cc_148 N_VPB_M1003_b N_A_1204_107#_M1023_g 0.0925197f $X=-0.33 $Y=1.885 $X2=2.72
+ $Y2=1.94
cc_149 N_VPB_M1003_b N_A_1204_107#_c_527_n 0.0187242f $X=-0.33 $Y=1.885
+ $X2=1.115 $Y2=1.58
cc_150 N_VPB_M1003_b N_A_1204_107#_c_528_n 0.0276693f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_151 VPB N_A_1204_107#_c_528_n 0.00195181f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_152 N_VPB_c_119_p N_A_1204_107#_c_528_n 0.0200897f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_153 N_VPB_M1003_b N_A_1204_107#_c_531_n 0.00507615f $X=-0.33 $Y=1.885
+ $X2=2.95 $Y2=0.745
cc_154 VPB N_A_1204_107#_c_531_n 0.00102583f $X=0 $Y=3.955 $X2=2.95 $Y2=0.745
cc_155 N_VPB_c_119_p N_A_1204_107#_c_531_n 0.0159324f $X=14.64 $Y=4.07 $X2=2.95
+ $Y2=0.745
cc_156 N_VPB_M1003_b N_A_1204_107#_c_534_n 0.00474079f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_157 N_VPB_M1003_b N_A_1204_107#_c_535_n 2.01647e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_158 N_VPB_M1003_b N_A_1204_107#_c_536_n 0.00405326f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_159 N_VPB_M1003_b N_A_1204_107#_c_524_n 0.0408535f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_160 N_VPB_M1003_b N_A_938_107#_c_659_n 0.150805f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.855
cc_161 N_VPB_M1003_b N_A_938_107#_M1020_g 0.0443533f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=3.175
cc_162 VPB N_A_938_107#_M1020_g 0.00970178f $X=0 $Y=3.955 $X2=0.685 $Y2=3.175
cc_163 N_VPB_c_119_p N_A_938_107#_M1020_g 0.016048f $X=14.64 $Y=4.07 $X2=0.685
+ $Y2=3.175
cc_164 N_VPB_M1003_b N_A_938_107#_c_660_n 0.0319491f $X=-0.33 $Y=1.885 $X2=1.465
+ $Y2=3.175
cc_165 N_VPB_M1003_b N_A_938_107#_M1024_g 0.0763458f $X=-0.33 $Y=1.885 $X2=2.885
+ $Y2=1.25
cc_166 N_VPB_M1003_b N_A_938_107#_c_679_n 0.0109342f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_167 VPB N_A_938_107#_c_679_n 0.00101808f $X=0 $Y=3.955 $X2=0.635 $Y2=1.58
cc_168 N_VPB_c_119_p N_A_938_107#_c_679_n 0.0158392f $X=14.64 $Y=4.07 $X2=0.635
+ $Y2=1.58
cc_169 N_VPB_M1003_b N_A_938_107#_c_682_n 0.0079008f $X=-0.33 $Y=1.885 $X2=2.95
+ $Y2=0.745
cc_170 N_VPB_M1003_b N_A_938_107#_c_683_n 0.00548137f $X=-0.33 $Y=1.885 $X2=2.95
+ $Y2=0.745
cc_171 N_VPB_M1003_b N_A_938_107#_c_684_n 0.0201955f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_172 N_VPB_c_119_p N_A_938_107#_c_684_n 0.0121557f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_173 N_VPB_M1003_b N_A_938_107#_c_686_n 0.00452024f $X=-0.33 $Y=1.885 $X2=1.68
+ $Y2=1.735
cc_174 N_VPB_c_119_p N_A_938_107#_c_686_n 0.00206641f $X=14.64 $Y=4.07 $X2=1.68
+ $Y2=1.735
cc_175 N_VPB_M1003_b N_A_938_107#_c_688_n 0.0113589f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_176 VPB N_A_938_107#_c_688_n 0.00224212f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_177 N_VPB_c_119_p N_A_938_107#_c_688_n 0.0197679f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_178 N_VPB_M1003_b N_A_938_107#_c_665_n 0.00175093f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_179 N_VPB_M1003_b N_A_938_107#_c_692_n 0.0839476f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_180 VPB N_A_938_107#_c_692_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_181 N_VPB_c_119_p N_A_938_107#_c_692_n 0.0151198f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_182 VPB N_A_938_107#_c_695_n 7.18582e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_183 N_VPB_c_119_p N_A_938_107#_c_695_n 0.00307385f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_184 N_VPB_M1003_b N_A_938_107#_c_672_n 0.05226f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_185 N_VPB_M1003_b N_A_1688_81#_M1026_g 0.0371353f $X=-0.33 $Y=1.885 $X2=1.465
+ $Y2=3.175
cc_186 N_VPB_M1003_b N_A_1688_81#_c_860_n 0.0159885f $X=-0.33 $Y=1.885 $X2=2.885
+ $Y2=1.25
cc_187 N_VPB_M1003_b N_A_1688_81#_c_861_n 0.00855036f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_188 N_VPB_M1003_b N_A_1688_81#_c_857_n 0.067254f $X=-0.33 $Y=1.885 $X2=0.77
+ $Y2=1.565
cc_189 N_VPB_M1003_b N_A_1688_81#_c_863_n 0.00222833f $X=-0.33 $Y=1.885 $X2=0.77
+ $Y2=1.565
cc_190 N_VPB_M1003_b N_A_1688_81#_c_864_n 0.0016195f $X=-0.33 $Y=1.885 $X2=0.692
+ $Y2=2.09
cc_191 N_VPB_M1003_b N_A_1688_81#_c_865_n 0.00613488f $X=-0.33 $Y=1.885
+ $X2=1.505 $Y2=1.735
cc_192 N_VPB_M1003_b N_A_1490_107#_c_942_n 0.00113231f $X=-0.33 $Y=1.885
+ $X2=1.465 $Y2=3.175
cc_193 N_VPB_M1003_b N_A_1490_107#_c_943_n 0.00351869f $X=-0.33 $Y=1.885
+ $X2=0.685 $Y2=2.605
cc_194 N_VPB_M1003_b N_A_1490_107#_c_944_n 0.0114219f $X=-0.33 $Y=1.885
+ $X2=1.595 $Y2=1.58
cc_195 N_VPB_M1003_b N_A_1490_107#_M1013_g 0.10283f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_196 VPB N_A_1490_107#_M1013_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_197 N_VPB_c_119_p N_A_1490_107#_M1013_g 0.013715f $X=14.64 $Y=4.07 $X2=0
+ $Y2=0
cc_198 N_VPB_M1003_b N_A_2352_81#_M1004_g 0.0748724f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.605
cc_199 N_VPB_M1003_b N_A_2352_81#_M1010_g 0.0462427f $X=-0.33 $Y=1.885 $X2=2.885
+ $Y2=1.25
cc_200 VPB N_A_2352_81#_M1010_g 0.00970178f $X=0 $Y=3.955 $X2=2.885 $Y2=1.25
cc_201 N_VPB_c_119_p N_A_2352_81#_M1010_g 0.0159423f $X=14.64 $Y=4.07 $X2=2.885
+ $Y2=1.25
cc_202 N_VPB_M1003_b N_A_2352_81#_c_1016_n 0.0377376f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=1.58
cc_203 N_VPB_M1003_b N_A_2352_81#_c_1017_n 0.0216672f $X=-0.33 $Y=1.885
+ $X2=1.115 $Y2=1.58
cc_204 N_VPB_M1003_b N_A_2352_81#_c_1029_n 0.0173924f $X=-0.33 $Y=1.885 $X2=0.77
+ $Y2=1.565
cc_205 VPB N_A_2352_81#_c_1029_n 0.00101808f $X=0 $Y=3.955 $X2=0.77 $Y2=1.565
cc_206 N_VPB_c_119_p N_A_2352_81#_c_1029_n 0.0158392f $X=14.64 $Y=4.07 $X2=0.77
+ $Y2=1.565
cc_207 N_VPB_M1003_b N_A_2352_81#_c_1022_n 0.0282418f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_208 N_VPB_M1003_b N_A_2123_543#_M1005_g 0.0427937f $X=-0.33 $Y=1.885
+ $X2=0.685 $Y2=2.605
cc_209 VPB N_A_2123_543#_M1005_g 0.00970178f $X=0 $Y=3.955 $X2=0.685 $Y2=2.605
cc_210 N_VPB_c_119_p N_A_2123_543#_M1005_g 0.0159423f $X=14.64 $Y=4.07 $X2=0.685
+ $Y2=2.605
cc_211 N_VPB_M1003_b N_A_2123_543#_c_1107_n 0.00861203f $X=-0.33 $Y=1.885
+ $X2=2.885 $Y2=1.855
cc_212 N_VPB_M1003_b N_A_2123_543#_c_1112_n 0.00274942f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_213 N_VPB_M1003_b N_A_2123_543#_c_1119_n 0.0120852f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=1.58
cc_214 N_VPB_M1003_b N_A_2123_543#_c_1120_n 0.00629486f $X=-0.33 $Y=1.885
+ $X2=1.115 $Y2=1.58
cc_215 N_VPB_M1003_b N_A_2123_543#_c_1113_n 0.071998f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_216 N_VPB_M1003_b N_A_2123_543#_c_1122_n 0.00445269f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_217 N_VPB_M1003_b N_VPWR_c_1201_n 0.0111733f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1201_n 0.0036893f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_219 N_VPB_c_119_p N_VPWR_c_1201_n 0.0389096f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_220 N_VPB_M1003_b N_VPWR_c_1204_n 0.0130587f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1204_n 0.00334907f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_222 N_VPB_c_119_p N_VPWR_c_1204_n 0.0448889f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_223 N_VPB_M1003_b N_VPWR_c_1207_n 0.00992943f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1207_n 0.00226124f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_225 N_VPB_c_119_p N_VPWR_c_1207_n 0.0274397f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_226 N_VPB_M1003_b N_VPWR_c_1210_n 0.00613063f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1210_n 0.00360667f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_228 N_VPB_c_119_p N_VPWR_c_1210_n 0.0475243f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_229 N_VPB_M1003_b N_VPWR_c_1213_n 0.0169208f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1213_n 0.00334907f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_231 N_VPB_c_119_p N_VPWR_c_1213_n 0.0448889f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_232 N_VPB_M1003_b N_VPWR_c_1216_n 0.0641347f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1216_n 0.00222504f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_234 N_VPB_c_119_p N_VPWR_c_1216_n 0.0275189f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_235 N_VPB_M1003_b N_VPWR_c_1219_n 0.168999f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1219_n 1.5853f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_237 N_VPB_c_119_p N_VPWR_c_1219_n 0.0749202f $X=14.64 $Y=4.07 $X2=0 $Y2=0
cc_238 N_VPB_M1003_b N_A_484_107#_c_1303_n 0.00117313f $X=-0.33 $Y=1.885
+ $X2=1.465 $Y2=2.855
cc_239 N_VPB_M1003_b N_A_484_107#_c_1304_n 0.0178262f $X=-0.33 $Y=1.885
+ $X2=2.885 $Y2=1.25
cc_240 N_VPB_M1003_b N_A_484_107#_c_1297_n 0.0335932f $X=-0.33 $Y=1.885
+ $X2=2.885 $Y2=1.25
cc_241 N_VPB_M1003_b N_A_484_107#_c_1306_n 0.00612984f $X=-0.33 $Y=1.885
+ $X2=2.95 $Y2=1.25
cc_242 N_VPB_c_119_p N_A_484_107#_c_1306_n 0.00494722f $X=14.64 $Y=4.07 $X2=2.95
+ $Y2=1.25
cc_243 N_VPB_M1003_b N_A_484_107#_c_1301_n 0.00152417f $X=-0.33 $Y=1.885
+ $X2=0.692 $Y2=1.38
cc_244 N_VPB_M1003_b N_A_484_107#_c_1309_n 0.00229761f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_245 N_VPB_M1003_b N_A_484_107#_c_1310_n 0.0111757f $X=-0.33 $Y=1.885 $X2=1.2
+ $Y2=1.735
cc_246 N_VPB_M1003_b N_A_484_107#_c_1311_n 0.016672f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_247 N_VPB_M1003_b N_Q_c_1396_n 0.0132716f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.605
cc_248 VPB N_Q_c_1396_n 0.00116152f $X=0 $Y=3.955 $X2=0.685 $Y2=2.605
cc_249 N_VPB_c_119_p N_Q_c_1396_n 0.0171777f $X=14.64 $Y=4.07 $X2=0.685
+ $Y2=2.605
cc_250 N_VPB_M1003_b N_Q_c_1399_n 0.00365505f $X=-0.33 $Y=1.885 $X2=2.885
+ $Y2=1.25
cc_251 N_VPB_M1003_b N_Q_c_1400_n 0.00143467f $X=-0.33 $Y=1.885 $X2=2.885
+ $Y2=1.25
cc_252 N_SCE_M1011_g N_D_M1025_g 0.0307827f $X=0.68 $Y=0.745 $X2=0 $Y2=0
cc_253 N_SCE_c_258_n N_D_c_326_n 0.0122112f $X=0.77 $Y=1.565 $X2=0 $Y2=0
cc_254 N_SCE_c_259_n N_D_c_326_n 0.0117584f $X=1.505 $Y=1.735 $X2=0 $Y2=0
cc_255 N_SCE_c_260_n N_D_c_326_n 0.010648f $X=1.795 $Y=1.735 $X2=0 $Y2=0
cc_256 N_SCE_c_265_n N_D_M1016_g 0.0286352f $X=1.465 $Y=2.855 $X2=0 $Y2=0
cc_257 N_SCE_c_258_n N_D_c_327_n 0.0115185f $X=0.77 $Y=1.565 $X2=0.24 $Y2=0
cc_258 N_SCE_c_259_n N_D_c_327_n 0.0129235f $X=1.505 $Y=1.735 $X2=0.24 $Y2=0
cc_259 N_SCE_c_260_n N_D_c_327_n 0.00627549f $X=1.795 $Y=1.735 $X2=0.24 $Y2=0
cc_260 N_SCE_c_261_n D 0.0585217f $X=0.695 $Y=2.355 $X2=14.64 $Y2=0
cc_261 N_SCE_c_254_n D 0.00265902f $X=2.72 $Y=1.94 $X2=14.64 $Y2=0
cc_262 N_SCE_c_259_n D 0.157772f $X=1.505 $Y=1.735 $X2=14.64 $Y2=0
cc_263 N_SCE_c_261_n N_D_c_333_n 0.0726299f $X=0.695 $Y=2.355 $X2=0 $Y2=0
cc_264 N_SCE_c_254_n N_D_c_333_n 0.00563519f $X=2.72 $Y=1.94 $X2=0 $Y2=0
cc_265 N_SCE_c_259_n N_D_c_333_n 0.00331157f $X=1.505 $Y=1.735 $X2=0 $Y2=0
cc_266 N_SCE_c_260_n N_D_c_333_n 0.00723605f $X=1.795 $Y=1.735 $X2=0 $Y2=0
cc_267 N_SCE_M1015_g N_A_30_593#_c_370_n 0.0147942f $X=2.95 $Y=0.745 $X2=0 $Y2=0
cc_268 N_SCE_M1011_g N_A_30_593#_c_372_n 0.0221394f $X=0.68 $Y=0.745 $X2=14.64
+ $Y2=0
cc_269 N_SCE_M1011_g N_A_30_593#_c_374_n 0.0287144f $X=0.68 $Y=0.745 $X2=0 $Y2=0
cc_270 N_SCE_c_261_n N_A_30_593#_c_374_n 0.0379951f $X=0.695 $Y=2.355 $X2=0
+ $Y2=0
cc_271 N_SCE_c_259_n N_A_30_593#_c_374_n 0.0384963f $X=1.505 $Y=1.735 $X2=0
+ $Y2=0
cc_272 N_SCE_M1011_g N_A_30_593#_c_375_n 0.030661f $X=0.68 $Y=0.745 $X2=0 $Y2=0
cc_273 N_SCE_c_254_n N_A_30_593#_c_375_n 0.00546307f $X=2.72 $Y=1.94 $X2=0 $Y2=0
cc_274 N_SCE_c_258_n N_A_30_593#_c_375_n 7.0593e-19 $X=0.77 $Y=1.565 $X2=0 $Y2=0
cc_275 N_SCE_c_259_n N_A_30_593#_c_375_n 0.0878811f $X=1.505 $Y=1.735 $X2=0
+ $Y2=0
cc_276 N_SCE_M1011_g N_A_30_593#_c_376_n 0.00513266f $X=0.68 $Y=0.745 $X2=0
+ $Y2=0
cc_277 N_SCE_c_254_n N_A_30_593#_c_394_n 0.0237472f $X=2.72 $Y=1.94 $X2=0 $Y2=0
cc_278 N_SCE_c_255_n N_A_30_593#_c_394_n 0.0215354f $X=2.885 $Y=1.25 $X2=0 $Y2=0
cc_279 N_SCE_M1015_g N_A_30_593#_c_394_n 0.0016635f $X=2.95 $Y=0.745 $X2=0 $Y2=0
cc_280 N_SCE_c_260_n N_A_30_593#_c_394_n 0.018497f $X=1.795 $Y=1.735 $X2=0 $Y2=0
cc_281 N_SCE_c_254_n N_A_30_593#_c_377_n 0.0576291f $X=2.72 $Y=1.94 $X2=0 $Y2=0
cc_282 N_SCE_c_255_n N_A_30_593#_c_377_n 0.00627304f $X=2.885 $Y=1.25 $X2=0
+ $Y2=0
cc_283 N_SCE_M1015_g N_A_30_593#_c_377_n 0.0845977f $X=2.95 $Y=0.745 $X2=0 $Y2=0
cc_284 N_SCE_c_260_n N_A_30_593#_c_377_n 0.00675269f $X=1.795 $Y=1.735 $X2=0
+ $Y2=0
cc_285 N_SCE_M1015_g N_SCD_M1018_g 0.0770814f $X=2.95 $Y=0.745 $X2=0 $Y2=0
cc_286 N_SCE_c_254_n N_SCD_c_437_n 6.38034e-19 $X=2.72 $Y=1.94 $X2=0 $Y2=0
cc_287 N_SCE_M1015_g N_SCD_c_437_n 0.00930842f $X=2.95 $Y=0.745 $X2=0 $Y2=0
cc_288 N_SCE_c_261_n N_VPWR_c_1201_n 0.00328723f $X=0.695 $Y=2.355 $X2=0 $Y2=0
cc_289 N_SCE_c_262_n N_VPWR_c_1201_n 0.0255844f $X=0.685 $Y=2.855 $X2=0 $Y2=0
cc_290 N_SCE_c_265_n N_VPWR_c_1201_n 0.0605197f $X=1.465 $Y=2.855 $X2=0 $Y2=0
cc_291 N_SCE_c_262_n N_VPWR_c_1219_n 0.0348123f $X=0.685 $Y=2.855 $X2=0 $Y2=0
cc_292 N_SCE_c_265_n N_VPWR_c_1219_n 0.00415815f $X=1.465 $Y=2.855 $X2=0 $Y2=0
cc_293 N_SCE_c_255_n N_A_484_107#_c_1295_n 0.0223991f $X=2.885 $Y=1.25 $X2=0
+ $Y2=0
cc_294 N_SCE_M1015_g N_A_484_107#_c_1295_n 0.0302092f $X=2.95 $Y=0.745 $X2=0
+ $Y2=0
cc_295 N_SCE_c_254_n N_A_484_107#_c_1296_n 7.74718e-19 $X=2.72 $Y=1.94 $X2=0
+ $Y2=0
cc_296 N_SCE_c_255_n N_A_484_107#_c_1296_n 0.0549953f $X=2.885 $Y=1.25 $X2=0
+ $Y2=0
cc_297 N_SCE_M1015_g N_A_484_107#_c_1296_n 0.00893478f $X=2.95 $Y=0.745 $X2=0
+ $Y2=0
cc_298 N_SCE_M1015_g N_A_484_107#_c_1299_n 0.00904648f $X=2.95 $Y=0.745 $X2=0
+ $Y2=0
cc_299 N_SCE_c_265_n N_A_484_107#_c_1306_n 2.95467e-19 $X=1.465 $Y=2.855 $X2=0
+ $Y2=0
cc_300 N_SCE_c_254_n N_A_484_107#_c_1301_n 0.0142079f $X=2.72 $Y=1.94 $X2=0
+ $Y2=0
cc_301 N_SCE_M1011_g N_VGND_c_1430_n 0.01513f $X=0.68 $Y=0.745 $X2=0 $Y2=0
cc_302 N_SCE_M1015_g N_VGND_c_1432_n 0.00260392f $X=2.95 $Y=0.745 $X2=0 $Y2=0
cc_303 N_SCE_M1011_g N_VGND_c_1442_n 0.0153615f $X=0.68 $Y=0.745 $X2=0 $Y2=0
cc_304 N_SCE_c_255_n N_VGND_c_1442_n 6.68981e-19 $X=2.885 $Y=1.25 $X2=0 $Y2=0
cc_305 N_SCE_M1015_g N_VGND_c_1442_n 0.0151022f $X=2.95 $Y=0.745 $X2=0 $Y2=0
cc_306 N_D_M1025_g N_A_30_593#_c_370_n 0.0467316f $X=1.46 $Y=0.745 $X2=0 $Y2=0
cc_307 D N_A_30_593#_M1006_g 0.012113f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_308 N_D_c_333_n N_A_30_593#_M1006_g 0.0394873f $X=1.635 $Y=2.29 $X2=0 $Y2=0
cc_309 D N_A_30_593#_c_374_n 0.0208131f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_310 N_D_M1025_g N_A_30_593#_c_375_n 0.0254861f $X=1.46 $Y=0.745 $X2=0 $Y2=0
cc_311 N_D_M1025_g N_A_30_593#_c_394_n 0.0011719f $X=1.46 $Y=0.745 $X2=0 $Y2=0
cc_312 N_D_c_327_n N_A_30_593#_c_394_n 2.20562e-19 $X=1.46 $Y=1.585 $X2=0 $Y2=0
cc_313 N_D_c_326_n N_A_30_593#_c_377_n 0.00795011f $X=1.532 $Y=1.985 $X2=0 $Y2=0
cc_314 N_D_c_327_n N_A_30_593#_c_377_n 0.0467316f $X=1.46 $Y=1.585 $X2=0 $Y2=0
cc_315 D N_A_30_593#_c_377_n 0.0177903f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_316 N_D_c_333_n N_A_30_593#_c_377_n 0.0310375f $X=1.635 $Y=2.29 $X2=0 $Y2=0
cc_317 N_D_M1016_g N_VPWR_c_1201_n 0.00943955f $X=2.175 $Y=3.175 $X2=0 $Y2=0
cc_318 D N_VPWR_c_1201_n 0.0422669f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_319 N_D_c_333_n N_VPWR_c_1201_n 0.00123599f $X=1.635 $Y=2.29 $X2=0 $Y2=0
cc_320 N_D_M1016_g N_VPWR_c_1219_n 0.0300945f $X=2.175 $Y=3.175 $X2=0 $Y2=0
cc_321 D N_A_484_107#_c_1303_n 8.83448e-19 $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_322 D N_A_484_107#_c_1304_n 0.0114316f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_323 N_D_M1025_g N_A_484_107#_c_1299_n 3.16053e-19 $X=1.46 $Y=0.745 $X2=0
+ $Y2=0
cc_324 N_D_M1016_g N_A_484_107#_c_1306_n 0.0142509f $X=2.175 $Y=3.175 $X2=0
+ $Y2=0
cc_325 D N_A_484_107#_c_1306_n 0.0150422f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_326 N_D_M1025_g N_VGND_c_1430_n 0.0432487f $X=1.46 $Y=0.745 $X2=0 $Y2=0
cc_327 N_A_30_593#_M1006_g N_SCD_M1007_g 0.0460415f $X=2.955 $Y=3.175 $X2=0
+ $Y2=0
cc_328 N_A_30_593#_c_377_n N_SCD_c_442_n 0.0460415f $X=2.17 $Y=1.525 $X2=14.64
+ $Y2=0
cc_329 N_A_30_593#_c_377_n N_SCD_c_437_n 0.00681621f $X=2.17 $Y=1.525 $X2=0
+ $Y2=0
cc_330 N_A_30_593#_c_374_n N_VPWR_c_1201_n 0.00966689f $X=0.295 $Y=3.175 $X2=0
+ $Y2=0
cc_331 N_A_30_593#_M1006_g N_VPWR_c_1204_n 0.00225495f $X=2.955 $Y=3.175 $X2=0
+ $Y2=0
cc_332 N_A_30_593#_M1006_g N_VPWR_c_1219_n 0.0145717f $X=2.955 $Y=3.175 $X2=0
+ $Y2=0
cc_333 N_A_30_593#_c_374_n N_VPWR_c_1219_n 0.0115855f $X=0.295 $Y=3.175 $X2=0
+ $Y2=0
cc_334 N_A_30_593#_M1006_g N_A_484_107#_c_1303_n 0.0379591f $X=2.955 $Y=3.175
+ $X2=0 $Y2=0
cc_335 N_A_30_593#_c_377_n N_A_484_107#_c_1304_n 0.0181359f $X=2.17 $Y=1.525
+ $X2=0 $Y2=0
cc_336 N_A_30_593#_c_370_n N_A_484_107#_c_1299_n 0.0115285f $X=2.17 $Y=1.065
+ $X2=0 $Y2=0
cc_337 N_A_30_593#_c_377_n N_A_484_107#_c_1299_n 0.00201476f $X=2.17 $Y=1.525
+ $X2=0 $Y2=0
cc_338 N_A_30_593#_M1006_g N_A_484_107#_c_1306_n 0.0111426f $X=2.955 $Y=3.175
+ $X2=0 $Y2=0
cc_339 N_A_30_593#_c_377_n N_A_484_107#_c_1306_n 0.00123442f $X=2.17 $Y=1.525
+ $X2=0 $Y2=0
cc_340 N_A_30_593#_c_377_n N_A_484_107#_c_1301_n 7.41409e-19 $X=2.17 $Y=1.525
+ $X2=0 $Y2=0
cc_341 N_A_30_593#_c_370_n N_VGND_c_1430_n 0.00760888f $X=2.17 $Y=1.065 $X2=0
+ $Y2=0
cc_342 N_A_30_593#_c_372_n N_VGND_c_1430_n 0.01253f $X=0.29 $Y=0.745 $X2=0 $Y2=0
cc_343 N_A_30_593#_c_375_n N_VGND_c_1430_n 0.0602349f $X=1.975 $Y=1.18 $X2=0
+ $Y2=0
cc_344 N_A_30_593#_c_370_n N_VGND_c_1442_n 0.0198175f $X=2.17 $Y=1.065 $X2=0
+ $Y2=0
cc_345 N_A_30_593#_c_372_n N_VGND_c_1442_n 0.033134f $X=0.29 $Y=0.745 $X2=0
+ $Y2=0
cc_346 N_A_30_593#_c_375_n N_VGND_c_1442_n 0.0213269f $X=1.975 $Y=1.18 $X2=0
+ $Y2=0
cc_347 N_A_30_593#_c_394_n N_VGND_c_1442_n 0.0114007f $X=2.14 $Y=1.25 $X2=0
+ $Y2=0
cc_348 N_SCD_M1007_g N_CLK_M1009_g 0.0152868f $X=3.665 $Y=3.175 $X2=0 $Y2=0
cc_349 SCD N_CLK_M1009_g 0.0144756f $X=3.995 $Y=2.32 $X2=0 $Y2=0
cc_350 N_SCD_c_437_n N_CLK_M1009_g 0.0414228f $X=3.682 $Y=2.115 $X2=0 $Y2=0
cc_351 N_SCD_c_436_n CLK 0.00270932f $X=3.68 $Y=1.585 $X2=0 $Y2=0
cc_352 N_SCD_c_436_n N_CLK_c_477_n 0.0470255f $X=3.68 $Y=1.585 $X2=0.24 $Y2=0
cc_353 N_SCD_M1018_g N_CLK_c_478_n 0.0145485f $X=3.66 $Y=0.745 $X2=0 $Y2=0
cc_354 SCD N_A_938_107#_c_683_n 0.00591205f $X=3.995 $Y=2.32 $X2=0 $Y2=0
cc_355 N_SCD_M1007_g N_VPWR_c_1204_n 0.042487f $X=3.665 $Y=3.175 $X2=0 $Y2=0
cc_356 SCD N_VPWR_c_1204_n 0.0466141f $X=3.995 $Y=2.32 $X2=0 $Y2=0
cc_357 N_SCD_c_442_n N_VPWR_c_1204_n 0.00103072f $X=3.765 $Y=2.3 $X2=0 $Y2=0
cc_358 N_SCD_M1007_g N_VPWR_c_1219_n 0.0134149f $X=3.665 $Y=3.175 $X2=0 $Y2=0
cc_359 N_SCD_M1007_g N_A_484_107#_c_1303_n 0.00146371f $X=3.665 $Y=3.175 $X2=0
+ $Y2=0
cc_360 N_SCD_M1018_g N_A_484_107#_c_1296_n 0.0155071f $X=3.66 $Y=0.745 $X2=0
+ $Y2=0
cc_361 N_SCD_c_437_n N_A_484_107#_c_1296_n 0.00875248f $X=3.682 $Y=2.115 $X2=0
+ $Y2=0
cc_362 SCD N_A_484_107#_c_1304_n 0.0382989f $X=3.995 $Y=2.32 $X2=0 $Y2=0
cc_363 N_SCD_c_442_n N_A_484_107#_c_1304_n 0.0110978f $X=3.765 $Y=2.3 $X2=0
+ $Y2=0
cc_364 N_SCD_c_437_n N_A_484_107#_c_1304_n 0.00195415f $X=3.682 $Y=2.115 $X2=0
+ $Y2=0
cc_365 N_SCD_c_436_n N_A_484_107#_c_1297_n 9.59793e-19 $X=3.68 $Y=1.585 $X2=7.44
+ $Y2=0
cc_366 SCD N_A_484_107#_c_1297_n 0.0443377f $X=3.995 $Y=2.32 $X2=7.44 $Y2=0
cc_367 N_SCD_c_442_n N_A_484_107#_c_1297_n 0.00101157f $X=3.765 $Y=2.3 $X2=7.44
+ $Y2=0
cc_368 N_SCD_c_437_n N_A_484_107#_c_1297_n 0.0465569f $X=3.682 $Y=2.115 $X2=7.44
+ $Y2=0
cc_369 N_SCD_M1018_g N_A_484_107#_c_1299_n 9.53229e-19 $X=3.66 $Y=0.745 $X2=0
+ $Y2=0
cc_370 N_SCD_M1007_g N_A_484_107#_c_1306_n 0.00101042f $X=3.665 $Y=3.175 $X2=0
+ $Y2=0
cc_371 N_SCD_M1018_g N_VGND_c_1432_n 0.0511636f $X=3.66 $Y=0.745 $X2=0 $Y2=0
cc_372 N_SCD_c_436_n N_VGND_c_1432_n 0.00207972f $X=3.68 $Y=1.585 $X2=0 $Y2=0
cc_373 N_SCD_M1018_g N_VGND_c_1442_n 0.0112937f $X=3.66 $Y=0.745 $X2=0 $Y2=0
cc_374 N_CLK_M1009_g N_A_938_107#_c_659_n 0.0217141f $X=4.54 $Y=3.34 $X2=0 $Y2=0
cc_375 N_CLK_M1009_g N_A_938_107#_c_679_n 0.0252223f $X=4.54 $Y=3.34 $X2=7.44
+ $Y2=0.057
cc_376 N_CLK_c_477_n N_A_938_107#_c_662_n 0.0036153f $X=4.51 $Y=1.26 $X2=0 $Y2=0
cc_377 N_CLK_c_478_n N_A_938_107#_c_662_n 0.00369253f $X=4.49 $Y=1.075 $X2=0
+ $Y2=0
cc_378 CLK N_A_938_107#_c_664_n 0.012115f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_379 N_CLK_c_477_n N_A_938_107#_c_664_n 0.00556357f $X=4.51 $Y=1.26 $X2=0
+ $Y2=0
cc_380 N_CLK_M1009_g N_A_938_107#_c_683_n 0.00803589f $X=4.54 $Y=3.34 $X2=0
+ $Y2=0
cc_381 N_CLK_M1009_g N_A_938_107#_c_706_n 0.00236779f $X=4.54 $Y=3.34 $X2=0
+ $Y2=0
cc_382 CLK N_A_938_107#_c_666_n 5.38903e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_383 N_CLK_c_477_n N_A_938_107#_c_666_n 0.00496743f $X=4.51 $Y=1.26 $X2=0
+ $Y2=0
cc_384 N_CLK_c_478_n N_A_938_107#_c_666_n 0.00955273f $X=4.49 $Y=1.075 $X2=0
+ $Y2=0
cc_385 N_CLK_M1009_g N_VPWR_c_1204_n 0.0502683f $X=4.54 $Y=3.34 $X2=0 $Y2=0
cc_386 N_CLK_M1009_g N_VPWR_c_1207_n 0.00150546f $X=4.54 $Y=3.34 $X2=0 $Y2=0
cc_387 N_CLK_M1009_g N_VPWR_c_1219_n 0.0120207f $X=4.54 $Y=3.34 $X2=0 $Y2=0
cc_388 N_CLK_M1009_g N_A_484_107#_c_1297_n 0.048309f $X=4.54 $Y=3.34 $X2=7.44
+ $Y2=0
cc_389 CLK N_A_484_107#_c_1297_n 0.0232944f $X=4.475 $Y=1.21 $X2=7.44 $Y2=0
cc_390 N_CLK_c_477_n N_A_484_107#_c_1297_n 0.00457782f $X=4.51 $Y=1.26 $X2=7.44
+ $Y2=0
cc_391 CLK N_VGND_c_1432_n 0.0104912f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_392 N_CLK_c_478_n N_VGND_c_1432_n 0.0417791f $X=4.49 $Y=1.075 $X2=0 $Y2=0
cc_393 N_CLK_c_478_n N_VGND_c_1434_n 0.00269622f $X=4.49 $Y=1.075 $X2=0 $Y2=0
cc_394 CLK N_VGND_c_1442_n 0.0062095f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_395 N_CLK_c_478_n N_VGND_c_1442_n 0.006838f $X=4.49 $Y=1.075 $X2=0 $Y2=0
cc_396 N_A_1204_107#_c_525_n N_A_938_107#_c_659_n 0.00489044f $X=7.2 $Y=2.605
+ $X2=0 $Y2=0
cc_397 N_A_1204_107#_c_513_n N_A_938_107#_c_659_n 0.00897608f $X=6.16 $Y=0.745
+ $X2=0 $Y2=0
cc_398 N_A_1204_107#_c_527_n N_A_938_107#_M1020_g 0.00886872f $X=6.26 $Y=3.11
+ $X2=0 $Y2=0
cc_399 N_A_1204_107#_c_531_n N_A_938_107#_M1020_g 0.00655318f $X=6.425 $Y=3.42
+ $X2=0 $Y2=0
cc_400 N_A_1204_107#_c_525_n N_A_938_107#_c_660_n 0.0365723f $X=7.2 $Y=2.605
+ $X2=0.24 $Y2=0
cc_401 N_A_1204_107#_c_513_n N_A_938_107#_M1028_g 0.00300225f $X=6.16 $Y=0.745
+ $X2=0 $Y2=0
cc_402 N_A_1204_107#_c_514_n N_A_938_107#_M1028_g 0.00616595f $X=7.075 $Y=0.35
+ $X2=0 $Y2=0
cc_403 N_A_1204_107#_c_518_n N_A_938_107#_M1028_g 0.00891555f $X=7.935 $Y=0.35
+ $X2=0 $Y2=0
cc_404 N_A_1204_107#_c_546_p N_A_938_107#_M1028_g 0.00125202f $X=8.045 $Y=1.25
+ $X2=0 $Y2=0
cc_405 N_A_1204_107#_c_536_n N_A_938_107#_M1028_g 0.0352906f $X=7.142 $Y=2.225
+ $X2=0 $Y2=0
cc_406 N_A_1204_107#_c_521_n N_A_938_107#_M1028_g 0.00339519f $X=7.16 $Y=0.35
+ $X2=0 $Y2=0
cc_407 N_A_1204_107#_M1021_g N_A_938_107#_M1028_g 0.0224793f $X=7.98 $Y=0.745
+ $X2=0 $Y2=0
cc_408 N_A_1204_107#_c_525_n N_A_938_107#_M1024_g 0.0288809f $X=7.2 $Y=2.605
+ $X2=0 $Y2=0
cc_409 N_A_1204_107#_c_534_n N_A_938_107#_M1024_g 7.04648e-19 $X=7.24 $Y=3.335
+ $X2=0 $Y2=0
cc_410 N_A_1204_107#_c_525_n N_A_938_107#_c_686_n 3.66173e-19 $X=7.2 $Y=2.605
+ $X2=0 $Y2=0
cc_411 N_A_1204_107#_M1023_g N_A_938_107#_c_725_n 0.00112355f $X=11.26 $Y=2.925
+ $X2=0 $Y2=0
cc_412 N_A_1204_107#_M1023_g N_A_938_107#_c_688_n 0.0103627f $X=11.26 $Y=2.925
+ $X2=0 $Y2=0
cc_413 N_A_1204_107#_M1023_g N_A_938_107#_c_665_n 0.0582338f $X=11.26 $Y=2.925
+ $X2=0 $Y2=0
cc_414 N_A_1204_107#_c_524_n N_A_938_107#_c_665_n 0.0153158f $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_415 N_A_1204_107#_M1023_g N_A_938_107#_c_692_n 0.02471f $X=11.26 $Y=2.925
+ $X2=0 $Y2=0
cc_416 N_A_1204_107#_c_524_n N_A_938_107#_c_692_n 0.0328866f $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_417 N_A_1204_107#_c_524_n N_A_938_107#_c_731_n 2.78903e-19 $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_418 N_A_1204_107#_c_513_n N_A_938_107#_M1019_g 0.0122632f $X=6.16 $Y=0.745
+ $X2=0 $Y2=0
cc_419 N_A_1204_107#_c_516_n N_A_938_107#_M1019_g 0.00149742f $X=6.325 $Y=0.35
+ $X2=0 $Y2=0
cc_420 N_A_1204_107#_M1029_g N_A_938_107#_M1000_g 0.0244496f $X=10.48 $Y=0.745
+ $X2=0 $Y2=0
cc_421 N_A_1204_107#_c_524_n N_A_938_107#_M1000_g 0.034511f $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_422 N_A_1204_107#_c_525_n N_A_938_107#_c_672_n 0.0103255f $X=7.2 $Y=2.605
+ $X2=0 $Y2=0
cc_423 N_A_1204_107#_c_565_p N_A_938_107#_c_672_n 3.98096e-19 $X=8.21 $Y=1.34
+ $X2=0 $Y2=0
cc_424 N_A_1204_107#_c_535_n N_A_938_107#_c_672_n 0.00167874f $X=7.125 $Y=2.39
+ $X2=0 $Y2=0
cc_425 N_A_1204_107#_c_536_n N_A_938_107#_c_672_n 0.038563f $X=7.142 $Y=2.225
+ $X2=0 $Y2=0
cc_426 N_A_1204_107#_M1021_g N_A_938_107#_c_672_n 0.0432867f $X=7.98 $Y=0.745
+ $X2=0 $Y2=0
cc_427 N_A_1204_107#_c_520_n N_A_1688_81#_M1013_d 0.00248714f $X=10.045 $Y=1.34
+ $X2=0 $Y2=0
cc_428 N_A_1204_107#_c_546_p N_A_1688_81#_c_851_n 0.00403512f $X=8.045 $Y=1.25
+ $X2=14.64 $Y2=0
cc_429 N_A_1204_107#_M1021_g N_A_1688_81#_c_851_n 0.0713016f $X=7.98 $Y=0.745
+ $X2=14.64 $Y2=0
cc_430 N_A_1204_107#_c_520_n N_A_1688_81#_c_853_n 0.0344075f $X=10.045 $Y=1.34
+ $X2=14.64 $Y2=0
cc_431 N_A_1204_107#_c_520_n N_A_1688_81#_c_860_n 0.00332639f $X=10.045 $Y=1.34
+ $X2=0 $Y2=0
cc_432 N_A_1204_107#_M1029_g N_A_1688_81#_c_854_n 0.0109765f $X=10.48 $Y=0.745
+ $X2=0 $Y2=0
cc_433 N_A_1204_107#_M1023_g N_A_1688_81#_c_861_n 6.64786e-19 $X=11.26 $Y=2.925
+ $X2=0 $Y2=0
cc_434 N_A_1204_107#_c_520_n N_A_1688_81#_c_861_n 0.00219243f $X=10.045 $Y=1.34
+ $X2=0 $Y2=0
cc_435 N_A_1204_107#_c_577_p N_A_1688_81#_c_861_n 0.0176411f $X=10.21 $Y=1.61
+ $X2=0 $Y2=0
cc_436 N_A_1204_107#_c_524_n N_A_1688_81#_c_861_n 0.0188235f $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_437 N_A_1204_107#_M1029_g N_A_1688_81#_c_856_n 0.0265449f $X=10.48 $Y=0.745
+ $X2=0 $Y2=0
cc_438 N_A_1204_107#_c_520_n N_A_1688_81#_c_856_n 0.0117287f $X=10.045 $Y=1.34
+ $X2=0 $Y2=0
cc_439 N_A_1204_107#_c_524_n N_A_1688_81#_c_856_n 4.14873e-19 $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_440 N_A_1204_107#_c_520_n N_A_1688_81#_c_879_n 0.0215544f $X=10.045 $Y=1.34
+ $X2=0 $Y2=0
cc_441 N_A_1204_107#_c_524_n N_A_1688_81#_c_879_n 4.85163e-19 $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_442 N_A_1204_107#_M1029_g N_A_1688_81#_c_881_n 0.0136617f $X=10.48 $Y=0.745
+ $X2=0 $Y2=0
cc_443 N_A_1204_107#_c_520_n N_A_1688_81#_c_881_n 0.0122935f $X=10.045 $Y=1.34
+ $X2=0 $Y2=0
cc_444 N_A_1204_107#_c_577_p N_A_1688_81#_c_881_n 0.0233177f $X=10.21 $Y=1.61
+ $X2=0 $Y2=0
cc_445 N_A_1204_107#_c_524_n N_A_1688_81#_c_881_n 0.0227168f $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_446 N_A_1204_107#_c_520_n N_A_1688_81#_c_863_n 0.0063041f $X=10.045 $Y=1.34
+ $X2=0 $Y2=0
cc_447 N_A_1204_107#_c_524_n N_A_1688_81#_c_864_n 3.38342e-19 $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_448 N_A_1204_107#_c_565_p N_A_1490_107#_c_937_n 0.0127038f $X=8.21 $Y=1.34
+ $X2=0 $Y2=0
cc_449 N_A_1204_107#_c_536_n N_A_1490_107#_c_937_n 0.0313952f $X=7.142 $Y=2.225
+ $X2=0 $Y2=0
cc_450 N_A_1204_107#_M1021_g N_A_1490_107#_c_937_n 0.0113799f $X=7.98 $Y=0.745
+ $X2=0 $Y2=0
cc_451 N_A_1204_107#_c_534_n N_A_1490_107#_c_942_n 0.0255453f $X=7.24 $Y=3.335
+ $X2=0.24 $Y2=0
cc_452 N_A_1204_107#_c_520_n N_A_1490_107#_c_938_n 0.100014f $X=10.045 $Y=1.34
+ $X2=14.64 $Y2=0
cc_453 N_A_1204_107#_c_565_p N_A_1490_107#_c_938_n 0.0210413f $X=8.21 $Y=1.34
+ $X2=14.64 $Y2=0
cc_454 N_A_1204_107#_c_577_p N_A_1490_107#_c_938_n 0.00717989f $X=10.21 $Y=1.61
+ $X2=14.64 $Y2=0
cc_455 N_A_1204_107#_M1021_g N_A_1490_107#_c_938_n 0.00554945f $X=7.98 $Y=0.745
+ $X2=14.64 $Y2=0
cc_456 N_A_1204_107#_c_524_n N_A_1490_107#_c_938_n 5.35661e-19 $X=10.48 $Y=1.71
+ $X2=14.64 $Y2=0
cc_457 N_A_1204_107#_c_518_n N_A_1490_107#_c_939_n 0.0199104f $X=7.935 $Y=0.35
+ $X2=7.44 $Y2=0
cc_458 N_A_1204_107#_c_546_p N_A_1490_107#_c_939_n 0.0446926f $X=8.045 $Y=1.25
+ $X2=7.44 $Y2=0
cc_459 N_A_1204_107#_c_536_n N_A_1490_107#_c_939_n 0.0258495f $X=7.142 $Y=2.225
+ $X2=7.44 $Y2=0
cc_460 N_A_1204_107#_M1021_g N_A_1490_107#_c_939_n 0.0067921f $X=7.98 $Y=0.745
+ $X2=7.44 $Y2=0
cc_461 N_A_1204_107#_c_536_n N_A_1490_107#_c_961_n 0.00920714f $X=7.142 $Y=2.225
+ $X2=0 $Y2=0
cc_462 N_A_1204_107#_c_525_n N_A_1490_107#_c_944_n 0.00493617f $X=7.2 $Y=2.605
+ $X2=0 $Y2=0
cc_463 N_A_1204_107#_c_535_n N_A_1490_107#_c_944_n 0.0255453f $X=7.125 $Y=2.39
+ $X2=0 $Y2=0
cc_464 N_A_1204_107#_c_536_n N_A_1490_107#_c_944_n 0.0233784f $X=7.142 $Y=2.225
+ $X2=0 $Y2=0
cc_465 N_A_1204_107#_M1029_g N_A_1490_107#_M1013_g 0.0261111f $X=10.48 $Y=0.745
+ $X2=0 $Y2=0
cc_466 N_A_1204_107#_c_520_n N_A_1490_107#_M1013_g 0.034223f $X=10.045 $Y=1.34
+ $X2=0 $Y2=0
cc_467 N_A_1204_107#_c_577_p N_A_1490_107#_M1013_g 0.00205069f $X=10.21 $Y=1.61
+ $X2=0 $Y2=0
cc_468 N_A_1204_107#_c_524_n N_A_1490_107#_M1013_g 0.0417964f $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_469 N_A_1204_107#_M1023_g N_A_2352_81#_M1004_g 0.043856f $X=11.26 $Y=2.925
+ $X2=0 $Y2=0
cc_470 N_A_1204_107#_c_524_n N_A_2352_81#_c_1022_n 0.043856f $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_471 N_A_1204_107#_M1029_g N_A_2123_543#_c_1107_n 0.0153717f $X=10.48 $Y=0.745
+ $X2=0 $Y2=0
cc_472 N_A_1204_107#_M1023_g N_A_2123_543#_c_1107_n 0.0227378f $X=11.26 $Y=2.925
+ $X2=0 $Y2=0
cc_473 N_A_1204_107#_c_524_n N_A_2123_543#_c_1107_n 0.0282093f $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_474 N_A_1204_107#_M1029_g N_A_2123_543#_c_1110_n 0.00370866f $X=10.48
+ $Y=0.745 $X2=0 $Y2=0
cc_475 N_A_1204_107#_c_524_n N_A_2123_543#_c_1112_n 0.00498566f $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_476 N_A_1204_107#_M1023_g N_A_2123_543#_c_1120_n 0.001351f $X=11.26 $Y=2.925
+ $X2=0 $Y2=0
cc_477 N_A_1204_107#_M1023_g N_A_2123_543#_c_1122_n 0.0165526f $X=11.26 $Y=2.925
+ $X2=0 $Y2=0
cc_478 N_A_1204_107#_c_524_n N_A_2123_543#_c_1122_n 0.00435738f $X=10.48 $Y=1.71
+ $X2=0 $Y2=0
cc_479 N_A_1204_107#_c_527_n N_VPWR_c_1207_n 0.0279815f $X=6.26 $Y=3.11 $X2=0
+ $Y2=0
cc_480 N_A_1204_107#_c_531_n N_VPWR_c_1207_n 0.0252545f $X=6.425 $Y=3.42 $X2=0
+ $Y2=0
cc_481 N_A_1204_107#_M1023_g N_VPWR_c_1213_n 0.00167554f $X=11.26 $Y=2.925 $X2=0
+ $Y2=0
cc_482 N_A_1204_107#_c_525_n N_VPWR_c_1219_n 0.00395199f $X=7.2 $Y=2.605 $X2=0
+ $Y2=0
cc_483 N_A_1204_107#_M1023_g N_VPWR_c_1219_n 0.00191492f $X=11.26 $Y=2.925 $X2=0
+ $Y2=0
cc_484 N_A_1204_107#_c_528_n N_VPWR_c_1219_n 0.0470743f $X=7.155 $Y=3.42 $X2=0
+ $Y2=0
cc_485 N_A_1204_107#_c_531_n N_VPWR_c_1219_n 0.0412003f $X=6.425 $Y=3.42 $X2=0
+ $Y2=0
cc_486 N_A_1204_107#_c_536_n N_A_484_107#_c_1298_n 0.0396884f $X=7.142 $Y=2.225
+ $X2=0 $Y2=0
cc_487 N_A_1204_107#_c_513_n N_A_484_107#_c_1302_n 0.023427f $X=6.16 $Y=0.745
+ $X2=0 $Y2=0
cc_488 N_A_1204_107#_c_514_n N_A_484_107#_c_1302_n 0.0219568f $X=7.075 $Y=0.35
+ $X2=0 $Y2=0
cc_489 N_A_1204_107#_c_536_n N_A_484_107#_c_1302_n 0.0140106f $X=7.142 $Y=2.225
+ $X2=0 $Y2=0
cc_490 N_A_1204_107#_c_536_n N_A_484_107#_c_1309_n 0.00866151f $X=7.142 $Y=2.225
+ $X2=0 $Y2=0
cc_491 N_A_1204_107#_c_525_n N_A_484_107#_c_1310_n 0.0163597f $X=7.2 $Y=2.605
+ $X2=0 $Y2=0
cc_492 N_A_1204_107#_c_527_n N_A_484_107#_c_1310_n 0.0166023f $X=6.26 $Y=3.11
+ $X2=0 $Y2=0
cc_493 N_A_1204_107#_c_528_n N_A_484_107#_c_1310_n 0.0263957f $X=7.155 $Y=3.42
+ $X2=0 $Y2=0
cc_494 N_A_1204_107#_c_534_n N_A_484_107#_c_1310_n 0.0316344f $X=7.24 $Y=3.335
+ $X2=0 $Y2=0
cc_495 N_A_1204_107#_c_535_n N_A_484_107#_c_1310_n 9.56356e-19 $X=7.125 $Y=2.39
+ $X2=0 $Y2=0
cc_496 N_A_1204_107#_c_525_n N_A_484_107#_c_1311_n 0.00899542f $X=7.2 $Y=2.605
+ $X2=0 $Y2=0
cc_497 N_A_1204_107#_c_534_n N_A_484_107#_c_1311_n 0.00707869f $X=7.24 $Y=3.335
+ $X2=0 $Y2=0
cc_498 N_A_1204_107#_c_535_n N_A_484_107#_c_1311_n 0.0210344f $X=7.125 $Y=2.39
+ $X2=0 $Y2=0
cc_499 N_A_1204_107#_c_536_n N_A_484_107#_c_1311_n 0.00963537f $X=7.142 $Y=2.225
+ $X2=0 $Y2=0
cc_500 N_A_1204_107#_c_520_n N_VGND_M1022_d 0.00248253f $X=10.045 $Y=1.34 $X2=0
+ $Y2=0
cc_501 N_A_1204_107#_c_513_n N_VGND_c_1434_n 0.0360977f $X=6.16 $Y=0.745 $X2=0
+ $Y2=0
cc_502 N_A_1204_107#_c_516_n N_VGND_c_1434_n 0.00439711f $X=6.325 $Y=0.35 $X2=0
+ $Y2=0
cc_503 N_A_1204_107#_M1029_g N_VGND_c_1436_n 7.65055e-19 $X=10.48 $Y=0.745 $X2=0
+ $Y2=0
cc_504 N_A_1204_107#_c_518_n N_VGND_c_1436_n 0.0015427f $X=7.935 $Y=0.35 $X2=0
+ $Y2=0
cc_505 N_A_1204_107#_c_546_p N_VGND_c_1436_n 0.0187255f $X=8.045 $Y=1.25 $X2=0
+ $Y2=0
cc_506 N_A_1204_107#_c_520_n N_VGND_c_1436_n 0.0669116f $X=10.045 $Y=1.34 $X2=0
+ $Y2=0
cc_507 N_A_1204_107#_M1021_g N_VGND_c_1436_n 0.00178354f $X=7.98 $Y=0.745 $X2=0
+ $Y2=0
cc_508 N_A_1204_107#_M1029_g N_VGND_c_1442_n 0.0213488f $X=10.48 $Y=0.745 $X2=0
+ $Y2=0
cc_509 N_A_1204_107#_c_513_n N_VGND_c_1442_n 0.0320609f $X=6.16 $Y=0.745 $X2=0
+ $Y2=0
cc_510 N_A_1204_107#_c_514_n N_VGND_c_1442_n 0.0292874f $X=7.075 $Y=0.35 $X2=0
+ $Y2=0
cc_511 N_A_1204_107#_c_516_n N_VGND_c_1442_n 0.0111249f $X=6.325 $Y=0.35 $X2=0
+ $Y2=0
cc_512 N_A_1204_107#_c_518_n N_VGND_c_1442_n 0.0345591f $X=7.935 $Y=0.35 $X2=0
+ $Y2=0
cc_513 N_A_1204_107#_c_546_p N_VGND_c_1442_n 0.0302286f $X=8.045 $Y=1.25 $X2=0
+ $Y2=0
cc_514 N_A_1204_107#_c_536_n N_VGND_c_1442_n 0.0229942f $X=7.142 $Y=2.225 $X2=0
+ $Y2=0
cc_515 N_A_1204_107#_c_521_n N_VGND_c_1442_n 0.00355762f $X=7.16 $Y=0.35 $X2=0
+ $Y2=0
cc_516 N_A_1204_107#_M1021_g N_VGND_c_1442_n 0.0112989f $X=7.98 $Y=0.745 $X2=0
+ $Y2=0
cc_517 N_A_938_107#_c_684_n N_A_1688_81#_M1017_d 0.00397455f $X=10.32 $Y=3.24
+ $X2=0 $Y2=0
cc_518 N_A_938_107#_M1024_g N_A_1688_81#_M1026_g 0.0492803f $X=7.98 $Y=2.925
+ $X2=0 $Y2=0
cc_519 N_A_938_107#_c_684_n N_A_1688_81#_M1026_g 0.0321434f $X=10.32 $Y=3.24
+ $X2=0 $Y2=0
cc_520 N_A_938_107#_c_744_p N_A_1688_81#_M1026_g 0.00337089f $X=8.045 $Y=2.495
+ $X2=0 $Y2=0
cc_521 N_A_938_107#_c_692_n N_A_1688_81#_c_861_n 0.00704942f $X=10.325 $Y=2.39
+ $X2=0 $Y2=0
cc_522 N_A_938_107#_c_731_n N_A_1688_81#_c_861_n 0.0228878f $X=10.405 $Y=2.4
+ $X2=0 $Y2=0
cc_523 N_A_938_107#_M1000_g N_A_1688_81#_c_881_n 2.87685e-19 $X=11.3 $Y=0.745
+ $X2=0 $Y2=0
cc_524 N_A_938_107#_c_748_p N_A_1688_81#_c_894_n 0.0223329f $X=8.045 $Y=2.05
+ $X2=0 $Y2=0
cc_525 N_A_938_107#_c_684_n N_A_1688_81#_c_894_n 0.00871826f $X=10.32 $Y=3.24
+ $X2=0 $Y2=0
cc_526 N_A_938_107#_c_672_n N_A_1688_81#_c_894_n 0.00175039f $X=7.98 $Y=1.725
+ $X2=0 $Y2=0
cc_527 N_A_938_107#_c_748_p N_A_1688_81#_c_857_n 0.00337089f $X=8.045 $Y=2.05
+ $X2=0 $Y2=0
cc_528 N_A_938_107#_c_684_n N_A_1688_81#_c_857_n 7.47771e-19 $X=10.32 $Y=3.24
+ $X2=0 $Y2=0
cc_529 N_A_938_107#_c_672_n N_A_1688_81#_c_857_n 0.0492803f $X=7.98 $Y=1.725
+ $X2=0 $Y2=0
cc_530 N_A_938_107#_c_684_n N_A_1688_81#_c_864_n 0.0150973f $X=10.32 $Y=3.24
+ $X2=0 $Y2=0
cc_531 N_A_938_107#_c_725_n N_A_1688_81#_c_864_n 0.020464f $X=10.405 $Y=3.155
+ $X2=0 $Y2=0
cc_532 N_A_938_107#_c_692_n N_A_1688_81#_c_864_n 0.00631361f $X=10.325 $Y=2.39
+ $X2=0 $Y2=0
cc_533 N_A_938_107#_c_725_n N_A_1688_81#_c_865_n 0.00765971f $X=10.405 $Y=3.155
+ $X2=0 $Y2=0
cc_534 N_A_938_107#_c_692_n N_A_1688_81#_c_865_n 0.005298f $X=10.325 $Y=2.39
+ $X2=0 $Y2=0
cc_535 N_A_938_107#_c_731_n N_A_1688_81#_c_865_n 0.013596f $X=10.405 $Y=2.4
+ $X2=0 $Y2=0
cc_536 N_A_938_107#_c_672_n N_A_1688_81#_c_858_n 0.0133713f $X=7.98 $Y=1.725
+ $X2=0 $Y2=0
cc_537 N_A_938_107#_M1028_g N_A_1490_107#_c_937_n 0.00278707f $X=7.2 $Y=0.745
+ $X2=0 $Y2=0
cc_538 N_A_938_107#_c_672_n N_A_1490_107#_c_937_n 0.0111989f $X=7.98 $Y=1.725
+ $X2=0 $Y2=0
cc_539 N_A_938_107#_M1024_g N_A_1490_107#_c_942_n 0.00420344f $X=7.98 $Y=2.925
+ $X2=0.24 $Y2=0
cc_540 N_A_938_107#_c_764_p N_A_1490_107#_c_942_n 0.0221386f $X=8.125 $Y=3.155
+ $X2=0.24 $Y2=0
cc_541 N_A_938_107#_c_672_n N_A_1490_107#_c_942_n 0.00166031f $X=7.98 $Y=1.725
+ $X2=0.24 $Y2=0
cc_542 N_A_938_107#_M1024_g N_A_1490_107#_c_943_n 0.00835881f $X=7.98 $Y=2.925
+ $X2=0 $Y2=0
cc_543 N_A_938_107#_c_686_n N_A_1490_107#_c_943_n 0.00103361f $X=8.21 $Y=3.24
+ $X2=0 $Y2=0
cc_544 N_A_938_107#_c_748_p N_A_1490_107#_c_938_n 0.0236391f $X=8.045 $Y=2.05
+ $X2=14.64 $Y2=0
cc_545 N_A_938_107#_c_672_n N_A_1490_107#_c_938_n 0.0193388f $X=7.98 $Y=1.725
+ $X2=14.64 $Y2=0
cc_546 N_A_938_107#_M1028_g N_A_1490_107#_c_939_n 0.00808788f $X=7.2 $Y=0.745
+ $X2=7.44 $Y2=0
cc_547 N_A_938_107#_c_672_n N_A_1490_107#_c_939_n 0.00220512f $X=7.98 $Y=1.725
+ $X2=7.44 $Y2=0
cc_548 N_A_938_107#_c_672_n N_A_1490_107#_c_961_n 0.0165579f $X=7.98 $Y=1.725
+ $X2=0 $Y2=0
cc_549 N_A_938_107#_M1024_g N_A_1490_107#_c_944_n 0.00542254f $X=7.98 $Y=2.925
+ $X2=0 $Y2=0
cc_550 N_A_938_107#_c_748_p N_A_1490_107#_c_944_n 0.0349414f $X=8.045 $Y=2.05
+ $X2=0 $Y2=0
cc_551 N_A_938_107#_c_764_p N_A_1490_107#_c_944_n 0.00724041f $X=8.125 $Y=3.155
+ $X2=0 $Y2=0
cc_552 N_A_938_107#_c_672_n N_A_1490_107#_c_944_n 0.0253395f $X=7.98 $Y=1.725
+ $X2=0 $Y2=0
cc_553 N_A_938_107#_c_684_n N_A_1490_107#_M1013_g 0.0411689f $X=10.32 $Y=3.24
+ $X2=0 $Y2=0
cc_554 N_A_938_107#_c_725_n N_A_1490_107#_M1013_g 9.00746e-19 $X=10.405 $Y=3.155
+ $X2=0 $Y2=0
cc_555 N_A_938_107#_c_692_n N_A_1490_107#_M1013_g 0.0626456f $X=10.325 $Y=2.39
+ $X2=0 $Y2=0
cc_556 N_A_938_107#_c_695_n N_A_1490_107#_M1013_g 9.72755e-19 $X=10.405 $Y=3.24
+ $X2=0 $Y2=0
cc_557 N_A_938_107#_c_665_n N_A_2352_81#_M1001_g 0.00136124f $X=11.355 $Y=1.25
+ $X2=0 $Y2=0
cc_558 N_A_938_107#_M1000_g N_A_2352_81#_M1001_g 0.0667482f $X=11.3 $Y=0.745
+ $X2=0 $Y2=0
cc_559 N_A_938_107#_c_665_n N_A_2352_81#_M1004_g 0.00347593f $X=11.355 $Y=1.25
+ $X2=0 $Y2=0
cc_560 N_A_938_107#_c_665_n N_A_2352_81#_c_1022_n 7.99646e-19 $X=11.355 $Y=1.25
+ $X2=0 $Y2=0
cc_561 N_A_938_107#_c_688_n N_A_2123_543#_M1031_d 0.00600953f $X=11.255 $Y=3.41
+ $X2=0 $Y2=0
cc_562 N_A_938_107#_c_725_n N_A_2123_543#_c_1107_n 0.00802745f $X=10.405
+ $Y=3.155 $X2=0 $Y2=0
cc_563 N_A_938_107#_c_665_n N_A_2123_543#_c_1107_n 0.108766f $X=11.355 $Y=1.25
+ $X2=0 $Y2=0
cc_564 N_A_938_107#_c_692_n N_A_2123_543#_c_1107_n 0.00594042f $X=10.325 $Y=2.39
+ $X2=0 $Y2=0
cc_565 N_A_938_107#_c_731_n N_A_2123_543#_c_1107_n 0.00880421f $X=10.405 $Y=2.4
+ $X2=0 $Y2=0
cc_566 N_A_938_107#_M1000_g N_A_2123_543#_c_1107_n 0.021061f $X=11.3 $Y=0.745
+ $X2=0 $Y2=0
cc_567 N_A_938_107#_c_665_n N_A_2123_543#_c_1108_n 0.00565817f $X=11.355 $Y=1.25
+ $X2=0 $Y2=0
cc_568 N_A_938_107#_M1000_g N_A_2123_543#_c_1108_n 0.0295284f $X=11.3 $Y=0.745
+ $X2=0 $Y2=0
cc_569 N_A_938_107#_M1000_g N_A_2123_543#_c_1110_n 0.00113377f $X=11.3 $Y=0.745
+ $X2=0 $Y2=0
cc_570 N_A_938_107#_c_665_n N_A_2123_543#_c_1112_n 0.0879404f $X=11.355 $Y=1.25
+ $X2=0 $Y2=0
cc_571 N_A_938_107#_M1000_g N_A_2123_543#_c_1112_n 0.00715659f $X=11.3 $Y=0.745
+ $X2=0 $Y2=0
cc_572 N_A_938_107#_c_665_n N_A_2123_543#_c_1120_n 0.0132568f $X=11.355 $Y=1.25
+ $X2=0 $Y2=0
cc_573 N_A_938_107#_c_725_n N_A_2123_543#_c_1122_n 0.0167913f $X=10.405 $Y=3.155
+ $X2=0 $Y2=0
cc_574 N_A_938_107#_c_688_n N_A_2123_543#_c_1122_n 0.0280676f $X=11.255 $Y=3.41
+ $X2=0 $Y2=0
cc_575 N_A_938_107#_c_665_n N_A_2123_543#_c_1122_n 0.0329407f $X=11.355 $Y=1.25
+ $X2=0 $Y2=0
cc_576 N_A_938_107#_c_692_n N_A_2123_543#_c_1122_n 7.17414e-19 $X=10.325 $Y=2.39
+ $X2=0 $Y2=0
cc_577 N_A_938_107#_c_684_n N_VPWR_M1026_d 0.011249f $X=10.32 $Y=3.24 $X2=0
+ $Y2=0
cc_578 N_A_938_107#_c_679_n N_VPWR_c_1204_n 0.0557548f $X=4.93 $Y=3.11 $X2=0
+ $Y2=0
cc_579 N_A_938_107#_c_659_n N_VPWR_c_1207_n 0.00928005f $X=5.87 $Y=2.835 $X2=0
+ $Y2=0
cc_580 N_A_938_107#_M1020_g N_VPWR_c_1207_n 0.0496358f $X=5.87 $Y=3.34 $X2=0
+ $Y2=0
cc_581 N_A_938_107#_c_679_n N_VPWR_c_1207_n 0.0527223f $X=4.93 $Y=3.11 $X2=0
+ $Y2=0
cc_582 N_A_938_107#_c_682_n N_VPWR_c_1207_n 0.0242975f $X=5.275 $Y=2.68 $X2=0
+ $Y2=0
cc_583 N_A_938_107#_c_684_n N_VPWR_c_1210_n 0.0498453f $X=10.32 $Y=3.24 $X2=0
+ $Y2=0
cc_584 N_A_938_107#_c_692_n N_VPWR_c_1210_n 0.00515298f $X=10.325 $Y=2.39 $X2=0
+ $Y2=0
cc_585 N_A_938_107#_c_688_n N_VPWR_c_1213_n 0.00615971f $X=11.255 $Y=3.41 $X2=0
+ $Y2=0
cc_586 N_A_938_107#_c_665_n N_VPWR_c_1213_n 0.019488f $X=11.355 $Y=1.25 $X2=0
+ $Y2=0
cc_587 N_A_938_107#_c_659_n N_VPWR_c_1219_n 0.00148679f $X=5.87 $Y=2.835 $X2=0
+ $Y2=0
cc_588 N_A_938_107#_M1020_g N_VPWR_c_1219_n 0.0124253f $X=5.87 $Y=3.34 $X2=0
+ $Y2=0
cc_589 N_A_938_107#_M1024_g N_VPWR_c_1219_n 0.00973252f $X=7.98 $Y=2.925 $X2=0
+ $Y2=0
cc_590 N_A_938_107#_c_679_n N_VPWR_c_1219_n 0.0382178f $X=4.93 $Y=3.11 $X2=0
+ $Y2=0
cc_591 N_A_938_107#_c_684_n N_VPWR_c_1219_n 0.0714868f $X=10.32 $Y=3.24 $X2=0
+ $Y2=0
cc_592 N_A_938_107#_c_686_n N_VPWR_c_1219_n 0.0071121f $X=8.21 $Y=3.24 $X2=0
+ $Y2=0
cc_593 N_A_938_107#_c_688_n N_VPWR_c_1219_n 0.0477764f $X=11.255 $Y=3.41 $X2=0
+ $Y2=0
cc_594 N_A_938_107#_c_692_n N_VPWR_c_1219_n 0.0163929f $X=10.325 $Y=2.39 $X2=0
+ $Y2=0
cc_595 N_A_938_107#_c_695_n N_VPWR_c_1219_n 0.0148841f $X=10.405 $Y=3.24 $X2=0
+ $Y2=0
cc_596 N_A_938_107#_c_659_n N_A_484_107#_c_1297_n 0.0598536f $X=5.87 $Y=2.835
+ $X2=7.44 $Y2=0
cc_597 N_A_938_107#_c_660_n N_A_484_107#_c_1297_n 0.0306974f $X=6.95 $Y=1.635
+ $X2=7.44 $Y2=0
cc_598 N_A_938_107#_c_663_n N_A_484_107#_c_1297_n 0.0172997f $X=5.54 $Y=1.24
+ $X2=7.44 $Y2=0
cc_599 N_A_938_107#_c_664_n N_A_484_107#_c_1297_n 0.00642736f $X=5.025 $Y=1.24
+ $X2=7.44 $Y2=0
cc_600 N_A_938_107#_c_682_n N_A_484_107#_c_1297_n 0.00581989f $X=5.275 $Y=2.68
+ $X2=7.44 $Y2=0
cc_601 N_A_938_107#_c_683_n N_A_484_107#_c_1297_n 0.0119473f $X=5.095 $Y=2.68
+ $X2=7.44 $Y2=0
cc_602 N_A_938_107#_c_706_n N_A_484_107#_c_1297_n 0.0246744f $X=5.44 $Y=2.3
+ $X2=7.44 $Y2=0
cc_603 N_A_938_107#_c_827_p N_A_484_107#_c_1297_n 0.0236659f $X=5.705 $Y=1.25
+ $X2=7.44 $Y2=0
cc_604 N_A_938_107#_c_660_n N_A_484_107#_c_1298_n 0.0545879f $X=6.95 $Y=1.635
+ $X2=0 $Y2=0
cc_605 N_A_938_107#_M1028_g N_A_484_107#_c_1298_n 0.00726813f $X=7.2 $Y=0.745
+ $X2=0 $Y2=0
cc_606 N_A_938_107#_c_660_n N_A_484_107#_c_1302_n 0.00320745f $X=6.95 $Y=1.635
+ $X2=0 $Y2=0
cc_607 N_A_938_107#_M1028_g N_A_484_107#_c_1302_n 0.00966503f $X=7.2 $Y=0.745
+ $X2=0 $Y2=0
cc_608 N_A_938_107#_M1019_g N_A_484_107#_c_1302_n 0.00892551f $X=5.77 $Y=0.745
+ $X2=0 $Y2=0
cc_609 N_A_938_107#_c_660_n N_A_484_107#_c_1309_n 0.0101148f $X=6.95 $Y=1.635
+ $X2=0 $Y2=0
cc_610 N_A_938_107#_M1020_g N_A_484_107#_c_1310_n 0.011734f $X=5.87 $Y=3.34
+ $X2=0 $Y2=0
cc_611 N_A_938_107#_c_660_n N_A_484_107#_c_1310_n 0.00100244f $X=6.95 $Y=1.635
+ $X2=0 $Y2=0
cc_612 N_A_938_107#_c_659_n N_A_484_107#_c_1311_n 0.0113593f $X=5.87 $Y=2.835
+ $X2=0 $Y2=0
cc_613 N_A_938_107#_c_662_n N_VGND_c_1432_n 8.65424e-19 $X=4.94 $Y=1.155 $X2=0
+ $Y2=0
cc_614 N_A_938_107#_c_666_n N_VGND_c_1432_n 0.0334873f $X=4.83 $Y=0.745 $X2=0
+ $Y2=0
cc_615 N_A_938_107#_c_663_n N_VGND_c_1434_n 0.0249965f $X=5.54 $Y=1.24 $X2=0
+ $Y2=0
cc_616 N_A_938_107#_c_666_n N_VGND_c_1434_n 0.0355362f $X=4.83 $Y=0.745 $X2=0
+ $Y2=0
cc_617 N_A_938_107#_c_827_p N_VGND_c_1434_n 0.0200253f $X=5.705 $Y=1.25 $X2=0
+ $Y2=0
cc_618 N_A_938_107#_M1019_g N_VGND_c_1434_n 0.0344571f $X=5.77 $Y=0.745 $X2=0
+ $Y2=0
cc_619 N_A_938_107#_M1000_g N_VGND_c_1438_n 0.00102038f $X=11.3 $Y=0.745 $X2=0
+ $Y2=0
cc_620 N_A_938_107#_M1028_g N_VGND_c_1442_n 0.0178578f $X=7.2 $Y=0.745 $X2=0
+ $Y2=0
cc_621 N_A_938_107#_c_663_n N_VGND_c_1442_n 0.00794827f $X=5.54 $Y=1.24 $X2=0
+ $Y2=0
cc_622 N_A_938_107#_c_665_n N_VGND_c_1442_n 0.00127079f $X=11.355 $Y=1.25 $X2=0
+ $Y2=0
cc_623 N_A_938_107#_c_666_n N_VGND_c_1442_n 0.0291907f $X=4.83 $Y=0.745 $X2=0
+ $Y2=0
cc_624 N_A_938_107#_c_827_p N_VGND_c_1442_n 0.00309009f $X=5.705 $Y=1.25 $X2=0
+ $Y2=0
cc_625 N_A_938_107#_M1019_g N_VGND_c_1442_n 0.00867625f $X=5.77 $Y=0.745 $X2=0
+ $Y2=0
cc_626 N_A_938_107#_M1000_g N_VGND_c_1442_n 0.0063847f $X=11.3 $Y=0.745 $X2=0
+ $Y2=0
cc_627 N_A_1688_81#_c_853_n N_A_1490_107#_c_937_n 0.00326231f $X=8.705 $Y=1.565
+ $X2=0 $Y2=0
cc_628 N_A_1688_81#_c_853_n N_A_1490_107#_c_938_n 2.88561e-19 $X=8.705 $Y=1.565
+ $X2=14.64 $Y2=0
cc_629 N_A_1688_81#_c_860_n N_A_1490_107#_c_938_n 0.0503224f $X=9.81 $Y=2.04
+ $X2=14.64 $Y2=0
cc_630 N_A_1688_81#_c_894_n N_A_1490_107#_c_938_n 0.0237561f $X=8.785 $Y=2.05
+ $X2=14.64 $Y2=0
cc_631 N_A_1688_81#_c_857_n N_A_1490_107#_c_938_n 7.46081e-19 $X=8.785 $Y=2.05
+ $X2=14.64 $Y2=0
cc_632 N_A_1688_81#_c_858_n N_A_1490_107#_c_938_n 0.0313261f $X=8.705 $Y=1.865
+ $X2=14.64 $Y2=0
cc_633 N_A_1688_81#_M1026_g N_A_1490_107#_M1013_g 0.0285736f $X=8.69 $Y=2.925
+ $X2=0 $Y2=0
cc_634 N_A_1688_81#_c_851_n N_A_1490_107#_M1013_g 0.0132547f $X=8.705 $Y=1.065
+ $X2=0 $Y2=0
cc_635 N_A_1688_81#_c_853_n N_A_1490_107#_M1013_g 0.0617038f $X=8.705 $Y=1.565
+ $X2=0 $Y2=0
cc_636 N_A_1688_81#_c_860_n N_A_1490_107#_M1013_g 0.0390248f $X=9.81 $Y=2.04
+ $X2=0 $Y2=0
cc_637 N_A_1688_81#_c_854_n N_A_1490_107#_M1013_g 0.00791276f $X=9.975 $Y=0.905
+ $X2=0 $Y2=0
cc_638 N_A_1688_81#_c_879_n N_A_1490_107#_M1013_g 0.00413441f $X=10.14 $Y=0.99
+ $X2=0 $Y2=0
cc_639 N_A_1688_81#_c_881_n N_A_1490_107#_M1013_g 0.00154662f $X=10.56 $Y=1.955
+ $X2=0 $Y2=0
cc_640 N_A_1688_81#_c_894_n N_A_1490_107#_M1013_g 0.00281989f $X=8.785 $Y=2.05
+ $X2=0 $Y2=0
cc_641 N_A_1688_81#_c_863_n N_A_1490_107#_M1013_g 0.00468122f $X=9.895 $Y=2.04
+ $X2=0 $Y2=0
cc_642 N_A_1688_81#_c_864_n N_A_1490_107#_M1013_g 0.0148952f $X=9.975 $Y=2.865
+ $X2=0 $Y2=0
cc_643 N_A_1688_81#_c_865_n N_A_1490_107#_M1013_g 0.0287908f $X=9.975 $Y=2.675
+ $X2=0 $Y2=0
cc_644 N_A_1688_81#_c_861_n N_A_2123_543#_c_1107_n 0.0138169f $X=10.475 $Y=2.04
+ $X2=0 $Y2=0
cc_645 N_A_1688_81#_c_856_n N_A_2123_543#_c_1107_n 0.0133059f $X=10.475 $Y=0.99
+ $X2=0 $Y2=0
cc_646 N_A_1688_81#_c_881_n N_A_2123_543#_c_1107_n 0.0608791f $X=10.56 $Y=1.955
+ $X2=0 $Y2=0
cc_647 N_A_1688_81#_M1017_d N_VPWR_c_1210_n 0.00401999f $X=9.835 $Y=2.715 $X2=0
+ $Y2=0
cc_648 N_A_1688_81#_M1017_d N_VPWR_c_1219_n 0.00231205f $X=9.835 $Y=2.715 $X2=0
+ $Y2=0
cc_649 N_A_1688_81#_c_851_n N_VGND_c_1436_n 0.0401918f $X=8.705 $Y=1.065 $X2=0
+ $Y2=0
cc_650 N_A_1688_81#_c_853_n N_VGND_c_1436_n 0.00562274f $X=8.705 $Y=1.565 $X2=0
+ $Y2=0
cc_651 N_A_1688_81#_c_854_n N_VGND_c_1436_n 0.029197f $X=9.975 $Y=0.905 $X2=0
+ $Y2=0
cc_652 N_A_1688_81#_c_879_n N_VGND_c_1436_n 0.0136768f $X=10.14 $Y=0.99 $X2=0
+ $Y2=0
cc_653 N_A_1688_81#_M1013_d N_VGND_c_1442_n 8.87201e-19 $X=9.835 $Y=0.535 $X2=0
+ $Y2=0
cc_654 N_A_1688_81#_c_851_n N_VGND_c_1442_n 0.0158717f $X=8.705 $Y=1.065 $X2=0
+ $Y2=0
cc_655 N_A_1688_81#_c_854_n N_VGND_c_1442_n 0.0324043f $X=9.975 $Y=0.905 $X2=0
+ $Y2=0
cc_656 N_A_1688_81#_c_856_n N_VGND_c_1442_n 0.0205294f $X=10.475 $Y=0.99 $X2=0
+ $Y2=0
cc_657 N_A_1490_107#_M1013_g N_VPWR_c_1210_n 0.0205123f $X=9.585 $Y=0.91 $X2=0
+ $Y2=0
cc_658 N_A_1490_107#_c_943_n N_VPWR_c_1219_n 0.0126529f $X=7.59 $Y=2.925 $X2=0
+ $Y2=0
cc_659 N_A_1490_107#_M1013_g N_VPWR_c_1219_n 0.00761806f $X=9.585 $Y=0.91 $X2=0
+ $Y2=0
cc_660 N_A_1490_107#_M1013_g N_VGND_c_1436_n 0.0409369f $X=9.585 $Y=0.91 $X2=0
+ $Y2=0
cc_661 N_A_1490_107#_c_939_n N_VGND_c_1442_n 0.0222434f $X=7.59 $Y=0.765 $X2=0
+ $Y2=0
cc_662 N_A_1490_107#_M1013_g N_VGND_c_1442_n 0.0111156f $X=9.585 $Y=0.91 $X2=0
+ $Y2=0
cc_663 N_A_2352_81#_M1001_g N_A_2123_543#_M1002_g 0.0247098f $X=12.01 $Y=0.745
+ $X2=0 $Y2=0
cc_664 N_A_2352_81#_c_1016_n N_A_2123_543#_M1002_g 0.0372017f $X=13.965 $Y=1.8
+ $X2=0 $Y2=0
cc_665 N_A_2352_81#_c_1018_n N_A_2123_543#_M1002_g 0.0339489f $X=13.11 $Y=1.57
+ $X2=0 $Y2=0
cc_666 N_A_2352_81#_c_1019_n N_A_2123_543#_M1002_g 0.0268945f $X=13.275 $Y=0.68
+ $X2=0 $Y2=0
cc_667 N_A_2352_81#_c_1021_n N_A_2123_543#_M1002_g 0.0121786f $X=13.275 $Y=2.015
+ $X2=0 $Y2=0
cc_668 N_A_2352_81#_c_1044_p N_A_2123_543#_M1002_g 0.00114094f $X=12.145 $Y=1.65
+ $X2=0 $Y2=0
cc_669 N_A_2352_81#_c_1022_n N_A_2123_543#_M1002_g 0.0165182f $X=12.145 $Y=1.65
+ $X2=0 $Y2=0
cc_670 N_A_2352_81#_M1004_g N_A_2123_543#_M1005_g 0.0142089f $X=12.01 $Y=2.925
+ $X2=0 $Y2=0
cc_671 N_A_2352_81#_c_1029_n N_A_2123_543#_M1005_g 0.0236877f $X=13.275 $Y=2.86
+ $X2=0 $Y2=0
cc_672 N_A_2352_81#_M1001_g N_A_2123_543#_c_1107_n 3.08458e-19 $X=12.01 $Y=0.745
+ $X2=0 $Y2=0
cc_673 N_A_2352_81#_M1001_g N_A_2123_543#_c_1108_n 0.00413314f $X=12.01 $Y=0.745
+ $X2=0 $Y2=0
cc_674 N_A_2352_81#_M1001_g N_A_2123_543#_c_1112_n 0.0229666f $X=12.01 $Y=0.745
+ $X2=0 $Y2=0
cc_675 N_A_2352_81#_M1004_g N_A_2123_543#_c_1112_n 0.00861921f $X=12.01 $Y=2.925
+ $X2=0 $Y2=0
cc_676 N_A_2352_81#_c_1044_p N_A_2123_543#_c_1112_n 0.046437f $X=12.145 $Y=1.65
+ $X2=0 $Y2=0
cc_677 N_A_2352_81#_c_1022_n N_A_2123_543#_c_1112_n 0.0200086f $X=12.145 $Y=1.65
+ $X2=0 $Y2=0
cc_678 N_A_2352_81#_M1004_g N_A_2123_543#_c_1119_n 0.0333672f $X=12.01 $Y=2.925
+ $X2=7.44 $Y2=0.057
cc_679 N_A_2352_81#_c_1029_n N_A_2123_543#_c_1119_n 0.0129587f $X=13.275 $Y=2.86
+ $X2=7.44 $Y2=0.057
cc_680 N_A_2352_81#_c_1044_p N_A_2123_543#_c_1119_n 0.0230012f $X=12.145 $Y=1.65
+ $X2=7.44 $Y2=0.057
cc_681 N_A_2352_81#_c_1022_n N_A_2123_543#_c_1119_n 0.00216891f $X=12.145
+ $Y=1.65 $X2=7.44 $Y2=0.057
cc_682 N_A_2352_81#_M1004_g N_A_2123_543#_c_1120_n 0.0037179f $X=12.01 $Y=2.925
+ $X2=0 $Y2=0
cc_683 N_A_2352_81#_M1004_g N_A_2123_543#_c_1170_n 0.00113312f $X=12.01 $Y=2.925
+ $X2=0 $Y2=0
cc_684 N_A_2352_81#_c_1018_n N_A_2123_543#_c_1170_n 0.0229442f $X=13.11 $Y=1.57
+ $X2=0 $Y2=0
cc_685 N_A_2352_81#_c_1021_n N_A_2123_543#_c_1170_n 0.0127596f $X=13.275
+ $Y=2.015 $X2=0 $Y2=0
cc_686 N_A_2352_81#_c_1029_n N_A_2123_543#_c_1170_n 0.0235836f $X=13.275 $Y=2.86
+ $X2=0 $Y2=0
cc_687 N_A_2352_81#_c_1044_p N_A_2123_543#_c_1170_n 0.0151792f $X=12.145 $Y=1.65
+ $X2=0 $Y2=0
cc_688 N_A_2352_81#_c_1022_n N_A_2123_543#_c_1170_n 0.00140038f $X=12.145
+ $Y=1.65 $X2=0 $Y2=0
cc_689 N_A_2352_81#_M1004_g N_A_2123_543#_c_1113_n 0.0183386f $X=12.01 $Y=2.925
+ $X2=0 $Y2=0
cc_690 N_A_2352_81#_c_1018_n N_A_2123_543#_c_1113_n 0.00177552f $X=13.11 $Y=1.57
+ $X2=0 $Y2=0
cc_691 N_A_2352_81#_c_1021_n N_A_2123_543#_c_1113_n 0.0056611f $X=13.275
+ $Y=2.015 $X2=0 $Y2=0
cc_692 N_A_2352_81#_c_1029_n N_A_2123_543#_c_1113_n 0.0223802f $X=13.275 $Y=2.86
+ $X2=0 $Y2=0
cc_693 N_A_2352_81#_c_1044_p N_A_2123_543#_c_1113_n 0.00139362f $X=12.145
+ $Y=1.65 $X2=0 $Y2=0
cc_694 N_A_2352_81#_c_1022_n N_A_2123_543#_c_1113_n 0.0191432f $X=12.145 $Y=1.65
+ $X2=0 $Y2=0
cc_695 N_A_2352_81#_M1004_g N_VPWR_c_1213_n 0.0437985f $X=12.01 $Y=2.925 $X2=0
+ $Y2=0
cc_696 N_A_2352_81#_c_1029_n N_VPWR_c_1213_n 0.0747268f $X=13.275 $Y=2.86 $X2=0
+ $Y2=0
cc_697 N_A_2352_81#_M1010_g N_VPWR_c_1216_n 0.0683883f $X=14.215 $Y=2.965 $X2=0
+ $Y2=0
cc_698 N_A_2352_81#_M1004_g N_VPWR_c_1219_n 0.00692603f $X=12.01 $Y=2.925 $X2=0
+ $Y2=0
cc_699 N_A_2352_81#_M1010_g N_VPWR_c_1219_n 0.0117682f $X=14.215 $Y=2.965 $X2=0
+ $Y2=0
cc_700 N_A_2352_81#_c_1029_n N_VPWR_c_1219_n 0.0382178f $X=13.275 $Y=2.86 $X2=0
+ $Y2=0
cc_701 N_A_2352_81#_M1012_g N_Q_c_1392_n 0.0161679f $X=14.215 $Y=1.01 $X2=0
+ $Y2=0
cc_702 N_A_2352_81#_c_1019_n N_Q_c_1392_n 0.049515f $X=13.275 $Y=0.68 $X2=0
+ $Y2=0
cc_703 N_A_2352_81#_M1010_g N_Q_c_1396_n 0.026167f $X=14.215 $Y=2.965 $X2=0
+ $Y2=0
cc_704 N_A_2352_81#_M1012_g N_Q_c_1394_n 0.0116277f $X=14.215 $Y=1.01 $X2=0
+ $Y2=0
cc_705 N_A_2352_81#_c_1016_n N_Q_c_1394_n 0.0215371f $X=13.965 $Y=1.8 $X2=0
+ $Y2=0
cc_706 N_A_2352_81#_c_1017_n N_Q_c_1394_n 0.00137245f $X=14.215 $Y=1.8 $X2=0
+ $Y2=0
cc_707 N_A_2352_81#_c_1019_n N_Q_c_1394_n 0.0112031f $X=13.275 $Y=0.68 $X2=0
+ $Y2=0
cc_708 N_A_2352_81#_c_1021_n N_Q_c_1394_n 0.0173465f $X=13.275 $Y=2.015 $X2=0
+ $Y2=0
cc_709 N_A_2352_81#_M1010_g N_Q_c_1399_n 0.00390564f $X=14.215 $Y=2.965 $X2=0
+ $Y2=0
cc_710 N_A_2352_81#_c_1016_n N_Q_c_1399_n 0.00930741f $X=13.965 $Y=1.8 $X2=0
+ $Y2=0
cc_711 N_A_2352_81#_c_1021_n N_Q_c_1399_n 7.30295e-19 $X=13.275 $Y=2.015 $X2=0
+ $Y2=0
cc_712 N_A_2352_81#_c_1029_n N_Q_c_1399_n 0.103686f $X=13.275 $Y=2.86 $X2=0
+ $Y2=0
cc_713 N_A_2352_81#_M1010_g N_Q_c_1400_n 0.00680362f $X=14.215 $Y=2.965 $X2=7.44
+ $Y2=0
cc_714 N_A_2352_81#_c_1016_n N_Q_c_1400_n 0.0109f $X=13.965 $Y=1.8 $X2=7.44
+ $Y2=0
cc_715 N_A_2352_81#_c_1017_n N_Q_c_1400_n 0.0141147f $X=14.215 $Y=1.8 $X2=7.44
+ $Y2=0
cc_716 N_A_2352_81#_c_1021_n N_Q_c_1400_n 0.0167868f $X=13.275 $Y=2.015 $X2=7.44
+ $Y2=0
cc_717 N_A_2352_81#_c_1029_n N_Q_c_1400_n 0.00716551f $X=13.275 $Y=2.86 $X2=7.44
+ $Y2=0
cc_718 N_A_2352_81#_M1012_g Q 0.0127006f $X=14.215 $Y=1.01 $X2=7.44 $Y2=0.057
cc_719 N_A_2352_81#_c_1017_n Q 0.0307464f $X=14.215 $Y=1.8 $X2=7.44 $Y2=0.057
cc_720 N_A_2352_81#_M1001_g N_VGND_c_1438_n 0.0577821f $X=12.01 $Y=0.745 $X2=0
+ $Y2=0
cc_721 N_A_2352_81#_c_1018_n N_VGND_c_1438_n 0.0476367f $X=13.11 $Y=1.57 $X2=0
+ $Y2=0
cc_722 N_A_2352_81#_c_1019_n N_VGND_c_1438_n 0.0583597f $X=13.275 $Y=0.68 $X2=0
+ $Y2=0
cc_723 N_A_2352_81#_c_1044_p N_VGND_c_1438_n 0.0267852f $X=12.145 $Y=1.65 $X2=0
+ $Y2=0
cc_724 N_A_2352_81#_c_1022_n N_VGND_c_1438_n 0.00193505f $X=12.145 $Y=1.65 $X2=0
+ $Y2=0
cc_725 N_A_2352_81#_M1012_g N_VGND_c_1440_n 0.0456523f $X=14.215 $Y=1.01 $X2=0
+ $Y2=0
cc_726 N_A_2352_81#_M1001_g N_VGND_c_1442_n 0.0109247f $X=12.01 $Y=0.745 $X2=0
+ $Y2=0
cc_727 N_A_2352_81#_M1012_g N_VGND_c_1442_n 0.0128764f $X=14.215 $Y=1.01 $X2=0
+ $Y2=0
cc_728 N_A_2352_81#_c_1019_n N_VGND_c_1442_n 0.0328648f $X=13.275 $Y=0.68 $X2=0
+ $Y2=0
cc_729 N_A_2123_543#_M1005_g N_VPWR_c_1213_n 0.0489731f $X=12.885 $Y=3.215 $X2=0
+ $Y2=0
cc_730 N_A_2123_543#_c_1119_n N_VPWR_c_1213_n 0.0744788f $X=12.6 $Y=2.43 $X2=0
+ $Y2=0
cc_731 N_A_2123_543#_c_1113_n N_VPWR_c_1213_n 0.00161905f $X=12.765 $Y=2.01
+ $X2=0 $Y2=0
cc_732 N_A_2123_543#_M1031_d N_VPWR_c_1219_n 4.27145e-19 $X=10.615 $Y=2.715
+ $X2=0 $Y2=0
cc_733 N_A_2123_543#_M1005_g N_VPWR_c_1219_n 0.0120207f $X=12.885 $Y=3.215 $X2=0
+ $Y2=0
cc_734 N_A_2123_543#_c_1122_n N_VPWR_c_1219_n 0.00242262f $X=10.95 $Y=2.91 $X2=0
+ $Y2=0
cc_735 N_A_2123_543#_M1002_g N_Q_c_1392_n 0.00145533f $X=12.885 $Y=0.91 $X2=0
+ $Y2=0
cc_736 N_A_2123_543#_M1005_g N_Q_c_1396_n 0.00180148f $X=12.885 $Y=3.215 $X2=0
+ $Y2=0
cc_737 N_A_2123_543#_M1002_g N_Q_c_1394_n 7.13177e-19 $X=12.885 $Y=0.91 $X2=0
+ $Y2=0
cc_738 N_A_2123_543#_c_1113_n N_Q_c_1399_n 0.00180148f $X=12.765 $Y=2.01 $X2=0
+ $Y2=0
cc_739 N_A_2123_543#_M1002_g N_VGND_c_1438_n 0.0501553f $X=12.885 $Y=0.91 $X2=0
+ $Y2=0
cc_740 N_A_2123_543#_c_1108_n N_VGND_c_1438_n 0.0112758f $X=11.63 $Y=0.58 $X2=0
+ $Y2=0
cc_741 N_A_2123_543#_c_1112_n N_VGND_c_1438_n 0.0463156f $X=11.715 $Y=2.345
+ $X2=0 $Y2=0
cc_742 N_A_2123_543#_M1029_d N_VGND_c_1442_n 0.00392019f $X=10.73 $Y=0.535 $X2=0
+ $Y2=0
cc_743 N_A_2123_543#_M1002_g N_VGND_c_1442_n 0.0122311f $X=12.885 $Y=0.91 $X2=0
+ $Y2=0
cc_744 N_A_2123_543#_c_1108_n N_VGND_c_1442_n 0.0519738f $X=11.63 $Y=0.58 $X2=0
+ $Y2=0
cc_745 N_A_2123_543#_c_1110_n N_VGND_c_1442_n 0.0260915f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_746 N_A_2123_543#_c_1108_n A_2310_107# 8.39422e-19 $X=11.63 $Y=0.58 $X2=0
+ $Y2=0
cc_747 N_A_2123_543#_c_1112_n A_2310_107# 0.00359332f $X=11.715 $Y=2.345 $X2=0
+ $Y2=0
cc_748 N_VPWR_c_1201_n A_343_593# 0.00579442f $X=1.075 $Y=3.175 $X2=0 $Y2=3.985
cc_749 N_VPWR_c_1204_n N_A_484_107#_c_1303_n 0.00557519f $X=4.15 $Y=3.11
+ $X2=14.64 $Y2=4.07
cc_750 N_VPWR_c_1219_n N_A_484_107#_c_1303_n 0.0255822f $X=14.675 $Y=3.59
+ $X2=14.64 $Y2=4.07
cc_751 N_VPWR_c_1201_n N_A_484_107#_c_1306_n 0.0168228f $X=1.075 $Y=3.175 $X2=0
+ $Y2=0
cc_752 N_VPWR_c_1219_n N_A_484_107#_c_1306_n 0.0144801f $X=14.675 $Y=3.59 $X2=0
+ $Y2=0
cc_753 N_VPWR_c_1219_n N_A_484_107#_c_1310_n 0.00227751f $X=14.675 $Y=3.59 $X2=0
+ $Y2=0
cc_754 N_VPWR_c_1219_n N_Q_c_1396_n 0.0411361f $X=14.675 $Y=3.59 $X2=14.64
+ $Y2=4.07
cc_755 N_VPWR_c_1216_n N_Q_c_1399_n 0.112136f $X=14.605 $Y=2.36 $X2=7.44
+ $Y2=4.013
cc_756 N_VPWR_c_1216_n Q 0.0237314f $X=14.605 $Y=2.36 $X2=0 $Y2=0
cc_757 N_A_484_107#_c_1303_n A_641_593# 0.00178739f $X=3.23 $Y=3.01 $X2=0 $Y2=0
cc_758 N_A_484_107#_c_1299_n N_VGND_c_1430_n 0.0117552f $X=2.56 $Y=0.745 $X2=0
+ $Y2=0
cc_759 N_A_484_107#_c_1296_n N_VGND_c_1432_n 0.00461294f $X=3.315 $Y=1.865 $X2=0
+ $Y2=0
cc_760 N_A_484_107#_M1028_s N_VGND_c_1442_n 0.00225203f $X=6.585 $Y=0.535 $X2=0
+ $Y2=0
cc_761 N_A_484_107#_c_1295_n N_VGND_c_1442_n 0.0239592f $X=3.23 $Y=0.83 $X2=0
+ $Y2=0
cc_762 N_A_484_107#_c_1299_n N_VGND_c_1442_n 0.0308296f $X=2.56 $Y=0.745 $X2=0
+ $Y2=0
cc_763 N_A_484_107#_c_1302_n N_VGND_c_1442_n 0.0220848f $X=6.73 $Y=0.765 $X2=0
+ $Y2=0
cc_764 N_A_484_107#_c_1295_n A_640_107# 0.00169137f $X=3.23 $Y=0.83 $X2=0 $Y2=0
cc_765 N_Q_c_1392_n N_VGND_c_1440_n 0.0534224f $X=13.825 $Y=0.78 $X2=0 $Y2=0
cc_766 Q N_VGND_c_1440_n 0.0412128f $X=14.555 $Y=1.58 $X2=0 $Y2=0
cc_767 N_Q_c_1392_n N_VGND_c_1442_n 0.0283453f $X=13.825 $Y=0.78 $X2=0 $Y2=0
cc_768 N_VGND_c_1430_n A_342_107# 0.00604574f $X=1.74 $Y=0.48 $X2=0 $Y2=0
cc_769 N_VGND_c_1442_n A_342_107# 8.10341e-19 $X=14.675 $Y=0.48 $X2=0 $Y2=0
cc_770 N_VGND_c_1442_n A_640_107# 0.00206734f $X=14.675 $Y=0.48 $X2=0 $Y2=0
cc_771 N_VGND_c_1442_n A_1646_107# 0.00875788f $X=14.675 $Y=0.48 $X2=0 $Y2=0
