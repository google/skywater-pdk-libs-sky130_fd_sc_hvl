* File: sky130_fd_sc_hvl__buf_8.pxi.spice
* Created: Fri Aug 28 09:33:32 2020
* 
x_PM_SKY130_FD_SC_HVL__BUF_8%VNB N_VNB_M1003_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__BUF_8%VNB
x_PM_SKY130_FD_SC_HVL__BUF_8%VPB N_VPB_M1006_b VPB N_VPB_c_43_p VPB
+ PM_SKY130_FD_SC_HVL__BUF_8%VPB
x_PM_SKY130_FD_SC_HVL__BUF_8%A N_A_M1006_g N_A_c_123_n N_A_M1003_g N_A_c_125_n
+ N_A_c_126_n N_A_M1008_g N_A_M1007_g N_A_c_127_n N_A_M1015_g N_A_M1019_g
+ N_A_c_128_n A A A A N_A_c_129_n PM_SKY130_FD_SC_HVL__BUF_8%A
x_PM_SKY130_FD_SC_HVL__BUF_8%A_45_443# N_A_45_443#_M1003_d N_A_45_443#_M1008_d
+ N_A_45_443#_M1006_s N_A_45_443#_M1007_s N_A_45_443#_M1001_g
+ N_A_45_443#_c_206_n N_A_45_443#_M1000_g N_A_45_443#_M1002_g
+ N_A_45_443#_c_209_n N_A_45_443#_M1004_g N_A_45_443#_M1009_g
+ N_A_45_443#_c_212_n N_A_45_443#_M1005_g N_A_45_443#_M1013_g
+ N_A_45_443#_c_215_n N_A_45_443#_M1010_g N_A_45_443#_M1014_g
+ N_A_45_443#_c_218_n N_A_45_443#_M1011_g N_A_45_443#_M1018_g
+ N_A_45_443#_c_221_n N_A_45_443#_M1012_g N_A_45_443#_M1020_g
+ N_A_45_443#_c_224_n N_A_45_443#_M1016_g N_A_45_443#_M1021_g
+ N_A_45_443#_c_227_n N_A_45_443#_M1017_g N_A_45_443#_c_240_n
+ N_A_45_443#_c_202_n N_A_45_443#_c_231_n N_A_45_443#_c_233_n
+ N_A_45_443#_c_248_n N_A_45_443#_c_374_p N_A_45_443#_c_250_n
+ N_A_45_443#_c_254_n N_A_45_443#_c_203_n N_A_45_443#_c_204_n
+ N_A_45_443#_c_235_n N_A_45_443#_c_236_n N_A_45_443#_c_261_n
+ N_A_45_443#_c_264_n N_A_45_443#_c_205_n PM_SKY130_FD_SC_HVL__BUF_8%A_45_443#
x_PM_SKY130_FD_SC_HVL__BUF_8%VPWR N_VPWR_M1006_d N_VPWR_M1019_d N_VPWR_M1004_s
+ N_VPWR_M1010_s N_VPWR_M1012_s N_VPWR_M1017_s N_VPWR_c_417_n N_VPWR_c_420_n
+ N_VPWR_c_423_n N_VPWR_c_426_n N_VPWR_c_429_n N_VPWR_c_430_n N_VPWR_c_431_n
+ N_VPWR_c_434_n N_VPWR_c_437_n N_VPWR_c_440_n VPWR N_VPWR_c_455_n
+ N_VPWR_c_485_n N_VPWR_c_490_n N_VPWR_c_495_n N_VPWR_c_443_n N_VPWR_c_446_n
+ N_VPWR_c_449_n PM_SKY130_FD_SC_HVL__BUF_8%VPWR
x_PM_SKY130_FD_SC_HVL__BUF_8%X N_X_M1001_d N_X_M1009_d N_X_M1014_d N_X_M1020_d
+ N_X_M1000_d N_X_M1005_d N_X_M1011_d N_X_M1016_d N_X_c_547_n N_X_c_540_n
+ N_X_c_552_n N_X_c_553_n N_X_c_544_n N_X_c_558_n N_X_c_561_n N_X_c_541_n
+ N_X_c_566_n N_X_c_545_n N_X_c_570_n N_X_c_542_n N_X_c_575_n N_X_c_546_n
+ N_X_c_631_p N_X_c_543_n N_X_c_582_n N_X_c_583_n N_X_c_586_n N_X_c_587_n
+ N_X_c_590_n X X X X X X X N_X_c_598_n N_X_c_599_n PM_SKY130_FD_SC_HVL__BUF_8%X
x_PM_SKY130_FD_SC_HVL__BUF_8%VGND N_VGND_M1003_s N_VGND_M1015_s N_VGND_M1002_s
+ N_VGND_M1013_s N_VGND_M1018_s N_VGND_M1021_s N_VGND_c_640_n N_VGND_c_641_n
+ VGND N_VGND_c_642_n N_VGND_c_644_n N_VGND_c_646_n N_VGND_c_648_n
+ N_VGND_c_649_n N_VGND_c_650_n N_VGND_c_651_n N_VGND_c_652_n N_VGND_c_653_n
+ N_VGND_c_654_n N_VGND_c_655_n PM_SKY130_FD_SC_HVL__BUF_8%VGND
cc_1 N_VNB_M1003_b N_A_c_123_n 0.0456634f $X=-0.33 $Y=-0.265 $X2=0.78 $Y2=1.565
cc_2 N_VNB_c_2_p N_A_c_123_n 5.58874e-19 $X=0.24 $Y=0 $X2=0.78 $Y2=1.565
cc_3 N_VNB_M1003_b N_A_c_125_n 0.0274014f $X=-0.33 $Y=-0.265 $X2=1.57 $Y2=1.815
cc_4 N_VNB_M1003_b N_A_c_126_n 0.0391903f $X=-0.33 $Y=-0.265 $X2=1.82 $Y2=1.565
cc_5 N_VNB_M1003_b N_A_c_127_n 0.0378062f $X=-0.33 $Y=-0.265 $X2=2.6 $Y2=1.565
cc_6 N_VNB_M1003_b N_A_c_128_n 0.0267973f $X=-0.33 $Y=-0.265 $X2=0.77 $Y2=1.815
cc_7 N_VNB_M1003_b N_A_c_129_n 0.0506531f $X=-0.33 $Y=-0.265 $X2=2.6 $Y2=1.815
cc_8 N_VNB_M1003_b N_A_45_443#_M1001_g 0.0409882f $X=-0.33 $Y=-0.265 $X2=1.82
+ $Y2=2.965
cc_9 N_VNB_M1003_b N_A_45_443#_M1002_g 0.0406374f $X=-0.33 $Y=-0.265 $X2=2.6
+ $Y2=2.965
cc_10 N_VNB_M1003_b N_A_45_443#_M1009_g 0.0406374f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1003_b N_A_45_443#_M1013_g 0.0406374f $X=-0.33 $Y=-0.265 $X2=1.82
+ $Y2=1.815
cc_12 N_VNB_M1003_b N_A_45_443#_M1014_g 0.0406374f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1003_b N_A_45_443#_M1018_g 0.0406374f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_M1003_b N_A_45_443#_M1020_g 0.0400078f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_15 N_VNB_M1003_b N_A_45_443#_M1021_g 0.0475743f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_16 N_VNB_M1003_b N_A_45_443#_c_202_n 0.0201484f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_17 N_VNB_M1003_b N_A_45_443#_c_203_n 0.00264768f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1003_b N_A_45_443#_c_204_n 0.00132121f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_19 N_VNB_M1003_b N_A_45_443#_c_205_n 0.215377f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_20 N_VNB_M1003_b N_X_c_540_n 0.00276601f $X=-0.33 $Y=-0.265 $X2=1.735
+ $Y2=1.815
cc_21 N_VNB_M1003_b N_X_c_541_n 0.00276601f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_22 N_VNB_M1003_b N_X_c_542_n 0.00276601f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_23 N_VNB_M1003_b N_X_c_543_n 0.00201572f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_24 N_VNB_M1003_b N_VGND_c_640_n 0.0113819f $X=-0.33 $Y=-0.265 $X2=2.6
+ $Y2=1.08
cc_25 N_VNB_M1003_b N_VGND_c_641_n 0.0421164f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_26 N_VNB_M1003_b N_VGND_c_642_n 0.090476f $X=-0.33 $Y=-0.265 $X2=1.68
+ $Y2=1.697
cc_27 N_VNB_c_2_p N_VGND_c_642_n 0.00538291f $X=0.24 $Y=0 $X2=1.68 $Y2=1.697
cc_28 N_VNB_M1003_b N_VGND_c_644_n 0.0421797f $X=-0.33 $Y=-0.265 $X2=2.16
+ $Y2=1.697
cc_29 N_VNB_c_2_p N_VGND_c_644_n 0.00247336f $X=0.24 $Y=0 $X2=2.16 $Y2=1.697
cc_30 N_VNB_M1003_b N_VGND_c_646_n 0.251101f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_31 N_VNB_c_2_p N_VGND_c_646_n 0.0168113f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_32 N_VNB_M1003_b N_VGND_c_648_n 0.00648157f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_33 N_VNB_M1003_b N_VGND_c_649_n 0.00846255f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_34 N_VNB_M1003_b N_VGND_c_650_n 0.00648157f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_35 N_VNB_M1003_b N_VGND_c_651_n 0.00846255f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_36 N_VNB_M1003_b N_VGND_c_652_n 0.00659769f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_37 N_VNB_M1003_b N_VGND_c_653_n 0.0125522f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_38 N_VNB_M1003_b N_VGND_c_654_n 0.00867563f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_39 N_VNB_M1003_b N_VGND_c_655_n 0.152445f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_40 N_VNB_c_2_p N_VGND_c_655_n 1.02625f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_41 N_VPB_M1006_b N_A_M1006_g 0.0429652f $X=-0.33 $Y=1.885 $X2=0.76 $Y2=2.965
cc_42 VPB N_A_M1006_g 0.00970178f $X=0 $Y=3.955 $X2=0.76 $Y2=2.965
cc_43 N_VPB_c_43_p N_A_M1006_g 0.0148199f $X=9.36 $Y=4.07 $X2=0.76 $Y2=2.965
cc_44 N_VPB_M1006_b N_A_c_125_n 0.0193995f $X=-0.33 $Y=1.885 $X2=1.57 $Y2=1.815
cc_45 N_VPB_M1006_b N_A_M1007_g 0.0378158f $X=-0.33 $Y=1.885 $X2=1.82 $Y2=2.965
cc_46 VPB N_A_M1007_g 0.00970178f $X=0 $Y=3.955 $X2=1.82 $Y2=2.965
cc_47 N_VPB_c_43_p N_A_M1007_g 0.013528f $X=9.36 $Y=4.07 $X2=1.82 $Y2=2.965
cc_48 N_VPB_M1006_b N_A_M1019_g 0.0364141f $X=-0.33 $Y=1.885 $X2=2.6 $Y2=2.965
cc_49 VPB N_A_M1019_g 0.00970178f $X=0 $Y=3.955 $X2=2.6 $Y2=2.965
cc_50 N_VPB_c_43_p N_A_M1019_g 0.0135178f $X=9.36 $Y=4.07 $X2=2.6 $Y2=2.965
cc_51 N_VPB_M1006_b N_A_c_128_n 0.0144517f $X=-0.33 $Y=1.885 $X2=0.77 $Y2=1.815
cc_52 N_VPB_M1006_b N_A_c_129_n 0.0299911f $X=-0.33 $Y=1.885 $X2=2.6 $Y2=1.815
cc_53 N_VPB_M1006_b N_A_45_443#_c_206_n 0.0328513f $X=-0.33 $Y=1.885 $X2=2.6
+ $Y2=1.565
cc_54 VPB N_A_45_443#_c_206_n 0.00970178f $X=0 $Y=3.955 $X2=2.6 $Y2=1.565
cc_55 N_VPB_c_43_p N_A_45_443#_c_206_n 0.0135156f $X=9.36 $Y=4.07 $X2=2.6
+ $Y2=1.565
cc_56 N_VPB_M1006_b N_A_45_443#_c_209_n 0.0321055f $X=-0.33 $Y=1.885 $X2=0.77
+ $Y2=1.815
cc_57 VPB N_A_45_443#_c_209_n 0.00970178f $X=0 $Y=3.955 $X2=0.77 $Y2=1.815
cc_58 N_VPB_c_43_p N_A_45_443#_c_209_n 0.0135156f $X=9.36 $Y=4.07 $X2=0.77
+ $Y2=1.815
cc_59 N_VPB_M1006_b N_A_45_443#_c_212_n 0.0321055f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_60 VPB N_A_45_443#_c_212_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_61 N_VPB_c_43_p N_A_45_443#_c_212_n 0.0135156f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_62 N_VPB_M1006_b N_A_45_443#_c_215_n 0.0321055f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_63 VPB N_A_45_443#_c_215_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_64 N_VPB_c_43_p N_A_45_443#_c_215_n 0.0135156f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_65 N_VPB_M1006_b N_A_45_443#_c_218_n 0.0321055f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_66 VPB N_A_45_443#_c_218_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_67 N_VPB_c_43_p N_A_45_443#_c_218_n 0.0135156f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_68 N_VPB_M1006_b N_A_45_443#_c_221_n 0.0321055f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_69 VPB N_A_45_443#_c_221_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_70 N_VPB_c_43_p N_A_45_443#_c_221_n 0.0135156f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_71 N_VPB_M1006_b N_A_45_443#_c_224_n 0.0321055f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_72 VPB N_A_45_443#_c_224_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_73 N_VPB_c_43_p N_A_45_443#_c_224_n 0.0135156f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_74 N_VPB_M1006_b N_A_45_443#_c_227_n 0.0390747f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_75 VPB N_A_45_443#_c_227_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_76 N_VPB_c_43_p N_A_45_443#_c_227_n 0.0135186f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_77 N_VPB_M1006_b N_A_45_443#_c_202_n 0.00998322f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_78 VPB N_A_45_443#_c_231_n 4.22267e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_79 N_VPB_c_43_p N_A_45_443#_c_231_n 0.00452125f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_80 N_VPB_M1006_b N_A_45_443#_c_233_n 0.00764217f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_81 N_VPB_M1006_b N_A_45_443#_c_203_n 0.00381808f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_82 N_VPB_M1006_b N_A_45_443#_c_235_n 0.00526456f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_83 N_VPB_M1006_b N_A_45_443#_c_236_n 0.00544073f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_84 N_VPB_M1006_b N_A_45_443#_c_205_n 0.17523f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_85 N_VPB_M1006_b N_VPWR_c_417_n 0.0010569f $X=-0.33 $Y=1.885 $X2=2.6 $Y2=1.08
cc_86 VPB N_VPWR_c_417_n 0.00362936f $X=0 $Y=3.955 $X2=2.6 $Y2=1.08
cc_87 N_VPB_c_43_p N_VPWR_c_417_n 0.054215f $X=9.36 $Y=4.07 $X2=2.6 $Y2=1.08
cc_88 N_VPB_M1006_b N_VPWR_c_420_n 0.0010569f $X=-0.33 $Y=1.885 $X2=2.6
+ $Y2=2.965
cc_89 VPB N_VPWR_c_420_n 0.00262607f $X=0 $Y=3.955 $X2=2.6 $Y2=2.965
cc_90 N_VPB_c_43_p N_VPWR_c_420_n 0.0405322f $X=9.36 $Y=4.07 $X2=2.6 $Y2=2.965
cc_91 N_VPB_M1006_b N_VPWR_c_423_n 0.0010569f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_423_n 0.00262607f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_93 N_VPB_c_43_p N_VPWR_c_423_n 0.0405322f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_94 N_VPB_M1006_b N_VPWR_c_426_n 0.0010569f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_95 VPB N_VPWR_c_426_n 0.00262607f $X=0 $Y=3.955 $X2=0.635 $Y2=1.58
cc_96 N_VPB_c_43_p N_VPWR_c_426_n 0.0405322f $X=9.36 $Y=4.07 $X2=0.635 $Y2=1.58
cc_97 N_VPB_M1006_b N_VPWR_c_429_n 0.00769488f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_98 N_VPB_M1006_b N_VPWR_c_430_n 0.0525239f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_99 N_VPB_M1006_b N_VPWR_c_431_n 0.00105831f $X=-0.33 $Y=1.885 $X2=1.82
+ $Y2=1.815
cc_100 VPB N_VPWR_c_431_n 0.00279423f $X=0 $Y=3.955 $X2=1.82 $Y2=1.815
cc_101 N_VPB_c_43_p N_VPWR_c_431_n 0.0413412f $X=9.36 $Y=4.07 $X2=1.82 $Y2=1.815
cc_102 N_VPB_M1006_b N_VPWR_c_434_n 0.00105831f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_434_n 0.00385318f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_104 N_VPB_c_43_p N_VPWR_c_434_n 0.0545489f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_105 N_VPB_M1006_b N_VPWR_c_437_n 0.00105831f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_437_n 0.00385318f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_107 N_VPB_c_43_p N_VPWR_c_437_n 0.0545489f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_108 N_VPB_M1006_b N_VPWR_c_440_n 0.00105831f $X=-0.33 $Y=1.885 $X2=1.2
+ $Y2=1.697
cc_109 VPB N_VPWR_c_440_n 0.00385318f $X=0 $Y=3.955 $X2=1.2 $Y2=1.697
cc_110 N_VPB_c_43_p N_VPWR_c_440_n 0.0545489f $X=9.36 $Y=4.07 $X2=1.2 $Y2=1.697
cc_111 N_VPB_M1006_b N_VPWR_c_443_n 0.00270841f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_443_n 0.00513943f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_113 N_VPB_c_43_p N_VPWR_c_443_n 0.0771568f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_114 N_VPB_M1006_b N_VPWR_c_446_n 0.0010569f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_446_n 0.00535847f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_116 N_VPB_c_43_p N_VPWR_c_446_n 0.0847751f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_117 N_VPB_M1006_b N_VPWR_c_449_n 0.0587432f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_449_n 1.01609f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_119 N_VPB_c_43_p N_VPWR_c_449_n 0.033555f $X=9.36 $Y=4.07 $X2=0 $Y2=0
cc_120 N_VPB_M1006_b N_X_c_544_n 0.00261732f $X=-0.33 $Y=1.885 $X2=2.6 $Y2=1.815
cc_121 N_VPB_M1006_b N_X_c_545_n 0.00261732f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_122 N_VPB_M1006_b N_X_c_546_n 0.00261732f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_123 N_A_c_127_n N_A_45_443#_M1001_g 0.0206089f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_124 N_A_M1019_g N_A_45_443#_c_206_n 0.0206089f $X=2.6 $Y=2.965 $X2=9.36 $Y2=0
cc_125 N_A_c_123_n N_A_45_443#_c_240_n 0.00436519f $X=0.78 $Y=1.565 $X2=0 $Y2=0
cc_126 N_A_c_123_n N_A_45_443#_c_202_n 0.00386514f $X=0.78 $Y=1.565 $X2=0 $Y2=0
cc_127 N_A_c_128_n N_A_45_443#_c_202_n 0.0206904f $X=0.77 $Y=1.815 $X2=0 $Y2=0
cc_128 A N_A_45_443#_c_202_n 0.0165919f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A_M1006_g N_A_45_443#_c_233_n 0.0358157f $X=0.76 $Y=2.965 $X2=0 $Y2=0
cc_130 N_A_c_125_n N_A_45_443#_c_233_n 0.011632f $X=1.57 $Y=1.815 $X2=0 $Y2=0
cc_131 N_A_M1007_g N_A_45_443#_c_233_n 0.0313016f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_132 A N_A_45_443#_c_233_n 0.0678558f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A_M1007_g N_A_45_443#_c_248_n 0.0260651f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_134 N_A_M1019_g N_A_45_443#_c_248_n 0.0459046f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_135 N_A_c_126_n N_A_45_443#_c_250_n 9.17632e-19 $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_136 N_A_c_127_n N_A_45_443#_c_250_n 0.00807427f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_137 A N_A_45_443#_c_250_n 0.00316816f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A_c_129_n N_A_45_443#_c_250_n 0.00326877f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_139 N_A_M1019_g N_A_45_443#_c_254_n 0.00132085f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_140 N_A_c_129_n N_A_45_443#_c_254_n 0.00843589f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_141 N_A_c_129_n N_A_45_443#_c_203_n 0.0311559f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_142 N_A_M1007_g N_A_45_443#_c_236_n 0.00229199f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_143 N_A_M1019_g N_A_45_443#_c_236_n 0.0126893f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_144 A N_A_45_443#_c_236_n 0.0112571f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_145 N_A_c_129_n N_A_45_443#_c_236_n 0.00355898f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_146 N_A_c_127_n N_A_45_443#_c_261_n 0.01573f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_147 A N_A_45_443#_c_261_n 0.00887026f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A_c_129_n N_A_45_443#_c_261_n 0.00269586f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_149 A N_A_45_443#_c_264_n 0.0152738f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A_c_129_n N_A_45_443#_c_264_n 0.0154167f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_151 N_A_c_129_n N_A_45_443#_c_205_n 0.0206089f $X=2.6 $Y=1.815 $X2=0 $Y2=0
cc_152 N_A_M1007_g N_VPWR_c_417_n 0.0103088f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_153 N_A_M1019_g N_VPWR_c_417_n 0.0156302f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_154 N_A_M1019_g N_VPWR_c_431_n 0.00249815f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_155 N_A_M1007_g N_VPWR_c_455_n 7.78697e-19 $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_156 N_A_M1019_g N_VPWR_c_455_n 0.030772f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_157 N_A_M1006_g N_VPWR_c_443_n 0.0716973f $X=0.76 $Y=2.965 $X2=0 $Y2=0
cc_158 N_A_M1007_g N_VPWR_c_443_n 0.0862897f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_159 N_A_M1019_g N_VPWR_c_443_n 0.00121482f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_160 N_A_M1006_g N_VPWR_c_449_n 0.00951892f $X=0.76 $Y=2.965 $X2=0 $Y2=0
cc_161 N_A_M1007_g N_VPWR_c_449_n 0.010513f $X=1.82 $Y=2.965 $X2=0 $Y2=0
cc_162 N_A_M1019_g N_VPWR_c_449_n 0.010744f $X=2.6 $Y=2.965 $X2=0 $Y2=0
cc_163 N_A_c_126_n N_VGND_c_640_n 0.00367492f $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_164 N_A_c_127_n N_VGND_c_640_n 0.00793008f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_165 N_A_c_123_n N_VGND_c_642_n 0.0572185f $X=0.78 $Y=1.565 $X2=0 $Y2=0
cc_166 N_A_c_125_n N_VGND_c_642_n 0.00914385f $X=1.57 $Y=1.815 $X2=0 $Y2=0
cc_167 N_A_c_126_n N_VGND_c_642_n 0.0624717f $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_168 N_A_c_127_n N_VGND_c_642_n 6.48731e-19 $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_169 A N_VGND_c_642_n 0.0836537f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_170 N_A_c_126_n N_VGND_c_644_n 4.13084e-19 $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_171 N_A_c_127_n N_VGND_c_644_n 0.0408201f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_172 N_A_c_123_n N_VGND_c_655_n 0.00915616f $X=0.78 $Y=1.565 $X2=0 $Y2=0
cc_173 N_A_c_126_n N_VGND_c_655_n 0.00865748f $X=1.82 $Y=1.565 $X2=0 $Y2=0
cc_174 N_A_c_127_n N_VGND_c_655_n 0.00795556f $X=2.6 $Y=1.565 $X2=0 $Y2=0
cc_175 N_A_45_443#_c_233_n N_VPWR_M1006_d 0.00539862f $X=2.045 $Y=2.18 $X2=0
+ $Y2=0
cc_176 N_A_45_443#_M1007_s N_VPWR_c_417_n 8.28689e-19 $X=2.07 $Y=2.215 $X2=0
+ $Y2=0
cc_177 N_A_45_443#_c_248_n N_VPWR_c_417_n 0.0314378f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_178 N_A_45_443#_c_206_n N_VPWR_c_420_n 0.00981852f $X=3.38 $Y=2.105 $X2=4.8
+ $Y2=0
cc_179 N_A_45_443#_c_209_n N_VPWR_c_420_n 0.00984257f $X=4.16 $Y=2.105 $X2=4.8
+ $Y2=0
cc_180 N_A_45_443#_c_212_n N_VPWR_c_423_n 0.00984257f $X=4.94 $Y=2.105 $X2=4.8
+ $Y2=0.057
cc_181 N_A_45_443#_c_215_n N_VPWR_c_423_n 0.00984257f $X=5.72 $Y=2.105 $X2=4.8
+ $Y2=0.057
cc_182 N_A_45_443#_c_218_n N_VPWR_c_426_n 0.00984257f $X=6.5 $Y=2.105 $X2=4.8
+ $Y2=0.058
cc_183 N_A_45_443#_c_221_n N_VPWR_c_426_n 0.00984257f $X=7.28 $Y=2.105 $X2=4.8
+ $Y2=0.058
cc_184 N_A_45_443#_c_224_n N_VPWR_c_429_n 7.80614e-19 $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_185 N_A_45_443#_c_227_n N_VPWR_c_429_n 0.014504f $X=8.84 $Y=2.105 $X2=0 $Y2=0
cc_186 N_A_45_443#_c_206_n N_VPWR_c_431_n 0.00656115f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_187 N_A_45_443#_c_209_n N_VPWR_c_434_n 0.00656544f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_188 N_A_45_443#_c_212_n N_VPWR_c_434_n 0.00656544f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_189 N_A_45_443#_c_215_n N_VPWR_c_437_n 0.00656544f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_190 N_A_45_443#_c_218_n N_VPWR_c_437_n 0.00656544f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_191 N_A_45_443#_c_221_n N_VPWR_c_440_n 0.00656544f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_192 N_A_45_443#_c_224_n N_VPWR_c_440_n 0.00656544f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_193 N_A_45_443#_c_206_n N_VPWR_c_455_n 0.0613454f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_194 N_A_45_443#_c_209_n N_VPWR_c_455_n 4.52391e-19 $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_195 N_A_45_443#_c_248_n N_VPWR_c_455_n 0.0873251f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_196 N_A_45_443#_c_203_n N_VPWR_c_455_n 0.0224182f $X=3.295 $Y=1.79 $X2=0
+ $Y2=0
cc_197 N_A_45_443#_c_206_n N_VPWR_c_485_n 4.54877e-19 $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_198 N_A_45_443#_c_209_n N_VPWR_c_485_n 0.0570434f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_199 N_A_45_443#_c_212_n N_VPWR_c_485_n 0.0570434f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_200 N_A_45_443#_c_215_n N_VPWR_c_485_n 4.54877e-19 $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_201 N_A_45_443#_c_205_n N_VPWR_c_485_n 6.12604e-19 $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_202 N_A_45_443#_c_212_n N_VPWR_c_490_n 4.54877e-19 $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_203 N_A_45_443#_c_215_n N_VPWR_c_490_n 0.0570434f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_204 N_A_45_443#_c_218_n N_VPWR_c_490_n 0.0570434f $X=6.5 $Y=2.105 $X2=0 $Y2=0
cc_205 N_A_45_443#_c_221_n N_VPWR_c_490_n 4.54877e-19 $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_206 N_A_45_443#_c_205_n N_VPWR_c_490_n 6.12604e-19 $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_207 N_A_45_443#_c_218_n N_VPWR_c_495_n 4.54877e-19 $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_208 N_A_45_443#_c_221_n N_VPWR_c_495_n 0.0570434f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_209 N_A_45_443#_c_224_n N_VPWR_c_495_n 0.0581256f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_210 N_A_45_443#_c_227_n N_VPWR_c_495_n 0.0011619f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_211 N_A_45_443#_c_205_n N_VPWR_c_495_n 6.12604e-19 $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_212 N_A_45_443#_c_231_n N_VPWR_c_443_n 0.0817667f $X=0.35 $Y=2.36 $X2=0 $Y2=0
cc_213 N_A_45_443#_c_233_n N_VPWR_c_443_n 0.0847738f $X=2.045 $Y=2.18 $X2=0
+ $Y2=0
cc_214 N_A_45_443#_c_248_n N_VPWR_c_443_n 0.0787997f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_215 N_A_45_443#_c_224_n N_VPWR_c_446_n 0.0098265f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_216 N_A_45_443#_c_227_n N_VPWR_c_446_n 0.0115186f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_217 N_A_45_443#_M1006_s N_VPWR_c_449_n 0.00425071f $X=0.225 $Y=2.215 $X2=0
+ $Y2=0
cc_218 N_A_45_443#_c_206_n N_VPWR_c_449_n 0.00994558f $X=3.38 $Y=2.105 $X2=0
+ $Y2=0
cc_219 N_A_45_443#_c_209_n N_VPWR_c_449_n 0.00994001f $X=4.16 $Y=2.105 $X2=0
+ $Y2=0
cc_220 N_A_45_443#_c_212_n N_VPWR_c_449_n 0.00994001f $X=4.94 $Y=2.105 $X2=0
+ $Y2=0
cc_221 N_A_45_443#_c_215_n N_VPWR_c_449_n 0.00994001f $X=5.72 $Y=2.105 $X2=0
+ $Y2=0
cc_222 N_A_45_443#_c_218_n N_VPWR_c_449_n 0.00994001f $X=6.5 $Y=2.105 $X2=0
+ $Y2=0
cc_223 N_A_45_443#_c_221_n N_VPWR_c_449_n 0.00994001f $X=7.28 $Y=2.105 $X2=0
+ $Y2=0
cc_224 N_A_45_443#_c_224_n N_VPWR_c_449_n 0.00989505f $X=8.06 $Y=2.105 $X2=0
+ $Y2=0
cc_225 N_A_45_443#_c_227_n N_VPWR_c_449_n 0.0107477f $X=8.84 $Y=2.105 $X2=0
+ $Y2=0
cc_226 N_A_45_443#_c_231_n N_VPWR_c_449_n 0.0196936f $X=0.35 $Y=2.36 $X2=0 $Y2=0
cc_227 N_A_45_443#_c_248_n N_VPWR_c_449_n 0.0205648f $X=2.21 $Y=2.34 $X2=0 $Y2=0
cc_228 N_A_45_443#_c_206_n N_X_c_547_n 0.0259143f $X=3.38 $Y=2.105 $X2=0 $Y2=0
cc_229 N_A_45_443#_c_209_n N_X_c_547_n 0.0259143f $X=4.16 $Y=2.105 $X2=0 $Y2=0
cc_230 N_A_45_443#_M1001_g N_X_c_540_n 0.00400399f $X=3.38 $Y=1.08 $X2=0 $Y2=0
cc_231 N_A_45_443#_M1002_g N_X_c_540_n 0.00400399f $X=4.16 $Y=1.08 $X2=0 $Y2=0
cc_232 N_A_45_443#_c_205_n N_X_c_540_n 0.00453979f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_233 N_A_45_443#_c_205_n N_X_c_552_n 0.0696897f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_234 N_A_45_443#_c_203_n N_X_c_553_n 0.00942964f $X=3.295 $Y=1.79 $X2=0 $Y2=0
cc_235 N_A_45_443#_c_205_n N_X_c_553_n 0.00967184f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_236 N_A_45_443#_c_209_n N_X_c_544_n 0.0173368f $X=4.16 $Y=2.105 $X2=0 $Y2=0
cc_237 N_A_45_443#_c_212_n N_X_c_544_n 0.0173368f $X=4.94 $Y=2.105 $X2=0 $Y2=0
cc_238 N_A_45_443#_c_205_n N_X_c_544_n 0.0279996f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_239 N_A_45_443#_c_206_n N_X_c_558_n 0.0062277f $X=3.38 $Y=2.105 $X2=0 $Y2=0
cc_240 N_A_45_443#_c_209_n N_X_c_558_n 0.00141551f $X=4.16 $Y=2.105 $X2=0 $Y2=0
cc_241 N_A_45_443#_c_205_n N_X_c_558_n 0.0151427f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_242 N_A_45_443#_c_212_n N_X_c_561_n 0.0259143f $X=4.94 $Y=2.105 $X2=0 $Y2=0
cc_243 N_A_45_443#_c_215_n N_X_c_561_n 0.0259143f $X=5.72 $Y=2.105 $X2=0 $Y2=0
cc_244 N_A_45_443#_M1009_g N_X_c_541_n 0.00400399f $X=4.94 $Y=1.08 $X2=0 $Y2=0
cc_245 N_A_45_443#_M1013_g N_X_c_541_n 0.00400399f $X=5.72 $Y=1.08 $X2=0 $Y2=0
cc_246 N_A_45_443#_c_205_n N_X_c_541_n 0.00458351f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_247 N_A_45_443#_c_205_n N_X_c_566_n 0.0696897f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_248 N_A_45_443#_c_215_n N_X_c_545_n 0.0173368f $X=5.72 $Y=2.105 $X2=0 $Y2=0
cc_249 N_A_45_443#_c_218_n N_X_c_545_n 0.0173368f $X=6.5 $Y=2.105 $X2=0 $Y2=0
cc_250 N_A_45_443#_c_205_n N_X_c_545_n 0.0279996f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_251 N_A_45_443#_c_218_n N_X_c_570_n 0.0259143f $X=6.5 $Y=2.105 $X2=0 $Y2=0
cc_252 N_A_45_443#_c_221_n N_X_c_570_n 0.0259143f $X=7.28 $Y=2.105 $X2=0 $Y2=0
cc_253 N_A_45_443#_M1014_g N_X_c_542_n 0.00400399f $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_254 N_A_45_443#_M1018_g N_X_c_542_n 0.00400399f $X=7.28 $Y=1.08 $X2=0 $Y2=0
cc_255 N_A_45_443#_c_205_n N_X_c_542_n 0.00458351f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_256 N_A_45_443#_c_205_n N_X_c_575_n 0.0786621f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_257 N_A_45_443#_c_221_n N_X_c_546_n 0.0173368f $X=7.28 $Y=2.105 $X2=0 $Y2=0
cc_258 N_A_45_443#_c_224_n N_X_c_546_n 0.0173368f $X=8.06 $Y=2.105 $X2=0 $Y2=0
cc_259 N_A_45_443#_c_205_n N_X_c_546_n 0.0279996f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_260 N_A_45_443#_M1020_g N_X_c_543_n 0.00400399f $X=8.06 $Y=1.08 $X2=0 $Y2=0
cc_261 N_A_45_443#_M1021_g N_X_c_543_n 0.00133825f $X=8.84 $Y=1.08 $X2=0 $Y2=0
cc_262 N_A_45_443#_c_205_n N_X_c_543_n 0.00399266f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_263 N_A_45_443#_M1021_g N_X_c_582_n 0.0103635f $X=8.84 $Y=1.08 $X2=0 $Y2=0
cc_264 N_A_45_443#_c_212_n N_X_c_583_n 0.00141551f $X=4.94 $Y=2.105 $X2=0 $Y2=0
cc_265 N_A_45_443#_c_215_n N_X_c_583_n 0.00141551f $X=5.72 $Y=2.105 $X2=0 $Y2=0
cc_266 N_A_45_443#_c_205_n N_X_c_583_n 0.00951392f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_267 N_A_45_443#_c_205_n N_X_c_586_n 0.00643395f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_268 N_A_45_443#_c_218_n N_X_c_587_n 0.00141551f $X=6.5 $Y=2.105 $X2=0 $Y2=0
cc_269 N_A_45_443#_c_221_n N_X_c_587_n 0.00141551f $X=7.28 $Y=2.105 $X2=0 $Y2=0
cc_270 N_A_45_443#_c_205_n N_X_c_587_n 0.00951392f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_271 N_A_45_443#_c_205_n N_X_c_590_n 0.00643395f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_272 N_A_45_443#_M1021_g X 0.0291857f $X=8.84 $Y=1.08 $X2=0 $Y2=0
cc_273 N_A_45_443#_c_205_n X 0.0394165f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_274 N_A_45_443#_c_224_n X 0.00141551f $X=8.06 $Y=2.105 $X2=0 $Y2=0
cc_275 N_A_45_443#_c_227_n X 0.00911503f $X=8.84 $Y=2.105 $X2=0 $Y2=0
cc_276 N_A_45_443#_c_205_n X 0.0234141f $X=8.84 $Y=1.855 $X2=0 $Y2=0
cc_277 N_A_45_443#_c_224_n X 0.0094348f $X=8.06 $Y=2.105 $X2=0 $Y2=0
cc_278 N_A_45_443#_c_227_n X 0.0275957f $X=8.84 $Y=2.105 $X2=0 $Y2=0
cc_279 N_A_45_443#_M1021_g N_X_c_598_n 0.00796307f $X=8.84 $Y=1.08 $X2=0 $Y2=0
cc_280 N_A_45_443#_c_224_n N_X_c_599_n 0.0176022f $X=8.06 $Y=2.105 $X2=0 $Y2=0
cc_281 N_A_45_443#_c_227_n N_X_c_599_n 0.0363847f $X=8.84 $Y=2.105 $X2=0 $Y2=0
cc_282 N_A_45_443#_c_374_p N_VGND_c_640_n 0.0122346f $X=2.21 $Y=0.895 $X2=0
+ $Y2=0
cc_283 N_A_45_443#_M1021_g N_VGND_c_641_n 0.00589056f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_284 N_A_45_443#_c_240_n N_VGND_c_642_n 0.0377885f $X=0.37 $Y=0.97 $X2=0 $Y2=0
cc_285 N_A_45_443#_M1001_g N_VGND_c_644_n 0.0568363f $X=3.38 $Y=1.08 $X2=0 $Y2=0
cc_286 N_A_45_443#_M1002_g N_VGND_c_644_n 9.11203e-19 $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_287 N_A_45_443#_c_250_n N_VGND_c_644_n 0.00342789f $X=2.51 $Y=1.625 $X2=0
+ $Y2=0
cc_288 N_A_45_443#_c_203_n N_VGND_c_644_n 0.0438358f $X=3.295 $Y=1.79 $X2=0
+ $Y2=0
cc_289 N_A_45_443#_c_261_n N_VGND_c_644_n 0.0138755f $X=2.51 $Y=1.315 $X2=0
+ $Y2=0
cc_290 N_A_45_443#_M1001_g N_VGND_c_646_n 0.00328808f $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_291 N_A_45_443#_M1002_g N_VGND_c_646_n 0.00328808f $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_292 N_A_45_443#_M1001_g N_VGND_c_648_n 9.10934e-19 $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_293 N_A_45_443#_M1002_g N_VGND_c_648_n 0.0525668f $X=4.16 $Y=1.08 $X2=0 $Y2=0
cc_294 N_A_45_443#_M1009_g N_VGND_c_648_n 0.0525668f $X=4.94 $Y=1.08 $X2=0 $Y2=0
cc_295 N_A_45_443#_M1013_g N_VGND_c_648_n 9.10934e-19 $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_296 N_A_45_443#_c_205_n N_VGND_c_648_n 0.00257674f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_297 N_A_45_443#_M1009_g N_VGND_c_649_n 0.00328808f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_298 N_A_45_443#_M1013_g N_VGND_c_649_n 0.00328808f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_299 N_A_45_443#_M1009_g N_VGND_c_650_n 9.10934e-19 $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_300 N_A_45_443#_M1013_g N_VGND_c_650_n 0.0525668f $X=5.72 $Y=1.08 $X2=0 $Y2=0
cc_301 N_A_45_443#_M1014_g N_VGND_c_650_n 0.0525668f $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_302 N_A_45_443#_M1018_g N_VGND_c_650_n 9.10934e-19 $X=7.28 $Y=1.08 $X2=0
+ $Y2=0
cc_303 N_A_45_443#_c_205_n N_VGND_c_650_n 0.00257674f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_304 N_A_45_443#_M1014_g N_VGND_c_651_n 0.00328808f $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_305 N_A_45_443#_M1018_g N_VGND_c_651_n 0.00328808f $X=7.28 $Y=1.08 $X2=0
+ $Y2=0
cc_306 N_A_45_443#_M1014_g N_VGND_c_652_n 9.10934e-19 $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_307 N_A_45_443#_M1018_g N_VGND_c_652_n 0.0525668f $X=7.28 $Y=1.08 $X2=0 $Y2=0
cc_308 N_A_45_443#_M1020_g N_VGND_c_652_n 0.0532979f $X=8.06 $Y=1.08 $X2=0 $Y2=0
cc_309 N_A_45_443#_M1021_g N_VGND_c_652_n 0.00130456f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_310 N_A_45_443#_c_205_n N_VGND_c_652_n 0.00257674f $X=8.84 $Y=1.855 $X2=0
+ $Y2=0
cc_311 N_A_45_443#_M1020_g N_VGND_c_653_n 0.00520463f $X=8.06 $Y=1.08 $X2=0
+ $Y2=0
cc_312 N_A_45_443#_M1021_g N_VGND_c_653_n 0.00965248f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_313 N_A_45_443#_M1021_g N_VGND_c_654_n 0.00617584f $X=8.84 $Y=1.08 $X2=0
+ $Y2=0
cc_314 N_A_45_443#_M1001_g N_VGND_c_655_n 0.00808151f $X=3.38 $Y=1.08 $X2=0
+ $Y2=0
cc_315 N_A_45_443#_M1002_g N_VGND_c_655_n 0.00808151f $X=4.16 $Y=1.08 $X2=0
+ $Y2=0
cc_316 N_A_45_443#_M1009_g N_VGND_c_655_n 0.00808151f $X=4.94 $Y=1.08 $X2=0
+ $Y2=0
cc_317 N_A_45_443#_M1013_g N_VGND_c_655_n 0.00808151f $X=5.72 $Y=1.08 $X2=0
+ $Y2=0
cc_318 N_A_45_443#_M1014_g N_VGND_c_655_n 0.00808151f $X=6.5 $Y=1.08 $X2=0 $Y2=0
cc_319 N_A_45_443#_M1018_g N_VGND_c_655_n 0.00808151f $X=7.28 $Y=1.08 $X2=0
+ $Y2=0
cc_320 N_A_45_443#_M1020_g N_VGND_c_655_n 0.00808151f $X=8.06 $Y=1.08 $X2=0
+ $Y2=0
cc_321 N_A_45_443#_M1021_g N_VGND_c_655_n 0.0148456f $X=8.84 $Y=1.08 $X2=0 $Y2=0
cc_322 N_A_45_443#_c_240_n N_VGND_c_655_n 0.0118041f $X=0.37 $Y=0.97 $X2=0 $Y2=0
cc_323 N_A_45_443#_c_374_p N_VGND_c_655_n 0.00689067f $X=2.21 $Y=0.895 $X2=0
+ $Y2=0
cc_324 N_A_45_443#_c_261_n N_VGND_c_655_n 0.00762664f $X=2.51 $Y=1.315 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_420_n N_X_M1000_d 8.28689e-19 $X=4.105 $Y=3.71 $X2=0 $Y2=0
cc_326 N_VPWR_c_423_n N_X_M1005_d 8.28689e-19 $X=5.665 $Y=3.71 $X2=0 $Y2=3.955
cc_327 N_VPWR_c_426_n N_X_M1011_d 8.28689e-19 $X=7.225 $Y=3.71 $X2=0 $Y2=0
cc_328 N_VPWR_c_446_n N_X_M1016_d 8.28689e-19 $X=8.905 $Y=3.635 $X2=0.24
+ $Y2=4.07
cc_329 N_VPWR_c_420_n N_X_c_547_n 0.0178796f $X=4.105 $Y=3.71 $X2=0 $Y2=0
cc_330 N_VPWR_c_455_n N_X_c_547_n 0.0840941f $X=2.99 $Y=2.55 $X2=0 $Y2=0
cc_331 N_VPWR_c_485_n N_X_c_547_n 0.0842143f $X=4.55 $Y=2.55 $X2=0 $Y2=0
cc_332 N_VPWR_c_449_n N_X_c_547_n 0.01238f $X=9.35 $Y=3.56 $X2=0 $Y2=0
cc_333 N_VPWR_c_485_n N_X_c_544_n 0.0614512f $X=4.55 $Y=2.55 $X2=0 $Y2=0
cc_334 N_VPWR_c_423_n N_X_c_561_n 0.0178796f $X=5.665 $Y=3.71 $X2=0 $Y2=0
cc_335 N_VPWR_c_485_n N_X_c_561_n 0.0842143f $X=4.55 $Y=2.55 $X2=0 $Y2=0
cc_336 N_VPWR_c_490_n N_X_c_561_n 0.0842143f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_337 N_VPWR_c_449_n N_X_c_561_n 0.01238f $X=9.35 $Y=3.56 $X2=0 $Y2=0
cc_338 N_VPWR_c_490_n N_X_c_545_n 0.0614512f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_339 N_VPWR_c_426_n N_X_c_570_n 0.0178796f $X=7.225 $Y=3.71 $X2=0 $Y2=0
cc_340 N_VPWR_c_490_n N_X_c_570_n 0.0842143f $X=6.11 $Y=2.55 $X2=0 $Y2=0
cc_341 N_VPWR_c_495_n N_X_c_570_n 0.0842143f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_342 N_VPWR_c_449_n N_X_c_570_n 0.01238f $X=9.35 $Y=3.56 $X2=0 $Y2=0
cc_343 N_VPWR_c_495_n N_X_c_546_n 0.0614512f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_344 N_VPWR_c_429_n X 0.0026211f $X=9.32 $Y=3.475 $X2=0 $Y2=0
cc_345 N_VPWR_c_495_n X 0.0462063f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_346 N_VPWR_c_446_n X 0.0292853f $X=8.905 $Y=3.635 $X2=0 $Y2=0
cc_347 N_VPWR_c_449_n X 0.0232887f $X=9.35 $Y=3.56 $X2=0 $Y2=0
cc_348 N_VPWR_c_495_n N_X_c_599_n 0.0422929f $X=7.67 $Y=2.55 $X2=0 $Y2=0
cc_349 N_X_c_540_n N_VGND_c_646_n 0.0086879f $X=3.77 $Y=0.97 $X2=0 $Y2=0
cc_350 N_X_c_552_n N_VGND_c_648_n 0.0689585f $X=5.225 $Y=1.71 $X2=0 $Y2=0
cc_351 N_X_c_541_n N_VGND_c_649_n 0.0086879f $X=5.33 $Y=0.97 $X2=0 $Y2=0
cc_352 N_X_c_566_n N_VGND_c_650_n 0.0689585f $X=6.785 $Y=1.71 $X2=0 $Y2=0
cc_353 N_X_c_542_n N_VGND_c_651_n 0.0086879f $X=6.89 $Y=0.97 $X2=0 $Y2=0
cc_354 N_X_c_575_n N_VGND_c_652_n 0.0689585f $X=8.345 $Y=1.71 $X2=0 $Y2=0
cc_355 N_X_c_631_p N_VGND_c_653_n 0.00873551f $X=8.45 $Y=0.975 $X2=0 $Y2=0
cc_356 N_X_c_582_n N_VGND_c_653_n 0.0066386f $X=8.735 $Y=0.89 $X2=0 $Y2=0
cc_357 N_X_c_598_n N_VGND_c_653_n 0.0102128f $X=8.85 $Y=0.975 $X2=0 $Y2=0
cc_358 N_X_c_540_n N_VGND_c_655_n 0.00668507f $X=3.77 $Y=0.97 $X2=0 $Y2=0
cc_359 N_X_c_541_n N_VGND_c_655_n 0.00668507f $X=5.33 $Y=0.97 $X2=0 $Y2=0
cc_360 N_X_c_542_n N_VGND_c_655_n 0.00668507f $X=6.89 $Y=0.97 $X2=0 $Y2=0
cc_361 N_X_c_631_p N_VGND_c_655_n 0.00674935f $X=8.45 $Y=0.975 $X2=0 $Y2=0
cc_362 N_X_c_582_n N_VGND_c_655_n 0.00486341f $X=8.735 $Y=0.89 $X2=0 $Y2=0
cc_363 N_X_c_598_n N_VGND_c_655_n 0.00631558f $X=8.85 $Y=0.975 $X2=0 $Y2=0
