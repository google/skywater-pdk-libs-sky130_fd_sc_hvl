* File: sky130_fd_sc_hvl__dlrtp_1.pex.spice
* Created: Wed Sep  2 09:05:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%VNB 5 7 11 25
r71 7 25 1.30208e-05 $w=9.6e-06 $l=1e-09 $layer=MET1_cond $X=4.8 $Y=0.057
+ $X2=4.8 $Y2=0.058
r72 7 11 0.000742187 $w=9.6e-06 $l=5.7e-08 $layer=MET1_cond $X=4.8 $Y=0.057
+ $X2=4.8 $Y2=0
r73 5 11 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r74 5 11 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%VPB 4 6 14 21
c63 4 0 1.91513e-19 $X=-0.33 $Y=1.885
r64 10 21 0.000742187 $w=9.6e-06 $l=5.7e-08 $layer=MET1_cond $X=4.8 $Y=4.07
+ $X2=4.8 $Y2=4.013
r65 10 14 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=9.36 $Y=4.07
+ $X2=9.36 $Y2=4.07
r66 9 14 594.995 $w=1.68e-07 $l=9.12e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=9.36 $Y2=4.07
r67 9 10 0.93 $w=1.7e-07 $l=1.7e-06 $layer=mcon $count=10 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r68 6 21 1.30208e-05 $w=9.6e-06 $l=1e-09 $layer=MET1_cond $X=4.8 $Y=4.012
+ $X2=4.8 $Y2=4.013
r69 4 14 18.2 $w=1.7e-07 $l=9.4024e-06 $layer=licon1_NTAP_notbjt $count=10 $X=0
+ $Y=3.985 $X2=9.36 $Y2=4.07
r70 4 9 18.2 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=10 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%D 1 2 6 12
r19 9 12 117.706 $w=5e-07 $l=1.1e-06 $layer=POLY_cond $X=0.695 $Y=2.095
+ $X2=0.695 $Y2=3.195
r20 6 9 144.458 $w=5e-07 $l=1.35e-06 $layer=POLY_cond $X=0.695 $Y=0.745
+ $X2=0.695 $Y2=2.095
r21 1 2 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.735 $Y=2.035
+ $X2=0.735 $Y2=2.405
r22 1 9 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.735
+ $Y=2.095 $X2=0.735 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%GATE 1 2 3 8 14
c33 3 0 3.46739e-20 $X=1.68 $Y=1.295
r34 11 14 203.846 $w=5e-07 $l=1.905e-06 $layer=POLY_cond $X=1.475 $Y=1.29
+ $X2=1.475 $Y2=3.195
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.41
+ $Y=1.29 $X2=1.41 $Y2=1.29
r36 8 11 58.3182 $w=5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.475 $Y=0.745
+ $X2=1.475 $Y2=1.29
r37 3 12 13.8293 $w=2.23e-07 $l=2.7e-07 $layer=LI1_cond $X=1.68 $Y=1.287
+ $X2=1.41 $Y2=1.287
r38 2 12 10.7561 $w=2.23e-07 $l=2.1e-07 $layer=LI1_cond $X=1.2 $Y=1.287 $X2=1.41
+ $Y2=1.287
r39 1 2 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.287 $X2=1.2
+ $Y2=1.287
.ends

.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%A_345_107# 1 2 7 8 11 16 19 20 21 25 26 30
+ 34 35 38 42 46
c112 34 0 1.60823e-19 $X=4.27 $Y=1.77
c113 21 0 3.46739e-20 $X=2.03 $Y=2.11
c114 8 0 1.87959e-19 $X=4.585 $Y=1.68
r115 35 46 113.426 $w=5e-07 $l=1.06e-06 $layer=POLY_cond $X=4.335 $Y=1.77
+ $X2=4.335 $Y2=2.83
r116 34 36 8.99783 $w=4.61e-07 $l=3.4e-07 $layer=LI1_cond $X=4.135 $Y=1.77
+ $X2=4.135 $Y2=2.11
r117 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.27
+ $Y=1.77 $X2=4.27 $Y2=1.77
r118 28 30 4.66471 $w=4.98e-07 $l=1.95e-07 $layer=LI1_cond $X=1.865 $Y=0.745
+ $X2=2.06 $Y2=0.745
r119 25 34 9.52711 $w=4.61e-07 $l=4.87442e-07 $layer=LI1_cond $X=3.835 $Y=1.41
+ $X2=4.135 $Y2=1.77
r120 25 26 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=3.835 $Y=1.41
+ $X2=2.145 $Y2=1.41
r121 24 42 77.0442 $w=5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.845 $Y=2.11
+ $X2=2.845 $Y2=2.83
r122 24 38 146.063 $w=5e-07 $l=1.365e-06 $layer=POLY_cond $X=2.845 $Y=2.11
+ $X2=2.845 $Y2=0.745
r123 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.78
+ $Y=2.11 $X2=2.78 $Y2=2.11
r124 21 23 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.03 $Y=2.11
+ $X2=2.78 $Y2=2.11
r125 20 36 6.64987 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=3.835 $Y=2.11
+ $X2=4.135 $Y2=2.11
r126 20 23 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=3.835 $Y=2.11
+ $X2=2.78 $Y2=2.11
r127 19 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.06 $Y=1.325
+ $X2=2.145 $Y2=1.41
r128 18 30 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=2.06 $Y=0.995
+ $X2=2.06 $Y2=0.745
r129 18 19 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.06 $Y=0.995
+ $X2=2.06 $Y2=1.325
r130 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.865 $Y=2.195
+ $X2=2.03 $Y2=2.11
r131 14 16 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=1.865 $Y=2.195
+ $X2=1.865 $Y2=2.945
r132 13 35 1.60509 $w=5e-07 $l=1.5e-08 $layer=POLY_cond $X=4.335 $Y=1.755
+ $X2=4.335 $Y2=1.77
r133 9 11 92.0251 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.23 $Y=1.605 $X2=5.23
+ $Y2=0.745
r134 8 13 38.6381 $w=1.5e-07 $l=2.85044e-07 $layer=POLY_cond $X=4.585 $Y=1.68
+ $X2=4.335 $Y2=1.755
r135 7 9 38.6381 $w=1.5e-07 $l=2.85044e-07 $layer=POLY_cond $X=4.98 $Y=1.68
+ $X2=5.23 $Y2=1.605
r136 7 8 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.98 $Y=1.68
+ $X2=4.585 $Y2=1.68
r137 2 16 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.725
+ $Y=2.82 $X2=1.865 $Y2=2.945
r138 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.725
+ $Y=0.535 $X2=1.865 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%A_32_107# 1 2 9 13 17 21 23 27 28 30 31
c65 27 0 9.83206e-20 $X=3.49 $Y=1.76
r66 31 33 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.76
r67 28 37 18.3095 $w=5.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.59 $Y=1.76
+ $X2=3.59 $Y2=1.945
r68 28 36 30.512 $w=5.7e-07 $l=3.15e-07 $layer=POLY_cond $X=3.59 $Y=1.76
+ $X2=3.59 $Y2=1.445
r69 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.49
+ $Y=1.76 $X2=3.49 $Y2=1.76
r70 25 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=1.76
+ $X2=1.71 $Y2=1.76
r71 25 27 110.583 $w=1.68e-07 $l=1.695e-06 $layer=LI1_cond $X=1.795 $Y=1.76
+ $X2=3.49 $Y2=1.76
r72 24 30 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.39 $Y=1.665
+ $X2=0.265 $Y2=1.665
r73 23 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=1.665
+ $X2=1.71 $Y2=1.665
r74 23 24 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=1.625 $Y=1.665
+ $X2=0.39 $Y2=1.665
r75 19 30 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=1.75
+ $X2=0.265 $Y2=1.665
r76 19 21 55.0868 $w=2.48e-07 $l=1.195e-06 $layer=LI1_cond $X=0.265 $Y=1.75
+ $X2=0.265 $Y2=2.945
r77 15 30 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=1.58
+ $X2=0.265 $Y2=1.665
r78 15 17 38.4916 $w=2.48e-07 $l=8.35e-07 $layer=LI1_cond $X=0.265 $Y=1.58
+ $X2=0.265 $Y2=0.745
r79 13 37 94.7002 $w=5e-07 $l=8.85e-07 $layer=POLY_cond $X=3.625 $Y=2.83
+ $X2=3.625 $Y2=1.945
r80 9 36 74.9041 $w=5e-07 $l=7e-07 $layer=POLY_cond $X=3.625 $Y=0.745 $X2=3.625
+ $Y2=1.445
r81 2 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=2.82 $X2=0.305 $Y2=2.945
r82 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.535 $X2=0.305 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%A_462_107# 1 2 9 12 16 18 19 20 21 23 25 29
+ 30 33 39
c99 30 0 3.81261e-19 $X=5.01 $Y=2.13
c100 18 0 8.96383e-20 $X=4.185 $Y=1.06
r101 30 39 20.6903 $w=6.55e-07 $l=2.15e-07 $layer=POLY_cond $X=5.152 $Y=2.13
+ $X2=5.152 $Y2=2.345
r102 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.01
+ $Y=2.13 $X2=5.01 $Y2=2.13
r103 26 33 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.335 $Y=1.23
+ $X2=4.335 $Y2=0.745
r104 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.34
+ $Y=1.23 $X2=4.34 $Y2=1.23
r105 23 29 9.11628 $w=3.91e-07 $l=2.64953e-07 $layer=LI1_cond $X=4.7 $Y=1.965
+ $X2=4.895 $Y2=2.13
r106 22 25 14.689 $w=2.99e-07 $l=4.5299e-07 $layer=LI1_cond $X=4.7 $Y=1.395
+ $X2=4.34 $Y2=1.185
r107 22 23 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.7 $Y=1.395
+ $X2=4.7 $Y2=1.965
r108 20 29 10.2967 $w=3.91e-07 $l=4.48665e-07 $layer=LI1_cond $X=4.615 $Y=2.46
+ $X2=4.895 $Y2=2.13
r109 20 21 130.155 $w=1.68e-07 $l=1.995e-06 $layer=LI1_cond $X=4.615 $Y=2.46
+ $X2=2.62 $Y2=2.46
r110 18 25 8.57648 $w=2.99e-07 $l=2.08327e-07 $layer=LI1_cond $X=4.185 $Y=1.06
+ $X2=4.34 $Y2=1.185
r111 18 19 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=4.185 $Y=1.06
+ $X2=2.62 $Y2=1.06
r112 14 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.495 $Y=0.975
+ $X2=2.62 $Y2=1.06
r113 14 16 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=2.495 $Y=0.975
+ $X2=2.495 $Y2=0.745
r114 10 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.455 $Y=2.545
+ $X2=2.62 $Y2=2.46
r115 10 12 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.455 $Y=2.545
+ $X2=2.455 $Y2=2.58
r116 9 39 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.23 $Y=2.665 $X2=5.23
+ $Y2=2.345
r117 2 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.31
+ $Y=2.455 $X2=2.455 $Y2=2.58
r118 1 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.31
+ $Y=0.535 $X2=2.455 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%A_1138_81# 1 2 7 9 12 16 19 20 22 23 25 27
+ 30 36 40 44 49
c91 22 0 1.91513e-19 $X=7.045 $Y=1.905
c92 20 0 1.06401e-19 $X=6.14 $Y=1.99
r93 48 49 43.3374 $w=5e-07 $l=4.05e-07 $layer=POLY_cond $X=8.51 $Y=1.855
+ $X2=8.915 $Y2=1.855
r94 37 48 4.81527 $w=5e-07 $l=4.5e-08 $layer=POLY_cond $X=8.465 $Y=1.855
+ $X2=8.51 $Y2=1.855
r95 36 38 13.2509 $w=2.67e-07 $l=2.9e-07 $layer=LI1_cond $X=8.465 $Y=1.83
+ $X2=8.465 $Y2=2.12
r96 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.465
+ $Y=1.83 $X2=8.465 $Y2=1.83
r97 30 32 11.1667 $w=3.73e-07 $l=2.5e-07 $layer=LI1_cond $X=6.942 $Y=0.745
+ $X2=6.942 $Y2=0.995
r98 28 34 4.38581 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=7.39 $Y=2.12
+ $X2=7.175 $Y2=2.12
r99 27 38 3.37873 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.3 $Y=2.12
+ $X2=8.465 $Y2=2.12
r100 27 28 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=8.3 $Y=2.12 $X2=7.39
+ $Y2=2.12
r101 23 34 3.27848 $w=4.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.175 $Y=2.205
+ $X2=7.175 $Y2=2.12
r102 23 25 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=7.175 $Y=2.205
+ $X2=7.175 $Y2=2.34
r103 22 32 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=7.045 $Y=1.905
+ $X2=7.045 $Y2=0.995
r104 19 34 5.00315 $w=3.17e-07 $l=2.72351e-07 $layer=LI1_cond $X=6.96 $Y=1.99
+ $X2=7.175 $Y2=2.12
r105 19 22 5.87851 $w=3.17e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.96 $Y=1.99
+ $X2=7.045 $Y2=1.905
r106 19 20 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=6.96 $Y=1.99
+ $X2=6.14 $Y2=1.99
r107 17 44 110.751 $w=5e-07 $l=1.035e-06 $layer=POLY_cond $X=5.94 $Y=1.63
+ $X2=5.94 $Y2=2.665
r108 17 40 94.7002 $w=5e-07 $l=8.85e-07 $layer=POLY_cond $X=5.94 $Y=1.63
+ $X2=5.94 $Y2=0.745
r109 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.975
+ $Y=1.63 $X2=5.975 $Y2=1.63
r110 14 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.975 $Y=1.905
+ $X2=6.14 $Y2=1.99
r111 14 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.975 $Y=1.905
+ $X2=5.975 $Y2=1.63
r112 10 49 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.915 $Y=1.605
+ $X2=8.915 $Y2=1.855
r113 10 12 74.3691 $w=5e-07 $l=6.95e-07 $layer=POLY_cond $X=8.915 $Y=1.605
+ $X2=8.915 $Y2=0.91
r114 7 48 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.51 $Y=2.105 $X2=8.51
+ $Y2=1.855
r115 7 9 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.51 $Y=2.105 $X2=8.51
+ $Y2=2.965
r116 2 25 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=7.085
+ $Y=2.215 $X2=7.225 $Y2=2.34
r117 1 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.775
+ $Y=0.535 $X2=6.92 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%A_917_107# 1 2 9 11 13 14 17 18 20 21 22 24
+ 25 32 34 36 39
c105 22 0 1.14037e-19 $X=5.135 $Y=1.26
r106 37 39 18.7019 $w=5.67e-07 $l=2.2e-07 $layer=POLY_cond $X=6.615 $Y=1.435
+ $X2=6.835 $Y2=1.435
r107 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.615
+ $Y=1.28 $X2=6.615 $Y2=1.28
r108 30 32 5.02353 $w=4.98e-07 $l=2.1e-07 $layer=LI1_cond $X=4.84 $Y=0.745
+ $X2=5.05 $Y2=0.745
r109 26 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.525 $Y=1.26
+ $X2=5.44 $Y2=1.26
r110 25 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.45 $Y=1.26
+ $X2=6.615 $Y2=1.26
r111 25 26 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=6.45 $Y=1.26
+ $X2=5.525 $Y2=1.26
r112 23 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=1.345
+ $X2=5.44 $Y2=1.26
r113 23 24 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.44 $Y=1.345
+ $X2=5.44 $Y2=2.725
r114 21 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.355 $Y=1.26
+ $X2=5.44 $Y2=1.26
r115 21 22 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.355 $Y=1.26
+ $X2=5.135 $Y2=1.26
r116 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.05 $Y=1.175
+ $X2=5.135 $Y2=1.26
r117 19 32 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=5.05 $Y=0.995
+ $X2=5.05 $Y2=0.745
r118 19 20 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.05 $Y=0.995
+ $X2=5.05 $Y2=1.175
r119 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.355 $Y=2.81
+ $X2=5.44 $Y2=2.725
r120 17 18 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=5.355 $Y=2.81
+ $X2=4.89 $Y2=2.81
r121 14 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.725 $Y=2.895
+ $X2=4.89 $Y2=2.81
r122 14 16 1.84848 $w=3.3e-07 $l=5e-08 $layer=LI1_cond $X=4.725 $Y=2.895
+ $X2=4.725 $Y2=2.945
r123 11 39 40.3792 $w=5.67e-07 $l=6.33542e-07 $layer=POLY_cond $X=7.31 $Y=1.065
+ $X2=6.835 $Y2=1.435
r124 11 13 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.31 $Y=1.065 $X2=7.31
+ $Y2=0.745
r125 7 39 5.81687 $w=5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.835 $Y=1.805
+ $X2=6.835 $Y2=1.435
r126 7 9 83.9996 $w=5e-07 $l=7.85e-07 $layer=POLY_cond $X=6.835 $Y=1.805
+ $X2=6.835 $Y2=2.59
r127 2 16 600 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=1 $X=4.585
+ $Y=2.455 $X2=4.725 $Y2=2.945
r128 1 30 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=4.585
+ $Y=0.535 $X2=4.84 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%RESET_B 1 2 3 8 12 15
r35 15 18 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=8.02 $Y=0.745
+ $X2=8.02 $Y2=1.23
r36 8 12 87.7448 $w=5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.615 $Y=1.77 $X2=7.615
+ $Y2=2.59
r37 8 9 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.68 $Y=1.77
+ $X2=7.68 $Y2=1.77
r38 3 9 2.32909 $w=5.5e-07 $l=1.05e-07 $layer=LI1_cond $X=7.817 $Y=1.665
+ $X2=7.817 $Y2=1.77
r39 3 21 3.89602 $w=6.05e-07 $l=1.87e-07 $layer=LI1_cond $X=7.817 $Y=1.665
+ $X2=7.817 $Y2=1.478
r40 2 21 4.90293 $w=6.03e-07 $l=2.48e-07 $layer=LI1_cond $X=7.817 $Y=1.23
+ $X2=7.817 $Y2=1.478
r41 2 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.955
+ $Y=1.23 $X2=7.955 $Y2=1.23
r42 1 2 6.02982 $w=6.03e-07 $l=3.05e-07 $layer=LI1_cond $X=7.817 $Y=0.925
+ $X2=7.817 $Y2=1.23
.ends

.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%VPWR 1 2 3 4 13 16 25 34 43 51
r60 49 51 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.685 $Y=3.63
+ $X2=8.405 $Y2=3.63
r61 48 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.405 $Y=3.59
+ $X2=8.405 $Y2=3.59
r62 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.685 $Y=3.59
+ $X2=7.685 $Y2=3.59
r63 46 48 4.75158 $w=9.48e-07 $l=3.7e-07 $layer=LI1_cond $X=8.045 $Y=3.22
+ $X2=8.045 $Y2=3.59
r64 43 46 9.63158 $w=9.48e-07 $l=7.5e-07 $layer=LI1_cond $X=8.045 $Y=2.47
+ $X2=8.045 $Y2=3.22
r65 40 49 0.439572 $w=3.7e-07 $l=1.145e-06 $layer=MET1_cond $X=6.54 $Y=3.63
+ $X2=7.685 $Y2=3.63
r66 38 40 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.82 $Y=3.63
+ $X2=6.54 $Y2=3.63
r67 37 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.54 $Y=3.59
+ $X2=6.54 $Y2=3.59
r68 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.82 $Y=3.59
+ $X2=5.82 $Y2=3.59
r69 34 37 16.0526 $w=9.48e-07 $l=1.25e-06 $layer=LI1_cond $X=6.18 $Y=2.34
+ $X2=6.18 $Y2=3.59
r70 29 31 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.915 $Y=3.63
+ $X2=3.635 $Y2=3.63
r71 28 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.635 $Y=3.59
+ $X2=3.635 $Y2=3.59
r72 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.915 $Y=3.59
+ $X2=2.915 $Y2=3.59
r73 25 28 8.28316 $w=9.48e-07 $l=6.45e-07 $layer=LI1_cond $X=3.275 $Y=2.945
+ $X2=3.275 $Y2=3.59
r74 22 29 0.579697 $w=3.7e-07 $l=1.51e-06 $layer=MET1_cond $X=1.405 $Y=3.63
+ $X2=2.915 $Y2=3.63
r75 20 22 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.685 $Y=3.63
+ $X2=1.405 $Y2=3.63
r76 19 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.405 $Y=3.59
+ $X2=1.405 $Y2=3.59
r77 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.685 $Y=3.59
+ $X2=0.685 $Y2=3.59
r78 16 19 8.28316 $w=9.48e-07 $l=6.45e-07 $layer=LI1_cond $X=1.045 $Y=2.945
+ $X2=1.045 $Y2=3.59
r79 13 38 0.391584 $w=3.7e-07 $l=1.02e-06 $layer=MET1_cond $X=4.8 $Y=3.63
+ $X2=5.82 $Y2=3.63
r80 13 31 0.44725 $w=3.7e-07 $l=1.165e-06 $layer=MET1_cond $X=4.8 $Y=3.63
+ $X2=3.635 $Y2=3.63
r81 4 46 300 $w=1.7e-07 $l=1.1253e-06 $layer=licon1_PDIFF $count=2 $X=7.865
+ $Y=2.215 $X2=8.12 $Y2=3.22
r82 4 43 300 $w=1.7e-07 $l=3.60624e-07 $layer=licon1_PDIFF $count=2 $X=7.865
+ $Y=2.215 $X2=8.12 $Y2=2.47
r83 3 34 300 $w=1.7e-07 $l=3.07164e-07 $layer=licon1_PDIFF $count=2 $X=6.19
+ $Y=2.455 $X2=6.445 $Y2=2.34
r84 2 25 600 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=2.455 $X2=3.235 $Y2=2.945
r85 1 16 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.945
+ $Y=2.82 $X2=1.085 $Y2=2.945
.ends

.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%Q 1 2 7 8 9 10 11 12 13 23 42
r19 42 43 6.29164 $w=7.38e-07 $l=1.65e-07 $layer=LI1_cond $X=9.105 $Y=2.34
+ $X2=9.105 $Y2=2.175
r20 13 39 7.19263 $w=7.38e-07 $l=4.45e-07 $layer=LI1_cond $X=9.105 $Y=3.145
+ $X2=9.105 $Y2=3.59
r21 12 13 5.98039 $w=7.38e-07 $l=3.7e-07 $layer=LI1_cond $X=9.105 $Y=2.775
+ $X2=9.105 $Y2=3.145
r22 12 33 3.71754 $w=7.38e-07 $l=2.3e-07 $layer=LI1_cond $X=9.105 $Y=2.775
+ $X2=9.105 $Y2=2.545
r23 11 33 2.26285 $w=7.38e-07 $l=1.4e-07 $layer=LI1_cond $X=9.105 $Y=2.405
+ $X2=9.105 $Y2=2.545
r24 11 42 1.05061 $w=7.38e-07 $l=6.5e-08 $layer=LI1_cond $X=9.105 $Y=2.405
+ $X2=9.105 $Y2=2.34
r25 10 43 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=9.307 $Y=2.035
+ $X2=9.307 $Y2=2.175
r26 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=9.307 $Y=1.665
+ $X2=9.307 $Y2=2.035
r27 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=9.307 $Y=1.295
+ $X2=9.307 $Y2=1.665
r28 7 8 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=9.307 $Y=0.925
+ $X2=9.307 $Y2=1.295
r29 7 23 9.11634 $w=3.33e-07 $l=2.65e-07 $layer=LI1_cond $X=9.307 $Y=0.925
+ $X2=9.307 $Y2=0.66
r30 2 42 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=8.76
+ $Y=2.215 $X2=8.9 $Y2=2.34
r31 2 39 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=8.76
+ $Y=2.215 $X2=8.9 $Y2=3.59
r32 1 23 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=9.165
+ $Y=0.535 $X2=9.305 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__DLRTP_1%VGND 1 2 3 4 13 16 25 40 44 45
r68 48 50 10.1363 $w=5.88e-07 $l=5e-07 $layer=LI1_cond $X=8.595 $Y=0.66
+ $X2=8.595 $Y2=1.16
r69 44 48 3.64905 $w=5.88e-07 $l=1.8e-07 $layer=LI1_cond $X=8.595 $Y=0.48
+ $X2=8.595 $Y2=0.66
r70 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.775 $Y=0.48
+ $X2=8.775 $Y2=0.48
r71 41 45 0.919453 $w=3.7e-07 $l=2.395e-06 $layer=MET1_cond $X=6.38 $Y=0.44
+ $X2=8.775 $Y2=0.44
r72 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.38 $Y=0.48
+ $X2=6.38 $Y2=0.48
r73 38 40 0.949269 $w=6.28e-07 $l=5e-08 $layer=LI1_cond $X=6.33 $Y=0.68 $X2=6.38
+ $Y2=0.68
r74 35 41 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.66 $Y=0.44
+ $X2=6.38 $Y2=0.44
r75 34 38 12.7202 $w=6.28e-07 $l=6.7e-07 $layer=LI1_cond $X=5.66 $Y=0.68
+ $X2=6.33 $Y2=0.68
r76 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.66 $Y=0.48
+ $X2=5.66 $Y2=0.48
r77 26 29 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.915 $Y=0.44
+ $X2=3.635 $Y2=0.44
r78 25 31 2.63263 $w=9.48e-07 $l=2.05e-07 $layer=LI1_cond $X=3.275 $Y=0.48
+ $X2=3.275 $Y2=0.685
r79 25 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.635 $Y=0.48
+ $X2=3.635 $Y2=0.48
r80 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.915 $Y=0.48
+ $X2=2.915 $Y2=0.48
r81 20 26 0.579697 $w=3.7e-07 $l=1.51e-06 $layer=MET1_cond $X=1.405 $Y=0.44
+ $X2=2.915 $Y2=0.44
r82 17 20 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.685 $Y=0.44
+ $X2=1.405 $Y2=0.44
r83 16 22 3.40316 $w=9.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.045 $Y=0.48
+ $X2=1.045 $Y2=0.745
r84 16 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.405 $Y=0.48
+ $X2=1.405 $Y2=0.48
r85 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.685 $Y=0.48
+ $X2=0.685 $Y2=0.48
r86 13 35 0.330159 $w=3.7e-07 $l=8.6e-07 $layer=MET1_cond $X=4.8 $Y=0.44
+ $X2=5.66 $Y2=0.44
r87 13 29 0.44725 $w=3.7e-07 $l=1.165e-06 $layer=MET1_cond $X=4.8 $Y=0.44
+ $X2=3.635 $Y2=0.44
r88 4 50 182 $w=1.7e-07 $l=7.4162e-07 $layer=licon1_NDIFF $count=1 $X=8.27
+ $Y=0.535 $X2=8.525 $Y2=1.16
r89 4 48 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=8.27
+ $Y=0.535 $X2=8.525 $Y2=0.66
r90 3 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.19
+ $Y=0.535 $X2=6.33 $Y2=0.745
r91 2 31 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=3.095
+ $Y=0.535 $X2=3.235 $Y2=0.685
r92 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.945
+ $Y=0.535 $X2=1.085 $Y2=0.745
.ends

