# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__sdfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  19.20000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.910000 2.660000 3.205000 3.260000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.820000 0.515000 19.075000 3.755000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  4.415000 2.290000  4.705000 2.335000 ;
        RECT  4.415000 2.335000 14.305000 2.475000 ;
        RECT  4.415000 2.475000  4.705000 2.520000 ;
        RECT  8.255000 2.290000  8.545000 2.335000 ;
        RECT  8.255000 2.475000  8.545000 2.520000 ;
        RECT 14.015000 2.290000 14.305000 2.335000 ;
        RECT 14.015000 2.475000 14.305000 2.520000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 1.115000 1.510000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.445000 2.245000 1.835000 ;
        RECT 1.995000 1.835000 3.175000 2.005000 ;
        RECT 1.995000 2.005000 2.380000 2.575000 ;
        RECT 3.005000 1.550000 5.635000 1.835000 ;
        RECT 4.880000 1.835000 5.635000 2.525000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 15.485000 1.955000 16.140000 2.495000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 19.200000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 19.200000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 19.200000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 19.200000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 19.530000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 19.200000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 19.200000 0.085000 ;
      RECT  0.000000  3.985000 19.200000 4.155000 ;
      RECT  0.305000  1.690000  1.465000 1.860000 ;
      RECT  0.305000  1.860000  0.475000 3.105000 ;
      RECT  0.305000  3.105000  2.730000 3.275000 ;
      RECT  0.305000  3.275000  0.635000 3.705000 ;
      RECT  0.665000  0.265000  3.975000 0.435000 ;
      RECT  0.665000  0.435000  0.995000 0.995000 ;
      RECT  0.730000  2.255000  1.060000 2.755000 ;
      RECT  0.730000  2.755000  2.730000 2.925000 ;
      RECT  1.295000  0.615000  2.485000 0.915000 ;
      RECT  1.295000  0.915000  1.465000 1.690000 ;
      RECT  1.420000  3.455000  2.370000 3.705000 ;
      RECT  1.645000  1.095000  2.810000 1.175000 ;
      RECT  1.645000  1.175000  5.535000 1.265000 ;
      RECT  1.645000  1.265000  1.815000 2.755000 ;
      RECT  2.480000  1.265000  5.535000 1.345000 ;
      RECT  2.480000  1.345000  2.810000 1.655000 ;
      RECT  2.560000  2.310000  3.555000 2.480000 ;
      RECT  2.560000  2.480000  2.730000 2.755000 ;
      RECT  2.560000  3.275000  2.730000 3.535000 ;
      RECT  2.560000  3.535000  3.555000 3.705000 ;
      RECT  3.385000  2.480000  3.555000 2.705000 ;
      RECT  3.385000  2.705000  5.485000 2.875000 ;
      RECT  3.385000  3.055000  4.975000 3.225000 ;
      RECT  3.385000  3.225000  3.555000 3.535000 ;
      RECT  3.645000  0.435000  3.975000 0.995000 ;
      RECT  3.735000  3.405000  4.625000 3.705000 ;
      RECT  3.965000  2.015000  4.300000 2.290000 ;
      RECT  3.965000  2.290000  4.675000 2.525000 ;
      RECT  4.155000  0.365000  5.105000 0.995000 ;
      RECT  4.805000  3.225000  4.975000 3.635000 ;
      RECT  4.805000  3.635000  6.005000 3.805000 ;
      RECT  5.155000  2.875000  5.485000 3.455000 ;
      RECT  5.285000  0.515000  5.535000 1.175000 ;
      RECT  5.755000  0.515000  6.005000 1.005000 ;
      RECT  5.755000  3.165000  6.005000 3.635000 ;
      RECT  5.835000  1.005000  6.005000 3.165000 ;
      RECT  6.185000  0.265000  7.255000 0.435000 ;
      RECT  6.185000  0.435000  6.355000 3.635000 ;
      RECT  6.185000  3.635000  7.215000 3.805000 ;
      RECT  6.535000  0.615000  6.865000 0.995000 ;
      RECT  6.535000  0.995000  6.705000 2.715000 ;
      RECT  6.535000  2.715000  9.215000 2.885000 ;
      RECT  6.535000  2.885000  6.865000 3.455000 ;
      RECT  6.950000  1.915000  7.605000 2.085000 ;
      RECT  6.950000  2.085000  7.280000 2.535000 ;
      RECT  7.045000  0.435000  7.255000 1.175000 ;
      RECT  7.045000  1.175000  9.635000 1.345000 ;
      RECT  7.045000  1.345000  7.255000 1.735000 ;
      RECT  7.045000  3.065000  8.705000 3.235000 ;
      RECT  7.045000  3.235000  7.215000 3.635000 ;
      RECT  7.405000  3.415000  8.355000 3.705000 ;
      RECT  7.435000  1.525000 10.780000 1.695000 ;
      RECT  7.435000  1.695000  7.605000 1.915000 ;
      RECT  7.785000  1.875000 11.130000 2.045000 ;
      RECT  7.785000  2.045000  8.115000 2.535000 ;
      RECT  8.115000  0.365000  9.065000 0.995000 ;
      RECT  8.295000  2.225000  8.760000 2.535000 ;
      RECT  8.535000  3.235000  8.705000 3.635000 ;
      RECT  8.535000  3.635000  9.785000 3.805000 ;
      RECT  8.885000  2.885000  9.215000 3.455000 ;
      RECT  9.045000  2.225000 10.780000 2.395000 ;
      RECT  9.045000  2.395000  9.215000 2.715000 ;
      RECT  9.305000  0.885000  9.635000 1.175000 ;
      RECT  9.455000  2.695000  9.785000 3.135000 ;
      RECT  9.455000  3.135000 12.810000 3.305000 ;
      RECT  9.455000  3.305000  9.785000 3.635000 ;
      RECT  9.840000  0.365000 10.430000 1.345000 ;
      RECT  9.965000  3.485000 10.915000 3.735000 ;
      RECT 10.490000  2.395000 10.780000 2.555000 ;
      RECT 10.610000  0.265000 12.455000 0.435000 ;
      RECT 10.610000  0.435000 10.780000 1.525000 ;
      RECT 10.960000  0.615000 11.325000 1.285000 ;
      RECT 10.960000  1.285000 11.130000 1.875000 ;
      RECT 10.960000  2.045000 11.130000 2.675000 ;
      RECT 10.960000  2.675000 11.440000 2.955000 ;
      RECT 11.310000  1.465000 11.480000 2.285000 ;
      RECT 11.310000  2.285000 11.790000 2.455000 ;
      RECT 11.620000  2.455000 11.790000 3.135000 ;
      RECT 11.660000  0.615000 12.105000 1.365000 ;
      RECT 11.660000  1.365000 11.830000 1.935000 ;
      RECT 11.660000  1.935000 13.200000 2.105000 ;
      RECT 11.970000  2.105000 12.300000 2.955000 ;
      RECT 12.010000  1.545000 14.395000 1.715000 ;
      RECT 12.010000  1.715000 13.020000 1.755000 ;
      RECT 12.285000  0.435000 12.455000 1.545000 ;
      RECT 12.480000  2.285000 12.810000 3.135000 ;
      RECT 13.015000  3.370000 13.965000 3.705000 ;
      RECT 13.030000  2.105000 13.200000 3.020000 ;
      RECT 13.030000  3.020000 14.315000 3.190000 ;
      RECT 13.085000  0.365000 14.035000 1.365000 ;
      RECT 13.380000  1.895000 13.710000 2.670000 ;
      RECT 13.380000  2.670000 14.745000 2.840000 ;
      RECT 14.040000  1.895000 14.370000 2.490000 ;
      RECT 14.145000  3.190000 14.315000 3.355000 ;
      RECT 14.145000  3.355000 15.095000 3.525000 ;
      RECT 14.225000  0.535000 16.085000 0.705000 ;
      RECT 14.225000  0.705000 14.395000 1.545000 ;
      RECT 14.495000  2.840000 14.745000 3.175000 ;
      RECT 14.575000  1.175000 15.535000 1.345000 ;
      RECT 14.575000  1.345000 14.745000 2.670000 ;
      RECT 14.925000  1.605000 16.850000 1.775000 ;
      RECT 14.925000  1.775000 15.255000 2.275000 ;
      RECT 14.925000  2.275000 15.095000 3.355000 ;
      RECT 15.205000  0.885000 15.535000 1.175000 ;
      RECT 15.275000  2.675000 16.165000 3.705000 ;
      RECT 15.755000  0.705000 16.085000 1.255000 ;
      RECT 15.755000  1.255000 17.200000 1.425000 ;
      RECT 16.275000  0.365000 16.865000 0.995000 ;
      RECT 16.345000  1.955000 17.200000 2.125000 ;
      RECT 16.345000  2.125000 16.595000 3.505000 ;
      RECT 17.030000  1.425000 17.200000 1.955000 ;
      RECT 17.065000  2.305000 17.550000 3.005000 ;
      RECT 17.105000  0.825000 17.550000 1.075000 ;
      RECT 17.380000  1.075000 17.550000 1.485000 ;
      RECT 17.380000  1.485000 18.615000 1.815000 ;
      RECT 17.380000  1.815000 17.550000 2.305000 ;
      RECT 17.730000  0.365000 18.640000 1.305000 ;
      RECT 17.730000  2.175000 18.640000 3.755000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.450000  3.505000  1.620000 3.675000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  1.810000  3.505000  1.980000 3.675000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.170000  3.505000  2.340000 3.675000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.735000  3.505000  3.905000 3.675000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.095000  3.505000  4.265000 3.675000 ;
      RECT  4.185000  0.395000  4.355000 0.565000 ;
      RECT  4.455000  3.505000  4.625000 3.675000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  2.320000  4.645000 2.490000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.545000  0.395000  4.715000 0.565000 ;
      RECT  4.905000  0.395000  5.075000 0.565000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.435000  3.505000  7.605000 3.675000 ;
      RECT  7.795000  3.505000  7.965000 3.675000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.145000  0.395000  8.315000 0.565000 ;
      RECT  8.155000  3.505000  8.325000 3.675000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  2.320000  8.485000 2.490000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.505000  0.395000  8.675000 0.565000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.865000  0.395000  9.035000 0.565000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.870000  0.395000 10.040000 0.565000 ;
      RECT  9.995000  3.515000 10.165000 3.685000 ;
      RECT 10.230000  0.395000 10.400000 0.565000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.355000  3.515000 10.525000 3.685000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.515000 10.885000 3.685000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 13.045000  3.505000 13.215000 3.675000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  0.395000 13.285000 0.565000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.405000  3.505000 13.575000 3.675000 ;
      RECT 13.475000  0.395000 13.645000 0.565000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.765000  3.505000 13.935000 3.675000 ;
      RECT 13.835000  0.395000 14.005000 0.565000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  2.320000 14.245000 2.490000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.275000  3.505000 15.445000 3.675000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.635000  3.505000 15.805000 3.675000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.505000 16.165000 3.675000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.305000  0.395000 16.475000 0.565000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.665000  0.395000 16.835000 0.565000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
      RECT 17.740000  0.395000 17.910000 0.565000 ;
      RECT 17.740000  3.505000 17.910000 3.675000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.985000 18.085000 4.155000 ;
      RECT 18.100000  0.395000 18.270000 0.565000 ;
      RECT 18.100000  3.505000 18.270000 3.675000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.985000 18.565000 4.155000 ;
      RECT 18.460000  0.395000 18.630000 0.565000 ;
      RECT 18.460000  3.505000 18.630000 3.675000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  3.985000 19.045000 4.155000 ;
  END
END sky130_fd_sc_hvl__sdfrtp_1
END LIBRARY
