* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_87_81# B2 a_533_443# VPB phv w=1.5e+06u l=500000u
+  ad=4.2e+11p pd=3.56e+06u as=3.15e+11p ps=3.42e+06u
M1001 VGND A2 a_354_107# VNB nhv w=750000u l=500000u
+  ad=4.65e+11p pd=4.24e+06u as=4.2e+11p ps=4.12e+06u
M1002 a_87_81# B1 a_354_107# VNB nhv w=750000u l=500000u
+  ad=2.4375e+11p pd=2.15e+06u as=0p ps=0u
M1003 VGND a_87_81# X VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=2.1375e+11p ps=2.07e+06u
M1004 a_354_107# B2 a_87_81# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_831_443# A2 a_87_81# VPB phv w=1.5e+06u l=500000u
+  ad=3.15e+11p pd=3.42e+06u as=0p ps=0u
M1006 VPWR A1 a_831_443# VPB phv w=1.5e+06u l=500000u
+  ad=2.2425e+12p pd=8.99e+06u as=0p ps=0u
M1007 a_354_107# A1 VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_87_81# X VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=4.275e+11p ps=3.57e+06u
M1009 a_533_443# B1 VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
