* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hvl__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
*.PININFO A0:I A1:I A2:I A3:I S0:I S1:I VGND:I VNB:I VPB:I VPWR:I X:O
MMNA00 sndNS0ba0 S0b VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMNA01 VGND A0 VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMNA10 sndNS0a1 S0 VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMNA11 VGND A1 VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMNA20 sndNS0ba2 S0b VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMNA21 VGND A2 VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMNA30 sndNS0a3 S0 VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMNA31 VGND A3 VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMNs1o xb S1b VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMNs2o xb S1 VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.028 perim=0.76
MMIN1 VGND S1 VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMIN2 VGND S0 VNB nhv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMIN4 VGND xb VNB nhv m=1 w=0.75 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMPA00 sndPA0a0 A0 VPB phv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMPA01 xlowb S0 VPB phv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMPA10 sndPA1a1 A1 VPB phv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMPA11 xlowb S0b VPB phv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMPA20 sndPA2a2 A2 VPB phv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMPA21 xhib S0 VPB phv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMPA30 sndPA3a3 A3 VPB phv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMPA31 xhib S0b VPB phv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMPs1o xb S1 VPB phv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.028 perim=0.76
MMPs2o xb S1b VPB phv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMIP1 VPWR S1 VPB phv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMIP2 VPWR S0 VPB phv m=1 w=0.42 l=0.5 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.028 perim=0.76
MMIP4 VPWR xb VPB phv m=1 w=1.5 l=0.5 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.028 perim=0.76
.ENDS sky130_fd_sc_hvl__mux4_1
