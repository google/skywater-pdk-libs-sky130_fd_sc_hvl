* File: sky130_fd_sc_hvl__dfxtp_1.pxi.spice
* Created: Wed Sep  2 09:05:34 2020
* 
x_PM_SKY130_FD_SC_HVL__DFXTP_1%VNB N_VNB_M1022_b VNB N_VNB_c_3_p VNB
+ PM_SKY130_FD_SC_HVL__DFXTP_1%VNB
x_PM_SKY130_FD_SC_HVL__DFXTP_1%VPB N_VPB_M1011_b VPB N_VPB_c_90_p VPB
+ PM_SKY130_FD_SC_HVL__DFXTP_1%VPB
x_PM_SKY130_FD_SC_HVL__DFXTP_1%CLK N_CLK_M1011_g N_CLK_M1022_g N_CLK_c_196_n
+ N_CLK_c_197_n N_CLK_c_203_n CLK CLK N_CLK_c_199_n
+ PM_SKY130_FD_SC_HVL__DFXTP_1%CLK
x_PM_SKY130_FD_SC_HVL__DFXTP_1%A_30_127# N_A_30_127#_M1022_s N_A_30_127#_M1011_s
+ N_A_30_127#_c_243_n N_A_30_127#_M1001_g N_A_30_127#_M1004_g
+ N_A_30_127#_M1013_g N_A_30_127#_c_229_n N_A_30_127#_M1000_g
+ N_A_30_127#_c_230_n N_A_30_127#_M1020_g N_A_30_127#_c_231_n
+ N_A_30_127#_c_232_n N_A_30_127#_M1002_g N_A_30_127#_c_235_n
+ N_A_30_127#_c_236_n N_A_30_127#_c_238_n N_A_30_127#_c_239_n
+ N_A_30_127#_c_286_p N_A_30_127#_c_272_n N_A_30_127#_c_257_n
+ N_A_30_127#_c_240_n N_A_30_127#_c_281_p N_A_30_127#_c_336_p
+ N_A_30_127#_c_259_n N_A_30_127#_c_323_p N_A_30_127#_c_241_n
+ N_A_30_127#_c_242_n N_A_30_127#_c_261_n N_A_30_127#_c_343_p
+ PM_SKY130_FD_SC_HVL__DFXTP_1%A_30_127#
x_PM_SKY130_FD_SC_HVL__DFXTP_1%D N_D_c_416_n N_D_M1017_g N_D_M1016_g N_D_c_424_n
+ D D N_D_c_419_n N_D_c_420_n PM_SKY130_FD_SC_HVL__DFXTP_1%D
x_PM_SKY130_FD_SC_HVL__DFXTP_1%A_339_559# N_A_339_559#_M1004_d
+ N_A_339_559#_M1001_d N_A_339_559#_c_490_n N_A_339_559#_M1014_g
+ N_A_339_559#_c_491_n N_A_339_559#_c_472_n N_A_339_559#_c_494_n
+ N_A_339_559#_c_495_n N_A_339_559#_c_474_n N_A_339_559#_c_475_n
+ N_A_339_559#_c_566_n N_A_339_559#_c_496_n N_A_339_559#_c_499_n
+ N_A_339_559#_c_528_n N_A_339_559#_c_476_n N_A_339_559#_c_478_n
+ N_A_339_559#_c_532_n N_A_339_559#_c_502_n N_A_339_559#_c_504_n
+ N_A_339_559#_c_542_n N_A_339_559#_c_480_n N_A_339_559#_c_580_p
+ N_A_339_559#_c_481_n N_A_339_559#_c_483_n N_A_339_559#_c_543_n
+ N_A_339_559#_c_485_n N_A_339_559#_c_506_n N_A_339_559#_c_507_n
+ N_A_339_559#_c_508_n N_A_339_559#_c_486_n N_A_339_559#_c_551_n
+ N_A_339_559#_M1012_g N_A_339_559#_M1005_g N_A_339_559#_M1010_g
+ PM_SKY130_FD_SC_HVL__DFXTP_1%A_339_559#
x_PM_SKY130_FD_SC_HVL__DFXTP_1%A_1024_371# N_A_1024_371#_M1021_d
+ N_A_1024_371#_M1003_d N_A_1024_371#_M1006_g N_A_1024_371#_M1007_g
+ N_A_1024_371#_c_690_n N_A_1024_371#_c_703_n N_A_1024_371#_c_691_n
+ N_A_1024_371#_c_696_n N_A_1024_371#_c_709_n N_A_1024_371#_c_692_n
+ N_A_1024_371#_c_693_n PM_SKY130_FD_SC_HVL__DFXTP_1%A_1024_371#
x_PM_SKY130_FD_SC_HVL__DFXTP_1%A_780_574# N_A_780_574#_M1013_d
+ N_A_780_574#_M1012_d N_A_780_574#_M1003_g N_A_780_574#_c_758_n
+ N_A_780_574#_M1021_g N_A_780_574#_c_760_n N_A_780_574#_c_761_n
+ N_A_780_574#_c_768_n N_A_780_574#_c_762_n N_A_780_574#_c_763_n
+ PM_SKY130_FD_SC_HVL__DFXTP_1%A_780_574#
x_PM_SKY130_FD_SC_HVL__DFXTP_1%A_1729_87# N_A_1729_87#_M1019_d
+ N_A_1729_87#_M1018_d N_A_1729_87#_M1008_g N_A_1729_87#_M1015_g
+ N_A_1729_87#_M1023_g N_A_1729_87#_M1009_g N_A_1729_87#_c_871_p
+ N_A_1729_87#_c_860_p N_A_1729_87#_c_834_n N_A_1729_87#_c_835_n
+ N_A_1729_87#_c_837_n N_A_1729_87#_c_845_n N_A_1729_87#_c_888_p
+ N_A_1729_87#_c_838_n N_A_1729_87#_c_839_n N_A_1729_87#_c_840_n
+ PM_SKY130_FD_SC_HVL__DFXTP_1%A_1729_87#
x_PM_SKY130_FD_SC_HVL__DFXTP_1%A_1455_543# N_A_1455_543#_M1010_d
+ N_A_1455_543#_M1020_d N_A_1455_543#_M1019_g N_A_1455_543#_c_911_n
+ N_A_1455_543#_M1018_g N_A_1455_543#_c_920_n N_A_1455_543#_c_921_n
+ N_A_1455_543#_c_912_n N_A_1455_543#_c_924_n N_A_1455_543#_c_913_n
+ N_A_1455_543#_c_947_n N_A_1455_543#_c_926_n N_A_1455_543#_c_978_n
+ N_A_1455_543#_c_914_n N_A_1455_543#_c_953_n
+ PM_SKY130_FD_SC_HVL__DFXTP_1%A_1455_543#
x_PM_SKY130_FD_SC_HVL__DFXTP_1%VPWR N_VPWR_M1011_d N_VPWR_M1017_s N_VPWR_M1006_d
+ N_VPWR_M1015_d N_VPWR_M1009_s VPWR N_VPWR_c_1002_n N_VPWR_c_1005_n
+ N_VPWR_c_1008_n N_VPWR_c_1011_n N_VPWR_c_1014_n N_VPWR_c_1017_n
+ PM_SKY130_FD_SC_HVL__DFXTP_1%VPWR
x_PM_SKY130_FD_SC_HVL__DFXTP_1%A_605_563# N_A_605_563#_M1016_d
+ N_A_605_563#_M1017_d N_A_605_563#_c_1077_n N_A_605_563#_c_1076_n
+ N_A_605_563#_c_1078_n N_A_605_563#_c_1079_n N_A_605_563#_c_1080_n
+ PM_SKY130_FD_SC_HVL__DFXTP_1%A_605_563#
x_PM_SKY130_FD_SC_HVL__DFXTP_1%Q N_Q_M1023_d N_Q_M1009_d Q Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_HVL__DFXTP_1%Q
x_PM_SKY130_FD_SC_HVL__DFXTP_1%VGND N_VGND_M1022_d N_VGND_M1016_s N_VGND_M1007_d
+ N_VGND_M1008_d N_VGND_M1023_s VGND N_VGND_c_1129_n N_VGND_c_1131_n
+ N_VGND_c_1133_n N_VGND_c_1135_n N_VGND_c_1137_n N_VGND_c_1139_n
+ PM_SKY130_FD_SC_HVL__DFXTP_1%VGND
cc_1 N_VNB_M1022_b N_CLK_c_196_n 0.0259098f $X=-0.33 $Y=-0.265 $X2=0.675
+ $Y2=1.425
cc_2 N_VNB_M1022_b N_CLK_c_197_n 0.0420396f $X=-0.33 $Y=-0.265 $X2=0.675
+ $Y2=1.165
cc_3 N_VNB_c_3_p N_CLK_c_197_n 5.23624e-19 $X=0.24 $Y=0 $X2=0.675 $Y2=1.165
cc_4 N_VNB_M1022_b N_CLK_c_199_n 0.0437014f $X=-0.33 $Y=-0.265 $X2=0.705
+ $Y2=2.07
cc_5 N_VNB_M1022_b N_A_30_127#_M1004_g 0.0459046f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=2.32
cc_6 N_VNB_c_3_p N_A_30_127#_M1004_g 8.56083e-19 $X=0.24 $Y=0 $X2=0.635 $Y2=2.32
cc_7 N_VNB_M1022_b N_A_30_127#_M1013_g 0.0418568f $X=-0.33 $Y=-0.265 $X2=0.705
+ $Y2=2.07
cc_8 N_VNB_M1022_b N_A_30_127#_c_229_n 0.12885f $X=-0.33 $Y=-0.265 $X2=0.705
+ $Y2=2.035
cc_9 N_VNB_M1022_b N_A_30_127#_c_230_n 0.0261797f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_10 N_VNB_M1022_b N_A_30_127#_c_231_n 0.0220865f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1022_b N_A_30_127#_c_232_n 0.0657023f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1022_b N_A_30_127#_M1002_g 0.0478232f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_c_3_p N_A_30_127#_M1002_g 0.00224751f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_14 N_VNB_M1022_b N_A_30_127#_c_235_n 0.0311952f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_15 N_VNB_M1022_b N_A_30_127#_c_236_n 0.0517247f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_16 N_VNB_c_3_p N_A_30_127#_c_236_n 5.46509e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_17 N_VNB_M1022_b N_A_30_127#_c_238_n 0.00797076f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1022_b N_A_30_127#_c_239_n 0.0124687f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_19 N_VNB_M1022_b N_A_30_127#_c_240_n 0.00734273f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_20 N_VNB_M1022_b N_A_30_127#_c_241_n 0.00852418f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_21 N_VNB_M1022_b N_A_30_127#_c_242_n 0.0397658f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_22 N_VNB_M1022_b N_D_c_416_n 0.0037955f $X=-0.33 $Y=-0.265 $X2=0.665 $Y2=3.17
cc_23 N_VNB_M1022_b N_D_M1016_g 0.0705126f $X=-0.33 $Y=-0.265 $X2=0.675
+ $Y2=1.165
cc_24 N_VNB_c_3_p N_D_M1016_g 8.13598e-19 $X=0.24 $Y=0 $X2=0.675 $Y2=1.165
cc_25 N_VNB_M1022_b N_D_c_419_n 0.00791993f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_26 N_VNB_M1022_b N_D_c_420_n 0.102661f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_27 N_VNB_M1022_b N_A_339_559#_c_472_n 0.0164506f $X=-0.33 $Y=-0.265 $X2=0.675
+ $Y2=2.07
cc_28 N_VNB_c_3_p N_A_339_559#_c_472_n 7.21284e-19 $X=0.24 $Y=0 $X2=0.675
+ $Y2=2.07
cc_29 N_VNB_M1022_b N_A_339_559#_c_474_n 0.00840579f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_30 N_VNB_M1022_b N_A_339_559#_c_475_n 0.00320349f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_31 N_VNB_M1022_b N_A_339_559#_c_476_n 0.155212f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_32 N_VNB_c_3_p N_A_339_559#_c_476_n 0.00653204f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_33 N_VNB_M1022_b N_A_339_559#_c_478_n 0.013657f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_c_3_p N_A_339_559#_c_478_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_35 N_VNB_M1022_b N_A_339_559#_c_480_n 0.00950699f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_36 N_VNB_M1022_b N_A_339_559#_c_481_n 0.0730402f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_37 N_VNB_c_3_p N_A_339_559#_c_481_n 0.00301162f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_38 N_VNB_M1022_b N_A_339_559#_c_483_n 0.013657f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_39 N_VNB_c_3_p N_A_339_559#_c_483_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_40 N_VNB_M1022_b N_A_339_559#_c_485_n 0.00493931f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_41 N_VNB_M1022_b N_A_339_559#_c_486_n 0.00357589f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_42 N_VNB_M1022_b N_A_339_559#_M1005_g 0.0894044f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_M1022_b N_A_339_559#_M1010_g 0.0829991f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_44 N_VNB_c_3_p N_A_339_559#_M1010_g 9.21478e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_45 N_VNB_M1022_b N_A_1024_371#_M1007_g 0.109849f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=2.32
cc_46 N_VNB_M1022_b N_A_1024_371#_c_690_n 0.00196674f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_47 N_VNB_M1022_b N_A_1024_371#_c_691_n 0.00744164f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_M1022_b N_A_1024_371#_c_692_n 0.00775097f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_49 N_VNB_M1022_b N_A_1024_371#_c_693_n 6.85236e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_M1022_b N_A_780_574#_c_758_n 0.10135f $X=-0.33 $Y=-0.265 $X2=0.675
+ $Y2=2.665
cc_51 N_VNB_c_3_p N_A_780_574#_c_758_n 5.61877e-19 $X=0.24 $Y=0 $X2=0.675
+ $Y2=2.665
cc_52 N_VNB_M1022_b N_A_780_574#_c_760_n 0.00505629f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=2.07
cc_53 N_VNB_M1022_b N_A_780_574#_c_761_n 0.0180813f $X=-0.33 $Y=-0.265 $X2=0.705
+ $Y2=2.405
cc_54 N_VNB_M1022_b N_A_780_574#_c_762_n 0.00580575f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_55 N_VNB_M1022_b N_A_780_574#_c_763_n 0.00181934f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_56 N_VNB_M1022_b N_A_1729_87#_M1008_g 0.062197f $X=-0.33 $Y=-0.265 $X2=0.675
+ $Y2=1.165
cc_57 N_VNB_c_3_p N_A_1729_87#_M1008_g 6.11322e-19 $X=0.24 $Y=0 $X2=0.675
+ $Y2=1.165
cc_58 N_VNB_M1022_b N_A_1729_87#_M1023_g 0.0518045f $X=-0.33 $Y=-0.265 $X2=0.705
+ $Y2=2.07
cc_59 N_VNB_c_3_p N_A_1729_87#_M1023_g 0.00117942f $X=0.24 $Y=0 $X2=0.705
+ $Y2=2.07
cc_60 N_VNB_M1022_b N_A_1729_87#_c_834_n 0.014362f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_61 N_VNB_M1022_b N_A_1729_87#_c_835_n 0.018024f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_62 N_VNB_c_3_p N_A_1729_87#_c_835_n 7.88607e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_63 N_VNB_M1022_b N_A_1729_87#_c_837_n 0.00200133f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_64 N_VNB_M1022_b N_A_1729_87#_c_838_n 0.0234112f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_65 N_VNB_M1022_b N_A_1729_87#_c_839_n 0.0693091f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_66 N_VNB_M1022_b N_A_1729_87#_c_840_n 0.0441286f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_67 N_VNB_M1022_b N_A_1455_543#_M1019_g 0.0543077f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=1.165
cc_68 N_VNB_c_3_p N_A_1455_543#_M1019_g 0.00213963f $X=0.24 $Y=0 $X2=0.675
+ $Y2=1.165
cc_69 N_VNB_M1022_b N_A_1455_543#_c_911_n 0.0424398f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=2.665
cc_70 N_VNB_M1022_b N_A_1455_543#_c_912_n 2.34417e-19 $X=-0.33 $Y=-0.265
+ $X2=0.705 $Y2=2.035
cc_71 N_VNB_M1022_b N_A_1455_543#_c_913_n 0.00857823f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_72 N_VNB_M1022_b N_A_1455_543#_c_914_n 0.0130523f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_73 N_VNB_c_3_p N_A_1455_543#_c_914_n 0.00103607f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_74 N_VNB_M1022_b N_A_605_563#_c_1076_n 0.00605009f $X=-0.33 $Y=-0.265
+ $X2=0.675 $Y2=2.665
cc_75 N_VNB_M1022_b Q 0.0581789f $X=-0.33 $Y=-0.265 $X2=0.685 $Y2=0.845
cc_76 N_VNB_M1022_b N_VGND_c_1129_n 0.053203f $X=-0.33 $Y=-0.265 $X2=0.705
+ $Y2=2.035
cc_77 N_VNB_c_3_p N_VGND_c_1129_n 0.00269049f $X=0.24 $Y=0 $X2=0.705 $Y2=2.035
cc_78 N_VNB_M1022_b N_VGND_c_1131_n 0.0431017f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_79 N_VNB_c_3_p N_VGND_c_1131_n 0.00159858f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_80 N_VNB_M1022_b N_VGND_c_1133_n 0.050587f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_81 N_VNB_c_3_p N_VGND_c_1133_n 0.00269373f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_82 N_VNB_M1022_b N_VGND_c_1135_n 0.0524215f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_83 N_VNB_c_3_p N_VGND_c_1135_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_84 N_VNB_M1022_b N_VGND_c_1137_n 0.0489282f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_85 N_VNB_c_3_p N_VGND_c_1137_n 0.00166879f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_86 N_VNB_M1022_b N_VGND_c_1139_n 0.167031f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_87 N_VNB_c_3_p N_VGND_c_1139_n 1.28268f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_88 N_VPB_M1011_b N_CLK_M1011_g 0.0401459f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=3.17
cc_89 VPB N_CLK_M1011_g 5.93461e-19 $X=0 $Y=3.955 $X2=0.665 $Y2=3.17
cc_90 N_VPB_c_90_p N_CLK_M1011_g 0.00487048f $X=11.76 $Y=4.07 $X2=0.665 $Y2=3.17
cc_91 N_VPB_M1011_b N_CLK_c_203_n 0.02554f $X=-0.33 $Y=1.885 $X2=0.675 $Y2=2.665
cc_92 N_VPB_M1011_b N_CLK_c_199_n 0.0499336f $X=-0.33 $Y=1.885 $X2=0.705
+ $Y2=2.07
cc_93 N_VPB_M1011_b N_A_30_127#_c_243_n 0.0696802f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=0.845
cc_94 N_VPB_M1011_b N_A_30_127#_M1001_g 0.0408157f $X=-0.33 $Y=1.885 $X2=0.675
+ $Y2=1.165
cc_95 VPB N_A_30_127#_M1001_g 9.70262e-19 $X=0 $Y=3.955 $X2=0.675 $Y2=1.165
cc_96 N_VPB_c_90_p N_A_30_127#_M1001_g 0.0061414f $X=11.76 $Y=4.07 $X2=0.675
+ $Y2=1.165
cc_97 N_VPB_M1011_b N_A_30_127#_c_229_n 0.111005f $X=-0.33 $Y=1.885 $X2=0.705
+ $Y2=2.035
cc_98 N_VPB_M1011_b N_A_30_127#_M1000_g 0.0375644f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_99 N_VPB_M1011_b N_A_30_127#_c_230_n 0.132015f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_100 VPB N_A_30_127#_c_230_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_101 N_VPB_c_90_p N_A_30_127#_c_230_n 0.0196751f $X=11.76 $Y=4.07 $X2=0 $Y2=0
cc_102 N_VPB_M1011_b N_A_30_127#_c_231_n 0.0160198f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_103 N_VPB_M1011_b N_A_30_127#_c_232_n 0.0177588f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_104 N_VPB_M1011_b N_A_30_127#_c_238_n 0.075195f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_105 VPB N_A_30_127#_c_238_n 5.72987e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_106 N_VPB_c_90_p N_A_30_127#_c_238_n 0.00676138f $X=11.76 $Y=4.07 $X2=0 $Y2=0
cc_107 N_VPB_M1011_b N_A_30_127#_c_257_n 0.00843062f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_108 N_VPB_M1011_b N_A_30_127#_c_240_n 0.00779299f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_109 N_VPB_M1011_b N_A_30_127#_c_259_n 0.0202436f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_110 N_VPB_M1011_b N_A_30_127#_c_242_n 0.00735241f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_111 N_VPB_M1011_b N_A_30_127#_c_261_n 0.00703994f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_112 N_VPB_M1011_b N_D_c_416_n 0.0287002f $X=-0.33 $Y=1.885 $X2=0.665 $Y2=3.17
cc_113 N_VPB_M1011_b N_D_M1017_g 0.0407787f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=1.165
cc_114 N_VPB_c_90_p N_D_M1017_g 0.00393173f $X=11.76 $Y=4.07 $X2=0.685 $Y2=1.165
cc_115 N_VPB_M1011_b N_D_c_424_n 0.0889384f $X=-0.33 $Y=1.885 $X2=0.635 $Y2=2.32
cc_116 N_VPB_M1011_b N_A_339_559#_c_490_n 0.108488f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=0.845
cc_117 N_VPB_M1011_b N_A_339_559#_c_491_n 0.0114392f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.95
cc_118 VPB N_A_339_559#_c_491_n 8.09367e-19 $X=0 $Y=3.955 $X2=0.635 $Y2=1.95
cc_119 N_VPB_c_90_p N_A_339_559#_c_491_n 0.00884658f $X=11.76 $Y=4.07 $X2=0.635
+ $Y2=1.95
cc_120 N_VPB_M1011_b N_A_339_559#_c_494_n 0.00528627f $X=-0.33 $Y=1.885
+ $X2=0.705 $Y2=2.07
cc_121 N_VPB_M1011_b N_A_339_559#_c_495_n 0.00348063f $X=-0.33 $Y=1.885
+ $X2=0.705 $Y2=2.035
cc_122 N_VPB_M1011_b N_A_339_559#_c_496_n 0.0108737f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_123 VPB N_A_339_559#_c_496_n 0.0014439f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_124 N_VPB_c_90_p N_A_339_559#_c_496_n 0.0140502f $X=11.76 $Y=4.07 $X2=0 $Y2=0
cc_125 N_VPB_M1011_b N_A_339_559#_c_499_n 0.00223349f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_126 VPB N_A_339_559#_c_499_n 3.46666e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_127 N_VPB_c_90_p N_A_339_559#_c_499_n 0.00355965f $X=11.76 $Y=4.07 $X2=0
+ $Y2=0
cc_128 N_VPB_M1011_b N_A_339_559#_c_502_n 0.100587f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_129 N_VPB_c_90_p N_A_339_559#_c_502_n 0.00607399f $X=11.76 $Y=4.07 $X2=0
+ $Y2=0
cc_130 N_VPB_M1011_b N_A_339_559#_c_504_n 0.0230895f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_131 N_VPB_M1011_b N_A_339_559#_c_485_n 0.00717989f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_132 N_VPB_M1011_b N_A_339_559#_c_506_n 0.00288281f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_133 N_VPB_M1011_b N_A_339_559#_c_507_n 0.01018f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_134 N_VPB_M1011_b N_A_339_559#_c_508_n 0.00277409f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_135 VPB N_A_339_559#_c_508_n 3.46666e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_136 N_VPB_c_90_p N_A_339_559#_c_508_n 0.00355965f $X=11.76 $Y=4.07 $X2=0
+ $Y2=0
cc_137 N_VPB_M1011_b N_A_1024_371#_M1006_g 0.0366896f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=1.165
cc_138 N_VPB_M1011_b N_A_1024_371#_c_690_n 0.00523406f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_139 N_VPB_M1011_b N_A_1024_371#_c_696_n 0.00102083f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_140 N_VPB_M1011_b N_A_1024_371#_c_692_n 0.0754549f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_141 N_VPB_M1011_b N_A_1024_371#_c_693_n 0.00171275f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_142 N_VPB_M1011_b N_A_780_574#_M1003_g 0.0956674f $X=-0.33 $Y=1.885 $X2=0.675
+ $Y2=1.165
cc_143 VPB N_A_780_574#_M1003_g 0.00970178f $X=0 $Y=3.955 $X2=0.675 $Y2=1.165
cc_144 N_VPB_c_90_p N_A_780_574#_M1003_g 0.0193818f $X=11.76 $Y=4.07 $X2=0.675
+ $Y2=1.165
cc_145 N_VPB_M1011_b N_A_780_574#_c_758_n 0.009104f $X=-0.33 $Y=1.885 $X2=0.675
+ $Y2=2.665
cc_146 N_VPB_M1011_b N_A_780_574#_c_768_n 0.00364229f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_147 N_VPB_M1011_b N_A_780_574#_c_762_n 0.00156584f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_148 N_VPB_M1011_b N_A_1729_87#_M1015_g 0.088314f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=2.32
cc_149 N_VPB_M1011_b N_A_1729_87#_M1009_g 0.0436128f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_150 VPB N_A_1729_87#_M1009_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_151 N_VPB_c_90_p N_A_1729_87#_M1009_g 0.0167053f $X=11.76 $Y=4.07 $X2=0 $Y2=0
cc_152 N_VPB_M1011_b N_A_1729_87#_c_845_n 0.0170873f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_153 VPB N_A_1729_87#_c_845_n 0.00101808f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_154 N_VPB_c_90_p N_A_1729_87#_c_845_n 0.0158392f $X=11.76 $Y=4.07 $X2=0 $Y2=0
cc_155 N_VPB_M1011_b N_A_1729_87#_c_838_n 0.0156074f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_156 N_VPB_M1011_b N_A_1729_87#_c_839_n 0.0210767f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_157 N_VPB_M1011_b N_A_1729_87#_c_840_n 0.0366139f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_158 N_VPB_M1011_b N_A_1455_543#_c_911_n 0.0598478f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=2.665
cc_159 N_VPB_M1011_b N_A_1455_543#_M1018_g 0.0554546f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=2.32
cc_160 VPB N_A_1455_543#_M1018_g 0.00970178f $X=0 $Y=3.955 $X2=0.635 $Y2=2.32
cc_161 N_VPB_c_90_p N_A_1455_543#_M1018_g 0.0191116f $X=11.76 $Y=4.07 $X2=0.635
+ $Y2=2.32
cc_162 N_VPB_M1011_b N_A_1455_543#_c_920_n 0.00190281f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_163 N_VPB_M1011_b N_A_1455_543#_c_921_n 0.0139166f $X=-0.33 $Y=1.885
+ $X2=0.705 $Y2=2.07
cc_164 VPB N_A_1455_543#_c_921_n 7.36921e-19 $X=0 $Y=3.955 $X2=0.705 $Y2=2.07
cc_165 N_VPB_c_90_p N_A_1455_543#_c_921_n 0.0120479f $X=11.76 $Y=4.07 $X2=0.705
+ $Y2=2.07
cc_166 N_VPB_M1011_b N_A_1455_543#_c_924_n 4.0946e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_167 N_VPB_M1011_b N_A_1455_543#_c_913_n 0.0125647f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_168 N_VPB_M1011_b N_A_1455_543#_c_926_n 0.022585f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_169 N_VPB_M1011_b N_VPWR_c_1002_n 0.0150148f $X=-0.33 $Y=1.885 $X2=0.705
+ $Y2=2.035
cc_170 VPB N_VPWR_c_1002_n 0.00269049f $X=0 $Y=3.955 $X2=0.705 $Y2=2.035
cc_171 N_VPB_c_90_p N_VPWR_c_1002_n 0.0409968f $X=11.76 $Y=4.07 $X2=0.705
+ $Y2=2.035
cc_172 N_VPB_M1011_b N_VPWR_c_1005_n 0.020083f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1005_n 7.03841e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_174 N_VPB_c_90_p N_VPWR_c_1005_n 0.0107249f $X=11.76 $Y=4.07 $X2=0 $Y2=0
cc_175 N_VPB_M1011_b N_VPWR_c_1008_n 0.0161267f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1008_n 0.00289756f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_177 N_VPB_c_90_p N_VPWR_c_1008_n 0.0451371f $X=11.76 $Y=4.07 $X2=0 $Y2=0
cc_178 N_VPB_M1011_b N_VPWR_c_1011_n 0.028542f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1011_n 0.00286038f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_180 N_VPB_c_90_p N_VPWR_c_1011_n 0.0459589f $X=11.76 $Y=4.07 $X2=0 $Y2=0
cc_181 N_VPB_M1011_b N_VPWR_c_1014_n 0.0197226f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1014_n 0.0021617f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_183 N_VPB_c_90_p N_VPWR_c_1014_n 0.0276576f $X=11.76 $Y=4.07 $X2=0 $Y2=0
cc_184 N_VPB_M1011_b N_VPWR_c_1017_n 0.14872f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1017_n 1.28053f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_186 N_VPB_c_90_p N_VPWR_c_1017_n 0.0676499f $X=11.76 $Y=4.07 $X2=0 $Y2=0
cc_187 N_VPB_M1011_b N_A_605_563#_c_1077_n 0.00603119f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=1.165
cc_188 N_VPB_M1011_b N_A_605_563#_c_1078_n 0.0131265f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_189 N_VPB_M1011_b N_A_605_563#_c_1079_n 0.00337234f $X=-0.33 $Y=1.885
+ $X2=0.675 $Y2=2.07
cc_190 N_VPB_M1011_b N_A_605_563#_c_1080_n 0.00774156f $X=-0.33 $Y=1.885
+ $X2=0.705 $Y2=2.07
cc_191 N_VPB_M1011_b Q 0.0151104f $X=-0.33 $Y=1.885 $X2=0.685 $Y2=0.845
cc_192 N_VPB_M1011_b Q 0.00872165f $X=-0.33 $Y=1.885 $X2=0.675 $Y2=2.665
cc_193 N_VPB_M1011_b Q 0.04802f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_194 VPB Q 0.00101808f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_195 N_VPB_c_90_p Q 0.0158392f $X=11.76 $Y=4.07 $X2=0 $Y2=0
cc_196 N_CLK_c_203_n N_A_30_127#_c_243_n 0.0360253f $X=0.675 $Y=2.665 $X2=0
+ $Y2=0
cc_197 N_CLK_M1011_g N_A_30_127#_M1001_g 0.0181863f $X=0.665 $Y=3.17 $X2=0 $Y2=0
cc_198 N_CLK_c_197_n N_A_30_127#_M1004_g 0.0145436f $X=0.675 $Y=1.165 $X2=0
+ $Y2=0
cc_199 N_CLK_c_196_n N_A_30_127#_c_235_n 0.0360253f $X=0.675 $Y=1.425 $X2=0
+ $Y2=0
cc_200 N_CLK_c_196_n N_A_30_127#_c_236_n 0.0188108f $X=0.675 $Y=1.425 $X2=0
+ $Y2=0
cc_201 N_CLK_c_197_n N_A_30_127#_c_236_n 0.00609542f $X=0.675 $Y=1.165 $X2=0
+ $Y2=0
cc_202 CLK N_A_30_127#_c_238_n 0.0496484f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_203 N_CLK_c_199_n N_A_30_127#_c_238_n 0.0394454f $X=0.705 $Y=2.07 $X2=0 $Y2=0
cc_204 CLK N_A_30_127#_c_239_n 0.0238298f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_205 N_CLK_c_199_n N_A_30_127#_c_239_n 0.041485f $X=0.705 $Y=2.07 $X2=0 $Y2=0
cc_206 CLK N_A_30_127#_c_272_n 0.0162565f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_207 N_CLK_c_199_n N_A_30_127#_c_272_n 0.00250189f $X=0.705 $Y=2.07 $X2=0
+ $Y2=0
cc_208 CLK N_A_30_127#_c_242_n 0.00337473f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_209 N_CLK_c_199_n N_A_30_127#_c_242_n 0.0360253f $X=0.705 $Y=2.07 $X2=0 $Y2=0
cc_210 N_CLK_M1011_g N_VPWR_c_1002_n 0.0570878f $X=0.665 $Y=3.17 $X2=0 $Y2=0
cc_211 N_CLK_c_203_n N_VPWR_c_1002_n 0.0010557f $X=0.675 $Y=2.665 $X2=0 $Y2=0
cc_212 CLK N_VPWR_c_1002_n 0.0264771f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_213 N_CLK_M1011_g N_VPWR_c_1017_n 0.00868732f $X=0.665 $Y=3.17 $X2=0 $Y2=0
cc_214 N_CLK_c_197_n N_VGND_c_1129_n 0.0449384f $X=0.675 $Y=1.165 $X2=0 $Y2=0
cc_215 N_CLK_c_196_n N_VGND_c_1139_n 5.07648e-19 $X=0.675 $Y=1.425 $X2=0 $Y2=0
cc_216 N_CLK_c_197_n N_VGND_c_1139_n 0.00879041f $X=0.675 $Y=1.165 $X2=0 $Y2=0
cc_217 N_A_30_127#_c_257_n N_D_c_416_n 0.0273086f $X=2.65 $Y=2.077 $X2=0 $Y2=0
cc_218 N_A_30_127#_c_242_n N_D_c_416_n 0.0105603f $X=1.33 $Y=1.72 $X2=0 $Y2=0
cc_219 N_A_30_127#_c_261_n N_D_c_416_n 0.00891161f $X=2.735 $Y=1.845 $X2=0 $Y2=0
cc_220 N_A_30_127#_M1013_g N_D_M1016_g 0.0145102f $X=3.85 $Y=0.775 $X2=0 $Y2=0
cc_221 N_A_30_127#_c_229_n N_D_M1016_g 0.0527675f $X=4.66 $Y=2.585 $X2=0 $Y2=0
cc_222 N_A_30_127#_c_281_p N_D_M1016_g 0.00348868f $X=3.595 $Y=1.37 $X2=0 $Y2=0
cc_223 N_A_30_127#_c_243_n N_D_c_424_n 0.0253057f $X=1.445 $Y=2.665 $X2=0 $Y2=0
cc_224 N_A_30_127#_c_257_n N_D_c_424_n 0.0112011f $X=2.65 $Y=2.077 $X2=0 $Y2=0
cc_225 N_A_30_127#_c_240_n N_D_c_424_n 0.00379844f $X=3.43 $Y=1.845 $X2=0 $Y2=0
cc_226 N_A_30_127#_c_261_n N_D_c_424_n 0.00573984f $X=2.735 $Y=1.845 $X2=0 $Y2=0
cc_227 N_A_30_127#_c_286_p N_D_c_419_n 0.0136575f $X=1.29 $Y=1.725 $X2=6 $Y2=0
cc_228 N_A_30_127#_c_272_n N_D_c_419_n 0.00175897f $X=1.29 $Y=1.93 $X2=6 $Y2=0
cc_229 N_A_30_127#_c_257_n N_D_c_419_n 0.062977f $X=2.65 $Y=2.077 $X2=6 $Y2=0
cc_230 N_A_30_127#_c_242_n N_D_c_419_n 0.0143312f $X=1.33 $Y=1.72 $X2=6 $Y2=0
cc_231 N_A_30_127#_c_235_n N_D_c_420_n 0.0105603f $X=1.43 $Y=1.47 $X2=6
+ $Y2=0.058
cc_232 N_A_30_127#_c_240_n N_D_c_420_n 0.0181489f $X=3.43 $Y=1.845 $X2=6
+ $Y2=0.058
cc_233 N_A_30_127#_c_261_n N_D_c_420_n 0.0103113f $X=2.735 $Y=1.845 $X2=6
+ $Y2=0.058
cc_234 N_A_30_127#_c_230_n N_A_339_559#_c_490_n 0.0107097f $X=7.025 $Y=2.605
+ $X2=0 $Y2=0
cc_235 N_A_30_127#_c_231_n N_A_339_559#_c_490_n 0.0381983f $X=7.905 $Y=1.845
+ $X2=0 $Y2=0
cc_236 N_A_30_127#_c_232_n N_A_339_559#_c_490_n 9.68265e-19 $X=8.185 $Y=1.115
+ $X2=0 $Y2=0
cc_237 N_A_30_127#_c_243_n N_A_339_559#_c_491_n 0.00298107f $X=1.445 $Y=2.665
+ $X2=0 $Y2=0
cc_238 N_A_30_127#_M1001_g N_A_339_559#_c_491_n 0.0213841f $X=1.445 $Y=3.17
+ $X2=0 $Y2=0
cc_239 N_A_30_127#_M1004_g N_A_339_559#_c_472_n 0.0165884f $X=1.465 $Y=0.845
+ $X2=11.76 $Y2=0
cc_240 N_A_30_127#_c_235_n N_A_339_559#_c_472_n 0.00128754f $X=1.43 $Y=1.47
+ $X2=11.76 $Y2=0
cc_241 N_A_30_127#_c_257_n N_A_339_559#_c_494_n 0.0383377f $X=2.65 $Y=2.077
+ $X2=0 $Y2=0
cc_242 N_A_30_127#_c_261_n N_A_339_559#_c_494_n 0.0112221f $X=2.735 $Y=1.845
+ $X2=0 $Y2=0
cc_243 N_A_30_127#_c_243_n N_A_339_559#_c_495_n 0.012452f $X=1.445 $Y=2.665
+ $X2=0 $Y2=0
cc_244 N_A_30_127#_c_257_n N_A_339_559#_c_495_n 0.0238516f $X=2.65 $Y=2.077
+ $X2=0 $Y2=0
cc_245 N_A_30_127#_c_229_n N_A_339_559#_c_474_n 6.06251e-19 $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_246 N_A_30_127#_c_257_n N_A_339_559#_c_474_n 0.00481908f $X=2.65 $Y=2.077
+ $X2=0 $Y2=0
cc_247 N_A_30_127#_c_240_n N_A_339_559#_c_474_n 0.0110634f $X=3.43 $Y=1.845
+ $X2=0 $Y2=0
cc_248 N_A_30_127#_c_281_p N_A_339_559#_c_474_n 0.00808838f $X=3.595 $Y=1.37
+ $X2=0 $Y2=0
cc_249 N_A_30_127#_c_261_n N_A_339_559#_c_474_n 0.00640737f $X=2.735 $Y=1.845
+ $X2=0 $Y2=0
cc_250 N_A_30_127#_c_235_n N_A_339_559#_c_475_n 0.0130384f $X=1.43 $Y=1.47 $X2=6
+ $Y2=0
cc_251 N_A_30_127#_M1013_g N_A_339_559#_c_528_n 0.00185727f $X=3.85 $Y=0.775
+ $X2=0 $Y2=0
cc_252 N_A_30_127#_c_229_n N_A_339_559#_c_528_n 5.71179e-19 $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_253 N_A_30_127#_M1013_g N_A_339_559#_c_476_n 0.0134651f $X=3.85 $Y=0.775
+ $X2=0 $Y2=0
cc_254 N_A_30_127#_c_229_n N_A_339_559#_c_476_n 0.00256128f $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_255 N_A_30_127#_c_229_n N_A_339_559#_c_532_n 4.87016e-19 $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_256 N_A_30_127#_M1000_g N_A_339_559#_c_532_n 7.75035e-19 $X=4.66 $Y=2.925
+ $X2=0 $Y2=0
cc_257 N_A_30_127#_c_229_n N_A_339_559#_c_502_n 0.0418557f $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_258 N_A_30_127#_M1000_g N_A_339_559#_c_502_n 0.0109668f $X=4.66 $Y=2.925
+ $X2=0 $Y2=0
cc_259 N_A_30_127#_c_240_n N_A_339_559#_c_502_n 8.99937e-19 $X=3.43 $Y=1.845
+ $X2=0 $Y2=0
cc_260 N_A_30_127#_c_229_n N_A_339_559#_c_504_n 0.00140203f $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_261 N_A_30_127#_M1000_g N_A_339_559#_c_504_n 0.0330598f $X=4.66 $Y=2.925
+ $X2=0 $Y2=0
cc_262 N_A_30_127#_c_230_n N_A_339_559#_c_504_n 0.032546f $X=7.025 $Y=2.605
+ $X2=0 $Y2=0
cc_263 N_A_30_127#_c_259_n N_A_339_559#_c_504_n 0.0414391f $X=6.705 $Y=2.47
+ $X2=0 $Y2=0
cc_264 N_A_30_127#_c_323_p N_A_339_559#_c_504_n 0.0089596f $X=4.89 $Y=2.47 $X2=0
+ $Y2=0
cc_265 N_A_30_127#_M1013_g N_A_339_559#_c_542_n 0.0011373f $X=3.85 $Y=0.775
+ $X2=0 $Y2=0
cc_266 N_A_30_127#_M1002_g N_A_339_559#_c_543_n 0.00122402f $X=8.185 $Y=0.775
+ $X2=0 $Y2=0
cc_267 N_A_30_127#_c_230_n N_A_339_559#_c_485_n 0.0138823f $X=7.025 $Y=2.605
+ $X2=0 $Y2=0
cc_268 N_A_30_127#_c_231_n N_A_339_559#_c_485_n 0.025093f $X=7.905 $Y=1.845
+ $X2=0 $Y2=0
cc_269 N_A_30_127#_c_232_n N_A_339_559#_c_485_n 0.00783183f $X=8.185 $Y=1.115
+ $X2=0 $Y2=0
cc_270 N_A_30_127#_c_230_n N_A_339_559#_c_506_n 0.0116461f $X=7.025 $Y=2.605
+ $X2=0 $Y2=0
cc_271 N_A_30_127#_c_231_n N_A_339_559#_c_507_n 0.0120526f $X=7.905 $Y=1.845
+ $X2=0 $Y2=0
cc_272 N_A_30_127#_c_230_n N_A_339_559#_c_486_n 0.0015337f $X=7.025 $Y=2.605
+ $X2=0 $Y2=0
cc_273 N_A_30_127#_c_232_n N_A_339_559#_c_486_n 0.00231809f $X=8.185 $Y=1.115
+ $X2=0 $Y2=0
cc_274 N_A_30_127#_c_230_n N_A_339_559#_c_551_n 0.00929005f $X=7.025 $Y=2.605
+ $X2=0 $Y2=0
cc_275 N_A_30_127#_M1013_g N_A_339_559#_M1005_g 0.0107188f $X=3.85 $Y=0.775
+ $X2=0 $Y2=0
cc_276 N_A_30_127#_c_229_n N_A_339_559#_M1005_g 0.041997f $X=4.66 $Y=2.585 $X2=0
+ $Y2=0
cc_277 N_A_30_127#_c_336_p N_A_339_559#_M1005_g 3.20975e-19 $X=4.725 $Y=2.05
+ $X2=0 $Y2=0
cc_278 N_A_30_127#_c_230_n N_A_339_559#_M1010_g 0.0364277f $X=7.025 $Y=2.605
+ $X2=0 $Y2=0
cc_279 N_A_30_127#_c_232_n N_A_339_559#_M1010_g 0.0187234f $X=8.185 $Y=1.115
+ $X2=0 $Y2=0
cc_280 N_A_30_127#_M1002_g N_A_339_559#_M1010_g 0.0146369f $X=8.185 $Y=0.775
+ $X2=0 $Y2=0
cc_281 N_A_30_127#_M1000_g N_A_1024_371#_M1006_g 0.0519903f $X=4.66 $Y=2.925
+ $X2=0 $Y2=0
cc_282 N_A_30_127#_c_230_n N_A_1024_371#_c_690_n 0.00821524f $X=7.025 $Y=2.605
+ $X2=0 $Y2=0
cc_283 N_A_30_127#_c_259_n N_A_1024_371#_c_690_n 0.039801f $X=6.705 $Y=2.47
+ $X2=0 $Y2=0
cc_284 N_A_30_127#_c_343_p N_A_1024_371#_c_690_n 0.0178975f $X=6.87 $Y=2.39
+ $X2=0 $Y2=0
cc_285 N_A_30_127#_c_230_n N_A_1024_371#_c_703_n 0.0316602f $X=7.025 $Y=2.605
+ $X2=11.76 $Y2=0
cc_286 N_A_30_127#_c_259_n N_A_1024_371#_c_703_n 0.0135778f $X=6.705 $Y=2.47
+ $X2=11.76 $Y2=0
cc_287 N_A_30_127#_c_343_p N_A_1024_371#_c_703_n 0.0140606f $X=6.87 $Y=2.39
+ $X2=11.76 $Y2=0
cc_288 N_A_30_127#_c_230_n N_A_1024_371#_c_691_n 0.00973775f $X=7.025 $Y=2.605
+ $X2=6 $Y2=0.057
cc_289 N_A_30_127#_c_230_n N_A_1024_371#_c_696_n 0.0340193f $X=7.025 $Y=2.605
+ $X2=0 $Y2=0
cc_290 N_A_30_127#_c_343_p N_A_1024_371#_c_696_n 0.0220177f $X=6.87 $Y=2.39
+ $X2=0 $Y2=0
cc_291 N_A_30_127#_c_229_n N_A_1024_371#_c_709_n 8.47675e-19 $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_292 N_A_30_127#_c_336_p N_A_1024_371#_c_709_n 0.0092138f $X=4.725 $Y=2.05
+ $X2=0 $Y2=0
cc_293 N_A_30_127#_c_259_n N_A_1024_371#_c_709_n 0.0224849f $X=6.705 $Y=2.47
+ $X2=0 $Y2=0
cc_294 N_A_30_127#_c_229_n N_A_1024_371#_c_692_n 0.0519903f $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_295 N_A_30_127#_c_336_p N_A_1024_371#_c_692_n 0.00276533f $X=4.725 $Y=2.05
+ $X2=0 $Y2=0
cc_296 N_A_30_127#_c_259_n N_A_1024_371#_c_692_n 0.0482355f $X=6.705 $Y=2.47
+ $X2=0 $Y2=0
cc_297 N_A_30_127#_c_230_n N_A_1024_371#_c_693_n 0.0226999f $X=7.025 $Y=2.605
+ $X2=0 $Y2=0
cc_298 N_A_30_127#_c_230_n N_A_780_574#_M1003_g 0.0889587f $X=7.025 $Y=2.605
+ $X2=0 $Y2=0
cc_299 N_A_30_127#_c_259_n N_A_780_574#_M1003_g 0.0340727f $X=6.705 $Y=2.47
+ $X2=0 $Y2=0
cc_300 N_A_30_127#_c_343_p N_A_780_574#_M1003_g 0.00130455f $X=6.87 $Y=2.39
+ $X2=0 $Y2=0
cc_301 N_A_30_127#_c_230_n N_A_780_574#_c_758_n 0.0165628f $X=7.025 $Y=2.605
+ $X2=0.24 $Y2=0
cc_302 N_A_30_127#_c_259_n N_A_780_574#_c_758_n 9.8514e-19 $X=6.705 $Y=2.47
+ $X2=0.24 $Y2=0
cc_303 N_A_30_127#_M1013_g N_A_780_574#_c_760_n 0.00531282f $X=3.85 $Y=0.775
+ $X2=11.76 $Y2=0
cc_304 N_A_30_127#_c_229_n N_A_780_574#_c_760_n 0.0163751f $X=4.66 $Y=2.585
+ $X2=11.76 $Y2=0
cc_305 N_A_30_127#_c_229_n N_A_780_574#_c_761_n 0.00376597f $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_306 N_A_30_127#_c_336_p N_A_780_574#_c_761_n 0.0236931f $X=4.725 $Y=2.05
+ $X2=0 $Y2=0
cc_307 N_A_30_127#_c_229_n N_A_780_574#_c_768_n 0.00500529f $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_308 N_A_30_127#_c_229_n N_A_780_574#_c_762_n 0.041961f $X=4.66 $Y=2.585 $X2=0
+ $Y2=0
cc_309 N_A_30_127#_M1000_g N_A_780_574#_c_762_n 0.00398626f $X=4.66 $Y=2.925
+ $X2=0 $Y2=0
cc_310 N_A_30_127#_c_336_p N_A_780_574#_c_762_n 0.034029f $X=4.725 $Y=2.05 $X2=0
+ $Y2=0
cc_311 N_A_30_127#_c_323_p N_A_780_574#_c_762_n 0.0123662f $X=4.89 $Y=2.47 $X2=0
+ $Y2=0
cc_312 N_A_30_127#_c_229_n N_A_780_574#_c_763_n 0.0154451f $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_313 N_A_30_127#_M1002_g N_A_1729_87#_M1008_g 0.0414208f $X=8.185 $Y=0.775
+ $X2=0 $Y2=0
cc_314 N_A_30_127#_c_232_n N_A_1729_87#_c_839_n 0.0600868f $X=8.185 $Y=1.115
+ $X2=0 $Y2=0
cc_315 N_A_30_127#_c_230_n N_A_1455_543#_c_921_n 0.00900964f $X=7.025 $Y=2.605
+ $X2=11.76 $Y2=0
cc_316 N_A_30_127#_M1002_g N_A_1455_543#_c_912_n 0.0330882f $X=8.185 $Y=0.775
+ $X2=0 $Y2=0
cc_317 N_A_30_127#_c_232_n N_A_1455_543#_c_924_n 5.14506e-19 $X=8.185 $Y=1.115
+ $X2=6 $Y2=0
cc_318 N_A_30_127#_c_232_n N_A_1455_543#_c_913_n 0.0358691f $X=8.185 $Y=1.115
+ $X2=6 $Y2=0.058
cc_319 N_A_30_127#_M1002_g N_A_1455_543#_c_913_n 0.00423294f $X=8.185 $Y=0.775
+ $X2=6 $Y2=0.058
cc_320 N_A_30_127#_c_231_n N_A_1455_543#_c_914_n 0.00180601f $X=7.905 $Y=1.845
+ $X2=0 $Y2=0
cc_321 N_A_30_127#_c_232_n N_A_1455_543#_c_914_n 0.00152035f $X=8.185 $Y=1.115
+ $X2=0 $Y2=0
cc_322 N_A_30_127#_M1002_g N_A_1455_543#_c_914_n 0.0155375f $X=8.185 $Y=0.775
+ $X2=0 $Y2=0
cc_323 N_A_30_127#_c_243_n N_VPWR_c_1002_n 0.00213573f $X=1.445 $Y=2.665 $X2=0
+ $Y2=0
cc_324 N_A_30_127#_M1001_g N_VPWR_c_1002_n 0.0545229f $X=1.445 $Y=3.17 $X2=0
+ $Y2=0
cc_325 N_A_30_127#_c_238_n N_VPWR_c_1002_n 0.0351665f $X=0.275 $Y=2.94 $X2=0
+ $Y2=0
cc_326 N_A_30_127#_c_272_n N_VPWR_c_1002_n 0.00841271f $X=1.29 $Y=1.93 $X2=0
+ $Y2=0
cc_327 N_A_30_127#_c_257_n N_VPWR_c_1002_n 0.00228811f $X=2.65 $Y=2.077 $X2=0
+ $Y2=0
cc_328 N_A_30_127#_M1001_g N_VPWR_c_1005_n 0.00309972f $X=1.445 $Y=3.17 $X2=0
+ $Y2=0
cc_329 N_A_30_127#_M1011_s N_VPWR_c_1017_n 0.00221032f $X=0.15 $Y=2.795 $X2=0
+ $Y2=0
cc_330 N_A_30_127#_M1001_g N_VPWR_c_1017_n 0.0121989f $X=1.445 $Y=3.17 $X2=0
+ $Y2=0
cc_331 N_A_30_127#_c_230_n N_VPWR_c_1017_n 0.0227204f $X=7.025 $Y=2.605 $X2=0
+ $Y2=0
cc_332 N_A_30_127#_c_238_n N_VPWR_c_1017_n 0.025732f $X=0.275 $Y=2.94 $X2=0
+ $Y2=0
cc_333 N_A_30_127#_M1013_g N_A_605_563#_c_1076_n 0.0329256f $X=3.85 $Y=0.775
+ $X2=0.24 $Y2=0
cc_334 N_A_30_127#_c_229_n N_A_605_563#_c_1076_n 0.00605548f $X=4.66 $Y=2.585
+ $X2=0.24 $Y2=0
cc_335 N_A_30_127#_c_281_p N_A_605_563#_c_1076_n 0.0196874f $X=3.595 $Y=1.37
+ $X2=0.24 $Y2=0
cc_336 N_A_30_127#_c_229_n N_A_605_563#_c_1078_n 0.00907974f $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_337 N_A_30_127#_c_240_n N_A_605_563#_c_1078_n 0.0278367f $X=3.43 $Y=1.845
+ $X2=0 $Y2=0
cc_338 N_A_30_127#_c_240_n N_A_605_563#_c_1079_n 0.0267624f $X=3.43 $Y=1.845
+ $X2=11.76 $Y2=0
cc_339 N_A_30_127#_c_261_n N_A_605_563#_c_1079_n 0.00899259f $X=2.735 $Y=1.845
+ $X2=11.76 $Y2=0
cc_340 N_A_30_127#_M1013_g N_A_605_563#_c_1080_n 0.00368729f $X=3.85 $Y=0.775
+ $X2=0 $Y2=0
cc_341 N_A_30_127#_c_229_n N_A_605_563#_c_1080_n 0.0440164f $X=4.66 $Y=2.585
+ $X2=0 $Y2=0
cc_342 N_A_30_127#_c_240_n N_A_605_563#_c_1080_n 0.0126589f $X=3.43 $Y=1.845
+ $X2=0 $Y2=0
cc_343 N_A_30_127#_c_281_p N_A_605_563#_c_1080_n 0.0370533f $X=3.595 $Y=1.37
+ $X2=0 $Y2=0
cc_344 N_A_30_127#_M1004_g N_VGND_c_1129_n 0.0427478f $X=1.465 $Y=0.845 $X2=0
+ $Y2=0
cc_345 N_A_30_127#_c_235_n N_VGND_c_1129_n 0.00244799f $X=1.43 $Y=1.47 $X2=0
+ $Y2=0
cc_346 N_A_30_127#_c_236_n N_VGND_c_1129_n 0.0226208f $X=0.295 $Y=0.845 $X2=0
+ $Y2=0
cc_347 N_A_30_127#_c_239_n N_VGND_c_1129_n 0.0223123f $X=1.165 $Y=1.64 $X2=0
+ $Y2=0
cc_348 N_A_30_127#_c_286_p N_VGND_c_1129_n 0.00959694f $X=1.29 $Y=1.725 $X2=0
+ $Y2=0
cc_349 N_A_30_127#_M1004_g N_VGND_c_1131_n 0.00246028f $X=1.465 $Y=0.845 $X2=0
+ $Y2=0
cc_350 N_A_30_127#_M1002_g N_VGND_c_1135_n 0.00325409f $X=8.185 $Y=0.775 $X2=0
+ $Y2=0
cc_351 N_A_30_127#_M1004_g N_VGND_c_1139_n 0.012127f $X=1.465 $Y=0.845 $X2=0
+ $Y2=0
cc_352 N_A_30_127#_M1013_g N_VGND_c_1139_n 0.011508f $X=3.85 $Y=0.775 $X2=0
+ $Y2=0
cc_353 N_A_30_127#_c_229_n N_VGND_c_1139_n 0.00303117f $X=4.66 $Y=2.585 $X2=0
+ $Y2=0
cc_354 N_A_30_127#_M1002_g N_VGND_c_1139_n 0.0143441f $X=8.185 $Y=0.775 $X2=0
+ $Y2=0
cc_355 N_A_30_127#_c_236_n N_VGND_c_1139_n 0.0225738f $X=0.295 $Y=0.845 $X2=0
+ $Y2=0
cc_356 N_A_30_127#_c_281_p N_VGND_c_1139_n 8.84094e-19 $X=3.595 $Y=1.37 $X2=0
+ $Y2=0
cc_357 N_D_M1017_g N_A_339_559#_c_491_n 0.00312296f $X=2.775 $Y=3.025 $X2=0
+ $Y2=0
cc_358 N_D_c_424_n N_A_339_559#_c_491_n 0.0011424f $X=2.775 $Y=2.435 $X2=0 $Y2=0
cc_359 N_D_M1016_g N_A_339_559#_c_472_n 0.00505137f $X=2.95 $Y=0.775 $X2=11.76
+ $Y2=0
cc_360 N_D_c_424_n N_A_339_559#_c_494_n 0.040436f $X=2.775 $Y=2.435 $X2=0 $Y2=0
cc_361 N_D_M1016_g N_A_339_559#_c_474_n 0.015006f $X=2.95 $Y=0.775 $X2=0 $Y2=0
cc_362 N_D_c_419_n N_A_339_559#_c_474_n 0.0301749f $X=2.305 $Y=1.655 $X2=0 $Y2=0
cc_363 N_D_c_420_n N_A_339_559#_c_474_n 0.0337202f $X=2.95 $Y=1.59 $X2=0 $Y2=0
cc_364 N_D_c_419_n N_A_339_559#_c_475_n 0.0267662f $X=2.305 $Y=1.655 $X2=6 $Y2=0
cc_365 N_D_M1017_g N_A_339_559#_c_566_n 0.0255287f $X=2.775 $Y=3.025 $X2=6
+ $Y2=0.057
cc_366 N_D_c_424_n N_A_339_559#_c_566_n 0.00381022f $X=2.775 $Y=2.435 $X2=6
+ $Y2=0.057
cc_367 N_D_M1017_g N_A_339_559#_c_496_n 0.0136684f $X=2.775 $Y=3.025 $X2=6
+ $Y2=0.058
cc_368 N_D_M1017_g N_A_339_559#_c_499_n 0.00428284f $X=2.775 $Y=3.025 $X2=6
+ $Y2=0.058
cc_369 N_D_M1016_g N_A_339_559#_c_528_n 0.035257f $X=2.95 $Y=0.775 $X2=0 $Y2=0
cc_370 N_D_M1016_g N_A_339_559#_c_476_n 0.00341775f $X=2.95 $Y=0.775 $X2=0 $Y2=0
cc_371 N_D_M1016_g N_A_339_559#_c_478_n 0.00298755f $X=2.95 $Y=0.775 $X2=0 $Y2=0
cc_372 N_D_c_424_n N_A_339_559#_c_532_n 3.25894e-19 $X=2.775 $Y=2.435 $X2=0
+ $Y2=0
cc_373 N_D_c_424_n N_A_339_559#_c_502_n 0.0279784f $X=2.775 $Y=2.435 $X2=0 $Y2=0
cc_374 N_D_M1017_g N_A_339_559#_c_508_n 7.4616e-19 $X=2.775 $Y=3.025 $X2=0 $Y2=0
cc_375 N_D_M1017_g N_VPWR_c_1005_n 0.00501023f $X=2.775 $Y=3.025 $X2=0 $Y2=0
cc_376 N_D_c_424_n N_VPWR_c_1005_n 0.00730335f $X=2.775 $Y=2.435 $X2=0 $Y2=0
cc_377 N_D_M1017_g N_VPWR_c_1017_n 0.00417456f $X=2.775 $Y=3.025 $X2=0 $Y2=0
cc_378 N_D_M1017_g N_A_605_563#_c_1077_n 0.00926978f $X=2.775 $Y=3.025 $X2=0
+ $Y2=0
cc_379 N_D_c_424_n N_A_605_563#_c_1077_n 0.0172693f $X=2.775 $Y=2.435 $X2=0
+ $Y2=0
cc_380 N_D_M1016_g N_A_605_563#_c_1076_n 0.00433951f $X=2.95 $Y=0.775 $X2=0.24
+ $Y2=0
cc_381 N_D_c_424_n N_A_605_563#_c_1079_n 0.00581375f $X=2.775 $Y=2.435 $X2=11.76
+ $Y2=0
cc_382 N_D_c_420_n N_A_605_563#_c_1079_n 0.00117618f $X=2.95 $Y=1.59 $X2=11.76
+ $Y2=0
cc_383 N_D_M1016_g N_A_605_563#_c_1080_n 7.63366e-19 $X=2.95 $Y=0.775 $X2=0
+ $Y2=0
cc_384 N_D_M1016_g N_VGND_c_1131_n 0.0174126f $X=2.95 $Y=0.775 $X2=0 $Y2=0
cc_385 N_D_c_420_n N_VGND_c_1131_n 0.00279723f $X=2.95 $Y=1.59 $X2=0 $Y2=0
cc_386 N_D_M1016_g N_VGND_c_1139_n 0.0112688f $X=2.95 $Y=0.775 $X2=0 $Y2=0
cc_387 N_A_339_559#_c_504_n N_A_1024_371#_M1003_d 0.00388169f $X=7.485 $Y=3.22
+ $X2=0 $Y2=0
cc_388 N_A_339_559#_c_504_n N_A_1024_371#_M1006_g 0.0299555f $X=7.485 $Y=3.22
+ $X2=0 $Y2=0
cc_389 N_A_339_559#_c_542_n N_A_1024_371#_M1007_g 0.00202902f $X=4.89 $Y=1.175
+ $X2=0 $Y2=0
cc_390 N_A_339_559#_c_480_n N_A_1024_371#_M1007_g 0.0263986f $X=6.385 $Y=1.26
+ $X2=0 $Y2=0
cc_391 N_A_339_559#_c_580_p N_A_1024_371#_M1007_g 0.00133585f $X=6.47 $Y=1.175
+ $X2=0 $Y2=0
cc_392 N_A_339_559#_M1005_g N_A_1024_371#_M1007_g 0.0798812f $X=4.825 $Y=0.775
+ $X2=0 $Y2=0
cc_393 N_A_339_559#_c_480_n N_A_1024_371#_c_690_n 0.00614436f $X=6.385 $Y=1.26
+ $X2=0 $Y2=0
cc_394 N_A_339_559#_c_504_n N_A_1024_371#_c_703_n 0.0449398f $X=7.485 $Y=3.22
+ $X2=11.76 $Y2=0
cc_395 N_A_339_559#_c_480_n N_A_1024_371#_c_691_n 0.0129587f $X=6.385 $Y=1.26
+ $X2=6 $Y2=0.057
cc_396 N_A_339_559#_c_580_p N_A_1024_371#_c_691_n 0.0380955f $X=6.47 $Y=1.175
+ $X2=6 $Y2=0.057
cc_397 N_A_339_559#_c_481_n N_A_1024_371#_c_691_n 0.0210178f $X=7.28 $Y=0.35
+ $X2=6 $Y2=0.057
cc_398 N_A_339_559#_c_543_n N_A_1024_371#_c_691_n 0.031641f $X=7.365 $Y=1.125
+ $X2=6 $Y2=0.057
cc_399 N_A_339_559#_c_485_n N_A_1024_371#_c_691_n 0.0165649f $X=7.57 $Y=2.225
+ $X2=6 $Y2=0.057
cc_400 N_A_339_559#_c_486_n N_A_1024_371#_c_691_n 0.0213871f $X=7.57 $Y=1.285
+ $X2=6 $Y2=0.057
cc_401 N_A_339_559#_M1010_g N_A_1024_371#_c_691_n 0.00912891f $X=7.405 $Y=0.775
+ $X2=6 $Y2=0.057
cc_402 N_A_339_559#_c_485_n N_A_1024_371#_c_696_n 0.0116215f $X=7.57 $Y=2.225
+ $X2=0 $Y2=0
cc_403 N_A_339_559#_c_506_n N_A_1024_371#_c_696_n 0.0151051f $X=7.57 $Y=3.135
+ $X2=0 $Y2=0
cc_404 N_A_339_559#_c_551_n N_A_1024_371#_c_696_n 0.0210953f $X=7.57 $Y=2.37
+ $X2=0 $Y2=0
cc_405 N_A_339_559#_c_504_n N_A_1024_371#_c_692_n 0.00322853f $X=7.485 $Y=3.22
+ $X2=0 $Y2=0
cc_406 N_A_339_559#_c_485_n N_A_1024_371#_c_693_n 0.0122207f $X=7.57 $Y=2.225
+ $X2=0 $Y2=0
cc_407 N_A_339_559#_c_486_n N_A_1024_371#_c_693_n 8.4087e-19 $X=7.57 $Y=1.285
+ $X2=0 $Y2=0
cc_408 N_A_339_559#_M1010_g N_A_1024_371#_c_693_n 7.1046e-19 $X=7.405 $Y=0.775
+ $X2=0 $Y2=0
cc_409 N_A_339_559#_c_504_n N_A_780_574#_M1012_d 0.007508f $X=7.485 $Y=3.22
+ $X2=0 $Y2=0
cc_410 N_A_339_559#_c_504_n N_A_780_574#_M1003_g 0.0330955f $X=7.485 $Y=3.22
+ $X2=0 $Y2=0
cc_411 N_A_339_559#_c_480_n N_A_780_574#_c_758_n 0.0275485f $X=6.385 $Y=1.26
+ $X2=0.24 $Y2=0
cc_412 N_A_339_559#_c_580_p N_A_780_574#_c_758_n 0.0301024f $X=6.47 $Y=1.175
+ $X2=0.24 $Y2=0
cc_413 N_A_339_559#_c_481_n N_A_780_574#_c_758_n 0.0078963f $X=7.28 $Y=0.35
+ $X2=0.24 $Y2=0
cc_414 N_A_339_559#_c_483_n N_A_780_574#_c_758_n 0.00298755f $X=6.555 $Y=0.35
+ $X2=0.24 $Y2=0
cc_415 N_A_339_559#_c_543_n N_A_780_574#_c_758_n 0.00127013f $X=7.365 $Y=1.125
+ $X2=0.24 $Y2=0
cc_416 N_A_339_559#_M1010_g N_A_780_574#_c_758_n 0.0198276f $X=7.405 $Y=0.775
+ $X2=0.24 $Y2=0
cc_417 N_A_339_559#_c_476_n N_A_780_574#_c_760_n 0.0215508f $X=4.725 $Y=0.35
+ $X2=11.76 $Y2=0
cc_418 N_A_339_559#_c_542_n N_A_780_574#_c_760_n 0.0413632f $X=4.89 $Y=1.175
+ $X2=11.76 $Y2=0
cc_419 N_A_339_559#_M1005_g N_A_780_574#_c_760_n 0.00887723f $X=4.825 $Y=0.775
+ $X2=11.76 $Y2=0
cc_420 N_A_339_559#_c_542_n N_A_780_574#_c_761_n 0.024005f $X=4.89 $Y=1.175
+ $X2=0 $Y2=0
cc_421 N_A_339_559#_c_480_n N_A_780_574#_c_761_n 0.0876699f $X=6.385 $Y=1.26
+ $X2=0 $Y2=0
cc_422 N_A_339_559#_M1005_g N_A_780_574#_c_761_n 0.0207807f $X=4.825 $Y=0.775
+ $X2=0 $Y2=0
cc_423 N_A_339_559#_c_532_n N_A_780_574#_c_768_n 0.0182088f $X=3.675 $Y=2.545
+ $X2=0 $Y2=0
cc_424 N_A_339_559#_c_502_n N_A_780_574#_c_768_n 0.0030304f $X=3.675 $Y=2.545
+ $X2=0 $Y2=0
cc_425 N_A_339_559#_c_504_n N_A_780_574#_c_768_n 0.0225062f $X=7.485 $Y=3.22
+ $X2=0 $Y2=0
cc_426 N_A_339_559#_c_532_n N_A_780_574#_c_762_n 0.00845055f $X=3.675 $Y=2.545
+ $X2=0 $Y2=0
cc_427 N_A_339_559#_c_502_n N_A_780_574#_c_762_n 0.00232142f $X=3.675 $Y=2.545
+ $X2=0 $Y2=0
cc_428 N_A_339_559#_c_490_n N_A_1729_87#_M1015_g 0.0701214f $X=8.405 $Y=2.605
+ $X2=0 $Y2=0
cc_429 N_A_339_559#_c_490_n N_A_1729_87#_c_839_n 7.67108e-19 $X=8.405 $Y=2.605
+ $X2=0 $Y2=0
cc_430 N_A_339_559#_c_504_n N_A_1455_543#_M1020_d 0.01046f $X=7.485 $Y=3.22
+ $X2=0 $Y2=0
cc_431 N_A_339_559#_c_506_n N_A_1455_543#_M1020_d 0.0115048f $X=7.57 $Y=3.135
+ $X2=0 $Y2=0
cc_432 N_A_339_559#_c_490_n N_A_1455_543#_c_920_n 0.00491958f $X=8.405 $Y=2.605
+ $X2=0 $Y2=0
cc_433 N_A_339_559#_c_506_n N_A_1455_543#_c_920_n 0.0133151f $X=7.57 $Y=3.135
+ $X2=0 $Y2=0
cc_434 N_A_339_559#_c_507_n N_A_1455_543#_c_920_n 0.0202828f $X=8.085 $Y=2.39
+ $X2=0 $Y2=0
cc_435 N_A_339_559#_c_490_n N_A_1455_543#_c_921_n 0.0183504f $X=8.405 $Y=2.605
+ $X2=11.76 $Y2=0
cc_436 N_A_339_559#_c_504_n N_A_1455_543#_c_921_n 0.0136054f $X=7.485 $Y=3.22
+ $X2=11.76 $Y2=0
cc_437 N_A_339_559#_c_506_n N_A_1455_543#_c_921_n 0.0192822f $X=7.57 $Y=3.135
+ $X2=11.76 $Y2=0
cc_438 N_A_339_559#_c_490_n N_A_1455_543#_c_924_n 0.0292564f $X=8.405 $Y=2.605
+ $X2=6 $Y2=0
cc_439 N_A_339_559#_c_507_n N_A_1455_543#_c_924_n 0.0113668f $X=8.085 $Y=2.39
+ $X2=6 $Y2=0
cc_440 N_A_339_559#_c_490_n N_A_1455_543#_c_913_n 0.00620249f $X=8.405 $Y=2.605
+ $X2=6 $Y2=0.058
cc_441 N_A_339_559#_c_507_n N_A_1455_543#_c_913_n 0.00353187f $X=8.085 $Y=2.39
+ $X2=6 $Y2=0.058
cc_442 N_A_339_559#_c_490_n N_A_1455_543#_c_947_n 0.0153624f $X=8.405 $Y=2.605
+ $X2=0 $Y2=0
cc_443 N_A_339_559#_c_507_n N_A_1455_543#_c_947_n 0.00498672f $X=8.085 $Y=2.39
+ $X2=0 $Y2=0
cc_444 N_A_339_559#_c_490_n N_A_1455_543#_c_926_n 0.00654621f $X=8.405 $Y=2.605
+ $X2=0 $Y2=0
cc_445 N_A_339_559#_c_543_n N_A_1455_543#_c_914_n 0.0320668f $X=7.365 $Y=1.125
+ $X2=0 $Y2=0
cc_446 N_A_339_559#_c_486_n N_A_1455_543#_c_914_n 0.00172065f $X=7.57 $Y=1.285
+ $X2=0 $Y2=0
cc_447 N_A_339_559#_M1010_g N_A_1455_543#_c_914_n 0.00838965f $X=7.405 $Y=0.775
+ $X2=0 $Y2=0
cc_448 N_A_339_559#_c_490_n N_A_1455_543#_c_953_n 0.00525246f $X=8.405 $Y=2.605
+ $X2=0 $Y2=0
cc_449 N_A_339_559#_c_507_n N_A_1455_543#_c_953_n 0.0137383f $X=8.085 $Y=2.39
+ $X2=0 $Y2=0
cc_450 N_A_339_559#_c_504_n N_VPWR_M1006_d 0.00608368f $X=7.485 $Y=3.22 $X2=0
+ $Y2=0
cc_451 N_A_339_559#_c_491_n N_VPWR_c_1002_n 0.0597328f $X=1.835 $Y=2.94 $X2=0
+ $Y2=0
cc_452 N_A_339_559#_c_491_n N_VPWR_c_1005_n 0.0509425f $X=1.835 $Y=2.94 $X2=0
+ $Y2=0
cc_453 N_A_339_559#_c_494_n N_VPWR_c_1005_n 0.019167f $X=2.65 $Y=2.53 $X2=0
+ $Y2=0
cc_454 N_A_339_559#_c_566_n N_VPWR_c_1005_n 0.0198489f $X=2.735 $Y=3.305 $X2=0
+ $Y2=0
cc_455 N_A_339_559#_c_499_n N_VPWR_c_1005_n 0.0134523f $X=2.82 $Y=3.39 $X2=0
+ $Y2=0
cc_456 N_A_339_559#_c_504_n N_VPWR_c_1008_n 0.0557468f $X=7.485 $Y=3.22 $X2=0
+ $Y2=0
cc_457 N_A_339_559#_c_490_n N_VPWR_c_1011_n 0.00519298f $X=8.405 $Y=2.605 $X2=0
+ $Y2=0
cc_458 N_A_339_559#_c_490_n N_VPWR_c_1017_n 0.0156697f $X=8.405 $Y=2.605 $X2=0
+ $Y2=0
cc_459 N_A_339_559#_c_491_n N_VPWR_c_1017_n 0.0311182f $X=1.835 $Y=2.94 $X2=0
+ $Y2=0
cc_460 N_A_339_559#_c_496_n N_VPWR_c_1017_n 0.0303048f $X=3.51 $Y=3.39 $X2=0
+ $Y2=0
cc_461 N_A_339_559#_c_499_n N_VPWR_c_1017_n 0.00889212f $X=2.82 $Y=3.39 $X2=0
+ $Y2=0
cc_462 N_A_339_559#_c_502_n N_VPWR_c_1017_n 0.00757667f $X=3.675 $Y=2.545 $X2=0
+ $Y2=0
cc_463 N_A_339_559#_c_504_n N_VPWR_c_1017_n 0.170576f $X=7.485 $Y=3.22 $X2=0
+ $Y2=0
cc_464 N_A_339_559#_c_508_n N_VPWR_c_1017_n 0.018431f $X=3.675 $Y=3.22 $X2=0
+ $Y2=0
cc_465 N_A_339_559#_c_494_n N_A_605_563#_c_1077_n 0.0129587f $X=2.65 $Y=2.53
+ $X2=0 $Y2=0
cc_466 N_A_339_559#_c_566_n N_A_605_563#_c_1077_n 0.0346881f $X=2.735 $Y=3.305
+ $X2=0 $Y2=0
cc_467 N_A_339_559#_c_496_n N_A_605_563#_c_1077_n 0.021706f $X=3.51 $Y=3.39
+ $X2=0 $Y2=0
cc_468 N_A_339_559#_c_532_n N_A_605_563#_c_1077_n 0.0500187f $X=3.675 $Y=2.545
+ $X2=0 $Y2=0
cc_469 N_A_339_559#_c_502_n N_A_605_563#_c_1077_n 0.0120713f $X=3.675 $Y=2.545
+ $X2=0 $Y2=0
cc_470 N_A_339_559#_c_528_n N_A_605_563#_c_1076_n 0.030777f $X=3.03 $Y=1.205
+ $X2=0.24 $Y2=0
cc_471 N_A_339_559#_c_476_n N_A_605_563#_c_1076_n 0.0472258f $X=4.725 $Y=0.35
+ $X2=0.24 $Y2=0
cc_472 N_A_339_559#_c_532_n N_A_605_563#_c_1078_n 0.0238596f $X=3.675 $Y=2.545
+ $X2=0 $Y2=0
cc_473 N_A_339_559#_c_502_n N_A_605_563#_c_1078_n 0.0195082f $X=3.675 $Y=2.545
+ $X2=0 $Y2=0
cc_474 N_A_339_559#_c_480_n N_VGND_M1007_d 0.00417851f $X=6.385 $Y=1.26 $X2=0
+ $Y2=0
cc_475 N_A_339_559#_c_472_n N_VGND_c_1129_n 0.0375099f $X=1.855 $Y=0.845 $X2=0
+ $Y2=0
cc_476 N_A_339_559#_c_472_n N_VGND_c_1131_n 0.0354046f $X=1.855 $Y=0.845 $X2=0
+ $Y2=0
cc_477 N_A_339_559#_c_474_n N_VGND_c_1131_n 0.043781f $X=2.945 $Y=1.29 $X2=0
+ $Y2=0
cc_478 N_A_339_559#_c_528_n N_VGND_c_1131_n 0.0401114f $X=3.03 $Y=1.205 $X2=0
+ $Y2=0
cc_479 N_A_339_559#_c_478_n N_VGND_c_1131_n 0.00488507f $X=3.115 $Y=0.35 $X2=0
+ $Y2=0
cc_480 N_A_339_559#_c_476_n N_VGND_c_1133_n 0.00441475f $X=4.725 $Y=0.35 $X2=0
+ $Y2=0
cc_481 N_A_339_559#_c_542_n N_VGND_c_1133_n 0.0227166f $X=4.89 $Y=1.175 $X2=0
+ $Y2=0
cc_482 N_A_339_559#_c_480_n N_VGND_c_1133_n 0.0690271f $X=6.385 $Y=1.26 $X2=0
+ $Y2=0
cc_483 N_A_339_559#_c_580_p N_VGND_c_1133_n 0.0232834f $X=6.47 $Y=1.175 $X2=0
+ $Y2=0
cc_484 N_A_339_559#_c_483_n N_VGND_c_1133_n 0.00489946f $X=6.555 $Y=0.35 $X2=0
+ $Y2=0
cc_485 N_A_339_559#_M1005_g N_VGND_c_1133_n 0.00207121f $X=4.825 $Y=0.775 $X2=0
+ $Y2=0
cc_486 N_A_339_559#_c_472_n N_VGND_c_1139_n 0.0269193f $X=1.855 $Y=0.845 $X2=0
+ $Y2=0
cc_487 N_A_339_559#_c_474_n N_VGND_c_1139_n 0.0128829f $X=2.945 $Y=1.29 $X2=0
+ $Y2=0
cc_488 N_A_339_559#_c_528_n N_VGND_c_1139_n 0.0199794f $X=3.03 $Y=1.205 $X2=0
+ $Y2=0
cc_489 N_A_339_559#_c_476_n N_VGND_c_1139_n 0.0706587f $X=4.725 $Y=0.35 $X2=0
+ $Y2=0
cc_490 N_A_339_559#_c_478_n N_VGND_c_1139_n 0.00777234f $X=3.115 $Y=0.35 $X2=0
+ $Y2=0
cc_491 N_A_339_559#_c_542_n N_VGND_c_1139_n 0.0328837f $X=4.89 $Y=1.175 $X2=0
+ $Y2=0
cc_492 N_A_339_559#_c_480_n N_VGND_c_1139_n 0.0153945f $X=6.385 $Y=1.26 $X2=0
+ $Y2=0
cc_493 N_A_339_559#_c_580_p N_VGND_c_1139_n 0.0199629f $X=6.47 $Y=1.175 $X2=0
+ $Y2=0
cc_494 N_A_339_559#_c_481_n N_VGND_c_1139_n 0.0388381f $X=7.28 $Y=0.35 $X2=0
+ $Y2=0
cc_495 N_A_339_559#_c_483_n N_VGND_c_1139_n 0.00777234f $X=6.555 $Y=0.35 $X2=0
+ $Y2=0
cc_496 N_A_339_559#_c_543_n N_VGND_c_1139_n 0.015066f $X=7.365 $Y=1.125 $X2=0
+ $Y2=0
cc_497 N_A_339_559#_c_486_n N_VGND_c_1139_n 0.0061093f $X=7.57 $Y=1.285 $X2=0
+ $Y2=0
cc_498 N_A_339_559#_M1005_g N_VGND_c_1139_n 0.0112992f $X=4.825 $Y=0.775 $X2=0
+ $Y2=0
cc_499 N_A_339_559#_M1010_g N_VGND_c_1139_n 0.0141679f $X=7.405 $Y=0.775 $X2=0
+ $Y2=0
cc_500 N_A_1024_371#_M1006_g N_A_780_574#_M1003_g 0.0297323f $X=5.37 $Y=2.925
+ $X2=0 $Y2=0
cc_501 N_A_1024_371#_c_690_n N_A_780_574#_M1003_g 0.0198599f $X=6.735 $Y=1.96
+ $X2=0 $Y2=0
cc_502 N_A_1024_371#_c_703_n N_A_780_574#_M1003_g 0.0107706f $X=7.135 $Y=2.855
+ $X2=0 $Y2=0
cc_503 N_A_1024_371#_c_696_n N_A_780_574#_M1003_g 0.0014072f $X=7.22 $Y=2.755
+ $X2=0 $Y2=0
cc_504 N_A_1024_371#_c_709_n N_A_780_574#_M1003_g 0.00113699f $X=5.6 $Y=1.96
+ $X2=0 $Y2=0
cc_505 N_A_1024_371#_c_692_n N_A_780_574#_M1003_g 0.042473f $X=5.6 $Y=2.04 $X2=0
+ $Y2=0
cc_506 N_A_1024_371#_M1007_g N_A_780_574#_c_758_n 0.0669233f $X=5.535 $Y=0.775
+ $X2=0.24 $Y2=0
cc_507 N_A_1024_371#_c_690_n N_A_780_574#_c_758_n 0.0246121f $X=6.735 $Y=1.96
+ $X2=0.24 $Y2=0
cc_508 N_A_1024_371#_c_691_n N_A_780_574#_c_758_n 0.0437548f $X=6.9 $Y=0.7
+ $X2=0.24 $Y2=0
cc_509 N_A_1024_371#_c_693_n N_A_780_574#_c_758_n 6.41849e-19 $X=7.22 $Y=1.96
+ $X2=0.24 $Y2=0
cc_510 N_A_1024_371#_M1007_g N_A_780_574#_c_761_n 0.0311566f $X=5.535 $Y=0.775
+ $X2=0 $Y2=0
cc_511 N_A_1024_371#_c_690_n N_A_780_574#_c_761_n 0.039144f $X=6.735 $Y=1.96
+ $X2=0 $Y2=0
cc_512 N_A_1024_371#_c_691_n N_A_780_574#_c_761_n 0.00685575f $X=6.9 $Y=0.7
+ $X2=0 $Y2=0
cc_513 N_A_1024_371#_c_709_n N_A_780_574#_c_761_n 0.0224849f $X=5.6 $Y=1.96
+ $X2=0 $Y2=0
cc_514 N_A_1024_371#_c_692_n N_A_780_574#_c_761_n 0.00692299f $X=5.6 $Y=2.04
+ $X2=0 $Y2=0
cc_515 N_A_1024_371#_M1006_g N_VPWR_c_1008_n 0.00287831f $X=5.37 $Y=2.925 $X2=0
+ $Y2=0
cc_516 N_A_1024_371#_M1003_d N_VPWR_c_1017_n 0.00235311f $X=6.495 $Y=2.715 $X2=0
+ $Y2=0
cc_517 N_A_1024_371#_M1007_g N_VGND_c_1133_n 0.0515876f $X=5.535 $Y=0.775 $X2=0
+ $Y2=0
cc_518 N_A_1024_371#_M1021_d N_VGND_c_1139_n 0.00379508f $X=6.76 $Y=0.565 $X2=0
+ $Y2=0
cc_519 N_A_1024_371#_c_691_n N_VGND_c_1139_n 0.0227766f $X=6.9 $Y=0.7 $X2=0
+ $Y2=0
cc_520 N_A_780_574#_M1003_g N_VPWR_c_1008_n 0.00700108f $X=6.245 $Y=3.215 $X2=0
+ $Y2=0
cc_521 N_A_780_574#_M1003_g N_VPWR_c_1017_n 0.015854f $X=6.245 $Y=3.215 $X2=0
+ $Y2=0
cc_522 N_A_780_574#_c_760_n N_A_605_563#_c_1076_n 0.032229f $X=4.38 $Y=0.78
+ $X2=0.24 $Y2=0
cc_523 N_A_780_574#_c_762_n N_A_605_563#_c_1078_n 0.013138f $X=4.22 $Y=2.675
+ $X2=0 $Y2=0
cc_524 N_A_780_574#_c_760_n N_A_605_563#_c_1080_n 0.0343771f $X=4.38 $Y=0.78
+ $X2=0 $Y2=0
cc_525 N_A_780_574#_c_762_n N_A_605_563#_c_1080_n 0.0276095f $X=4.22 $Y=2.675
+ $X2=0 $Y2=0
cc_526 N_A_780_574#_c_763_n N_A_605_563#_c_1080_n 0.0123662f $X=4.38 $Y=1.61
+ $X2=0 $Y2=0
cc_527 N_A_780_574#_c_758_n N_VGND_c_1133_n 0.004926f $X=6.51 $Y=1.425 $X2=0
+ $Y2=0
cc_528 N_A_780_574#_M1013_d N_VGND_c_1139_n 0.00337793f $X=4.1 $Y=0.565 $X2=0
+ $Y2=0
cc_529 N_A_780_574#_c_758_n N_VGND_c_1139_n 0.0166345f $X=6.51 $Y=1.425 $X2=0
+ $Y2=0
cc_530 N_A_780_574#_c_760_n N_VGND_c_1139_n 0.0195569f $X=4.38 $Y=0.78 $X2=0
+ $Y2=0
cc_531 N_A_1729_87#_M1008_g N_A_1455_543#_M1019_g 0.00931748f $X=8.895 $Y=0.775
+ $X2=0 $Y2=0
cc_532 N_A_1729_87#_c_834_n N_A_1455_543#_M1019_g 0.021294f $X=10.18 $Y=1.51
+ $X2=0 $Y2=0
cc_533 N_A_1729_87#_c_835_n N_A_1455_543#_M1019_g 0.0319752f $X=10.345 $Y=0.69
+ $X2=0 $Y2=0
cc_534 N_A_1729_87#_c_837_n N_A_1455_543#_M1019_g 4.28593e-19 $X=10.38 $Y=2.005
+ $X2=0 $Y2=0
cc_535 N_A_1729_87#_c_839_n N_A_1455_543#_M1019_g 0.0185844f $X=9.165 $Y=1.51
+ $X2=0 $Y2=0
cc_536 N_A_1729_87#_c_860_p N_A_1455_543#_c_911_n 0.00219288f $X=9.165 $Y=1.85
+ $X2=0.24 $Y2=0
cc_537 N_A_1729_87#_c_834_n N_A_1455_543#_c_911_n 0.0205835f $X=10.18 $Y=1.51
+ $X2=0.24 $Y2=0
cc_538 N_A_1729_87#_c_837_n N_A_1455_543#_c_911_n 0.0229867f $X=10.38 $Y=2.005
+ $X2=0.24 $Y2=0
cc_539 N_A_1729_87#_c_845_n N_A_1455_543#_c_911_n 0.0166694f $X=10.38 $Y=2.86
+ $X2=0.24 $Y2=0
cc_540 N_A_1729_87#_c_839_n N_A_1455_543#_c_911_n 0.0305959f $X=9.165 $Y=1.51
+ $X2=0.24 $Y2=0
cc_541 N_A_1729_87#_c_840_n N_A_1455_543#_c_911_n 0.0326705f $X=11.085 $Y=1.835
+ $X2=0.24 $Y2=0
cc_542 N_A_1729_87#_M1015_g N_A_1455_543#_M1018_g 0.0198241f $X=9.115 $Y=2.925
+ $X2=0 $Y2=0
cc_543 N_A_1729_87#_c_845_n N_A_1455_543#_M1018_g 0.0414425f $X=10.38 $Y=2.86
+ $X2=0 $Y2=0
cc_544 N_A_1729_87#_M1008_g N_A_1455_543#_c_912_n 9.06764e-19 $X=8.895 $Y=0.775
+ $X2=0 $Y2=0
cc_545 N_A_1729_87#_M1008_g N_A_1455_543#_c_913_n 0.0125683f $X=8.895 $Y=0.775
+ $X2=6 $Y2=0.058
cc_546 N_A_1729_87#_M1015_g N_A_1455_543#_c_913_n 0.00781148f $X=9.115 $Y=2.925
+ $X2=6 $Y2=0.058
cc_547 N_A_1729_87#_c_871_p N_A_1455_543#_c_913_n 0.00711398f $X=9.165 $Y=1.595
+ $X2=6 $Y2=0.058
cc_548 N_A_1729_87#_c_860_p N_A_1455_543#_c_913_n 0.0165951f $X=9.165 $Y=1.85
+ $X2=6 $Y2=0.058
cc_549 N_A_1729_87#_M1015_g N_A_1455_543#_c_947_n 0.00163196f $X=9.115 $Y=2.925
+ $X2=0 $Y2=0
cc_550 N_A_1729_87#_M1015_g N_A_1455_543#_c_926_n 0.0332931f $X=9.115 $Y=2.925
+ $X2=0 $Y2=0
cc_551 N_A_1729_87#_c_860_p N_A_1455_543#_c_926_n 0.0175544f $X=9.165 $Y=1.85
+ $X2=0 $Y2=0
cc_552 N_A_1729_87#_c_845_n N_A_1455_543#_c_926_n 0.0129587f $X=10.38 $Y=2.86
+ $X2=0 $Y2=0
cc_553 N_A_1729_87#_c_839_n N_A_1455_543#_c_926_n 0.00798344f $X=9.165 $Y=1.51
+ $X2=0 $Y2=0
cc_554 N_A_1729_87#_c_860_p N_A_1455_543#_c_978_n 0.00953527f $X=9.165 $Y=1.85
+ $X2=0 $Y2=0
cc_555 N_A_1729_87#_c_834_n N_A_1455_543#_c_978_n 0.0238298f $X=10.18 $Y=1.51
+ $X2=0 $Y2=0
cc_556 N_A_1729_87#_c_837_n N_A_1455_543#_c_978_n 0.0175323f $X=10.38 $Y=2.005
+ $X2=0 $Y2=0
cc_557 N_A_1729_87#_c_845_n N_A_1455_543#_c_978_n 0.0192826f $X=10.38 $Y=2.86
+ $X2=0 $Y2=0
cc_558 N_A_1729_87#_c_839_n N_A_1455_543#_c_978_n 0.00284323f $X=9.165 $Y=1.51
+ $X2=0 $Y2=0
cc_559 N_A_1729_87#_M1008_g N_A_1455_543#_c_914_n 0.00124578f $X=8.895 $Y=0.775
+ $X2=0 $Y2=0
cc_560 N_A_1729_87#_M1015_g N_VPWR_c_1011_n 0.0569717f $X=9.115 $Y=2.925 $X2=0
+ $Y2=0
cc_561 N_A_1729_87#_c_845_n N_VPWR_c_1011_n 0.0325308f $X=10.38 $Y=2.86 $X2=0
+ $Y2=0
cc_562 N_A_1729_87#_M1009_g N_VPWR_c_1014_n 0.0645467f $X=11.335 $Y=2.965 $X2=0
+ $Y2=0
cc_563 N_A_1729_87#_c_845_n N_VPWR_c_1014_n 0.124474f $X=10.38 $Y=2.86 $X2=0
+ $Y2=0
cc_564 N_A_1729_87#_c_888_p N_VPWR_c_1014_n 0.0445218f $X=11.295 $Y=1.84 $X2=0
+ $Y2=0
cc_565 N_A_1729_87#_c_840_n N_VPWR_c_1014_n 0.0098749f $X=11.085 $Y=1.835 $X2=0
+ $Y2=0
cc_566 N_A_1729_87#_M1009_g N_VPWR_c_1017_n 0.01547f $X=11.335 $Y=2.965 $X2=0
+ $Y2=0
cc_567 N_A_1729_87#_c_845_n N_VPWR_c_1017_n 0.0404709f $X=10.38 $Y=2.86 $X2=0
+ $Y2=0
cc_568 N_A_1729_87#_M1023_g Q 0.030856f $X=11.335 $Y=1.08 $X2=0 $Y2=0
cc_569 N_A_1729_87#_c_888_p Q 0.0258106f $X=11.295 $Y=1.84 $X2=0 $Y2=0
cc_570 N_A_1729_87#_M1009_g Q 0.00529377f $X=11.335 $Y=2.965 $X2=0.24 $Y2=0
cc_571 N_A_1729_87#_M1009_g Q 0.0261682f $X=11.335 $Y=2.965 $X2=0 $Y2=0
cc_572 N_A_1729_87#_M1008_g N_VGND_c_1135_n 0.0731291f $X=8.895 $Y=0.775 $X2=0
+ $Y2=0
cc_573 N_A_1729_87#_c_871_p N_VGND_c_1135_n 0.0272246f $X=9.165 $Y=1.595 $X2=0
+ $Y2=0
cc_574 N_A_1729_87#_c_834_n N_VGND_c_1135_n 0.0290266f $X=10.18 $Y=1.51 $X2=0
+ $Y2=0
cc_575 N_A_1729_87#_c_835_n N_VGND_c_1135_n 0.0242648f $X=10.345 $Y=0.69 $X2=0
+ $Y2=0
cc_576 N_A_1729_87#_c_839_n N_VGND_c_1135_n 0.0067158f $X=9.165 $Y=1.51 $X2=0
+ $Y2=0
cc_577 N_A_1729_87#_M1023_g N_VGND_c_1137_n 0.0468575f $X=11.335 $Y=1.08 $X2=0
+ $Y2=0
cc_578 N_A_1729_87#_c_835_n N_VGND_c_1137_n 0.073746f $X=10.345 $Y=0.69 $X2=0
+ $Y2=0
cc_579 N_A_1729_87#_c_837_n N_VGND_c_1137_n 0.006204f $X=10.38 $Y=2.005 $X2=0
+ $Y2=0
cc_580 N_A_1729_87#_c_888_p N_VGND_c_1137_n 0.0465751f $X=11.295 $Y=1.84 $X2=0
+ $Y2=0
cc_581 N_A_1729_87#_c_840_n N_VGND_c_1137_n 0.0110338f $X=11.085 $Y=1.835 $X2=0
+ $Y2=0
cc_582 N_A_1729_87#_M1008_g N_VGND_c_1139_n 0.00886702f $X=8.895 $Y=0.775 $X2=0
+ $Y2=0
cc_583 N_A_1729_87#_M1023_g N_VGND_c_1139_n 0.0187561f $X=11.335 $Y=1.08 $X2=0
+ $Y2=0
cc_584 N_A_1729_87#_c_835_n N_VGND_c_1139_n 0.030995f $X=10.345 $Y=0.69 $X2=0
+ $Y2=0
cc_585 N_A_1455_543#_c_911_n N_VPWR_c_1011_n 0.00145793f $X=9.99 $Y=2.465 $X2=0
+ $Y2=0
cc_586 N_A_1455_543#_M1018_g N_VPWR_c_1011_n 0.0270513f $X=9.99 $Y=3.215 $X2=0
+ $Y2=0
cc_587 N_A_1455_543#_c_924_n N_VPWR_c_1011_n 0.00667962f $X=8.43 $Y=2.78 $X2=0
+ $Y2=0
cc_588 N_A_1455_543#_c_926_n N_VPWR_c_1011_n 0.0567394f $X=9.705 $Y=2.36 $X2=0
+ $Y2=0
cc_589 N_A_1455_543#_c_911_n N_VPWR_c_1014_n 0.0036694f $X=9.99 $Y=2.465 $X2=0
+ $Y2=0
cc_590 N_A_1455_543#_M1020_d N_VPWR_c_1017_n 0.0132914f $X=7.275 $Y=2.715 $X2=0
+ $Y2=0
cc_591 N_A_1455_543#_M1018_g N_VPWR_c_1017_n 0.0283383f $X=9.99 $Y=3.215 $X2=0
+ $Y2=0
cc_592 N_A_1455_543#_c_921_n N_VPWR_c_1017_n 0.043012f $X=7.92 $Y=3.215 $X2=0
+ $Y2=0
cc_593 N_A_1455_543#_c_924_n N_VPWR_c_1017_n 0.0166808f $X=8.43 $Y=2.78 $X2=0
+ $Y2=0
cc_594 N_A_1455_543#_M1019_g N_VGND_c_1135_n 0.0252328f $X=9.955 $Y=0.94 $X2=0
+ $Y2=0
cc_595 N_A_1455_543#_c_912_n N_VGND_c_1135_n 0.00858417f $X=8.43 $Y=0.94 $X2=0
+ $Y2=0
cc_596 N_A_1455_543#_c_913_n N_VGND_c_1135_n 0.0167237f $X=8.515 $Y=2.275 $X2=0
+ $Y2=0
cc_597 N_A_1455_543#_M1019_g N_VGND_c_1137_n 0.00379188f $X=9.955 $Y=0.94 $X2=0
+ $Y2=0
cc_598 N_A_1455_543#_c_911_n N_VGND_c_1137_n 2.13991e-19 $X=9.99 $Y=2.465 $X2=0
+ $Y2=0
cc_599 N_A_1455_543#_M1019_g N_VGND_c_1139_n 0.0292045f $X=9.955 $Y=0.94 $X2=0
+ $Y2=0
cc_600 N_A_1455_543#_c_912_n N_VGND_c_1139_n 0.0258996f $X=8.43 $Y=0.94 $X2=0
+ $Y2=0
cc_601 N_A_1455_543#_c_914_n N_VGND_c_1139_n 0.0316806f $X=7.795 $Y=0.775 $X2=0
+ $Y2=0
cc_602 N_A_1455_543#_c_912_n A_1687_113# 0.00156314f $X=8.43 $Y=0.94 $X2=0 $Y2=0
cc_603 N_VPWR_c_1017_n N_A_605_563#_c_1077_n 0.00196592f $X=11.2 $Y=3.59
+ $X2=0.24 $Y2=4.07
cc_604 N_VPWR_c_1014_n Q 0.085876f $X=10.945 $Y=2.36 $X2=0 $Y2=0
cc_605 N_VPWR_c_1017_n Q 0.0425942f $X=11.2 $Y=3.59 $X2=0 $Y2=0
cc_606 N_A_605_563#_M1016_d N_VGND_c_1139_n 0.0039619f $X=3.2 $Y=0.565 $X2=0
+ $Y2=0
cc_607 N_A_605_563#_c_1076_n N_VGND_c_1139_n 0.0390958f $X=3.865 $Y=0.82 $X2=0
+ $Y2=0
cc_608 Q N_VGND_c_1137_n 0.0195601f $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_609 Q N_VGND_c_1139_n 0.0109542f $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_610 N_VGND_c_1139_n A_1015_113# 0.00244025f $X=11.165 $Y=0.48 $X2=0 $Y2=0
cc_611 N_VGND_c_1139_n A_1687_113# 0.00340398f $X=11.165 $Y=0.48 $X2=0 $Y2=0
