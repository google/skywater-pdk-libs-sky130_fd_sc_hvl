* File: sky130_fd_sc_hvl__lsbufhv2hv_lh_1.pex.spice
* Created: Wed Sep  2 09:07:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%VNB 9 11 12 23 35 42 49
r77 29 49 2.92572 $w=2.3e-07 $l=4.56e-06 $layer=MET1_cond $X=0.24 $Y=8.14
+ $X2=4.8 $Y2=8.14
r78 17 42 2.92572 $w=2.3e-07 $l=4.56e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.8
+ $Y2=0
r79 12 35 3.23369 $w=2.3e-07 $l=5.04e-06 $layer=MET1_cond $X=5.28 $Y=8.14
+ $X2=10.32 $Y2=8.14
r80 12 49 0.30797 $w=2.3e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=8.14 $X2=4.8
+ $Y2=8.14
r81 11 23 3.23369 $w=2.3e-07 $l=5.04e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=10.32
+ $Y2=0
r82 11 42 0.30797 $w=2.3e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=0 $X2=4.8
+ $Y2=0
r83 9 35 0.845455 $w=1.7e-07 $l=1.87e-06 $layer=mcon $count=11 $X=10.32 $Y=8.14
+ $X2=10.32 $Y2=8.14
r84 9 29 0.845455 $w=1.7e-07 $l=1.87e-06 $layer=mcon $count=11 $X=0.24 $Y=8.14
+ $X2=0.24 $Y2=8.14
r85 9 23 0.845455 $w=1.7e-07 $l=1.87e-06 $layer=mcon $count=11 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r86 9 17 0.845455 $w=1.7e-07 $l=1.87e-06 $layer=mcon $count=11 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%VPB 7 8 11 14 25 26 32
r58 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=4.07
+ $X2=10.32 $Y2=4.07
r59 21 26 0.92391 $w=2.3e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=4.07
+ $X2=10.32 $Y2=4.07
r60 20 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=4.07
+ $X2=10.32 $Y2=4.07
r61 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=4.07
+ $X2=8.88 $Y2=4.07
r62 15 32 2.92572 $w=2.3e-07 $l=4.56e-06 $layer=MET1_cond $X=0.24 $Y=4.07
+ $X2=4.8 $Y2=4.07
r63 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r64 11 21 2.30978 $w=2.3e-07 $l=3.6e-06 $layer=MET1_cond $X=5.28 $Y=4.07
+ $X2=8.88 $Y2=4.07
r65 11 32 0.30797 $w=2.3e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=4.07 $X2=4.8
+ $Y2=4.07
r66 8 25 91 $w=1.7e-07 $l=1.68696e-06 $layer=licon1_NTAP_notbjt $count=2
+ $X=8.675 $Y=3.985 $X2=10.32 $Y2=4.07
r67 8 20 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=8.675 $Y=3.985 $X2=8.88 $Y2=4.07
r68 7 14 182 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=1 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%LOWHVPWR 1 7 15 17 20 28
r48 24 28 0.291566 $w=2.85e-07 $l=5.85e-07 $layer=MET1_cond $X=4.215 $Y=3.162
+ $X2=4.8 $Y2=3.162
r49 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.215 $Y=3.135
+ $X2=4.215 $Y2=3.135
r50 20 23 13.0758 $w=5.88e-07 $l=6.45e-07 $layer=LI1_cond $X=4.035 $Y=2.49
+ $X2=4.035 $Y2=3.135
r51 17 28 0.239234 $w=2.85e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=3.162
+ $X2=4.8 $Y2=3.162
r52 13 23 4.45995 $w=5.88e-07 $l=2.2e-07 $layer=LI1_cond $X=4.035 $Y=3.355
+ $X2=4.035 $Y2=3.135
r53 12 15 11.7823 $w=6.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.035 $Y=3.69
+ $X2=4.695 $Y2=3.69
r54 12 13 1.48065 $w=5.9e-07 $l=3.35e-07 $layer=LI1_cond $X=4.035 $Y=3.69
+ $X2=4.035 $Y2=3.355
r55 10 12 6.42669 $w=6.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.675 $Y=3.69
+ $X2=4.035 $Y2=3.69
r56 7 15 45.5 $w=1.7e-07 $l=1.6263e-06 $layer=licon1_NTAP_notbjt $count=4
+ $X=3.13 $Y=3.395 $X2=4.695 $Y2=3.52
r57 7 10 45.5 $w=1.7e-07 $l=6.04276e-07 $layer=licon1_NTAP_notbjt $count=4
+ $X=3.13 $Y=3.395 $X2=3.675 $Y2=3.52
r58 1 20 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.895
+ $Y=2.345 $X2=4.035 $Y2=2.49
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A 1 5 9 11 12 13 17
r33 17 20 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.66 $Y=1.695
+ $X2=2.66 $Y2=1.87
r34 12 13 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.65 $Y=1.665
+ $X2=2.65 $Y2=2.035
r35 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.66
+ $Y=1.695 $X2=2.66 $Y2=1.695
r36 7 11 14.2643 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.645 $Y=2.035
+ $X2=3.645 $Y2=1.87
r37 7 9 73.299 $w=5e-07 $l=6.85e-07 $layer=POLY_cond $X=3.645 $Y=2.035 $X2=3.645
+ $Y2=2.72
r38 3 11 14.2643 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.645 $Y=1.705
+ $X2=3.645 $Y2=1.87
r39 3 5 66.8787 $w=5e-07 $l=6.25e-07 $layer=POLY_cond $X=3.645 $Y=1.705
+ $X2=3.645 $Y2=1.08
r40 2 20 2.83073 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.825 $Y=1.87
+ $X2=2.66 $Y2=1.87
r41 1 11 11.3528 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.395 $Y=1.87
+ $X2=3.645 $Y2=1.87
r42 1 2 99.6709 $w=3.3e-07 $l=5.7e-07 $layer=POLY_cond $X=3.395 $Y=1.87
+ $X2=2.825 $Y2=1.87
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A_626_141# 1 2 7 9 12 16 18 20 21
+ 23 24 26 29 34 37 38 40 45 48 56
r95 46 56 4.75345 $w=5.07e-07 $l=5e-08 $layer=POLY_cond $X=5.495 $Y=5.58
+ $X2=5.545 $Y2=5.58
r96 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.495
+ $Y=5.33 $X2=5.495 $Y2=5.33
r97 43 46 64.6469 $w=5.07e-07 $l=6.8e-07 $layer=POLY_cond $X=4.815 $Y=5.58
+ $X2=5.495 $Y2=5.58
r98 43 53 4.75345 $w=5.07e-07 $l=5e-08 $layer=POLY_cond $X=4.815 $Y=5.58
+ $X2=4.765 $Y2=5.58
r99 42 45 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.815 $Y=5.33
+ $X2=5.495 $Y2=5.33
r100 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.815
+ $Y=5.33 $X2=4.815 $Y2=5.33
r101 40 42 48.7169 $w=3.28e-07 $l=1.395e-06 $layer=LI1_cond $X=3.42 $Y=5.33
+ $X2=4.815 $Y2=5.33
r102 38 51 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.51 $Y=1.87
+ $X2=4.51 $Y2=2.035
r103 38 50 16.7369 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.51 $Y=1.87
+ $X2=4.51 $Y2=1.705
r104 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.68
+ $Y=1.87 $X2=4.68 $Y2=1.87
r105 35 48 2.3589 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.42 $Y=1.87
+ $X2=3.255 $Y2=1.87
r106 35 37 58.0831 $w=2.48e-07 $l=1.26e-06 $layer=LI1_cond $X=3.42 $Y=1.87
+ $X2=4.68 $Y2=1.87
r107 32 40 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=3.255 $Y=5.165
+ $X2=3.42 $Y2=5.33
r108 32 34 93.4177 $w=3.28e-07 $l=2.675e-06 $layer=LI1_cond $X=3.255 $Y=5.165
+ $X2=3.255 $Y2=2.49
r109 31 48 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=3.255 $Y=1.995
+ $X2=3.255 $Y2=1.87
r110 31 34 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.255 $Y=1.995
+ $X2=3.255 $Y2=2.49
r111 27 48 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=3.255 $Y=1.745
+ $X2=3.255 $Y2=1.87
r112 27 29 31.2557 $w=3.28e-07 $l=8.95e-07 $layer=LI1_cond $X=3.255 $Y=1.745
+ $X2=3.255 $Y2=0.85
r113 24 56 74.1538 $w=5.07e-07 $l=9.65453e-07 $layer=POLY_cond $X=6.325 $Y=5.995
+ $X2=5.545 $Y2=5.58
r114 24 26 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.325 $Y=5.995
+ $X2=6.325 $Y2=6.855
r115 21 56 3.16516 $w=5e-07 $l=4.15e-07 $layer=POLY_cond $X=5.545 $Y=5.995
+ $X2=5.545 $Y2=5.58
r116 21 23 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.545 $Y=5.995
+ $X2=5.545 $Y2=6.855
r117 18 53 3.16516 $w=5e-07 $l=4.15e-07 $layer=POLY_cond $X=4.765 $Y=5.995
+ $X2=4.765 $Y2=5.58
r118 18 20 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.765 $Y=5.995
+ $X2=4.765 $Y2=6.855
r119 16 51 73.299 $w=5e-07 $l=6.85e-07 $layer=POLY_cond $X=4.425 $Y=2.72
+ $X2=4.425 $Y2=2.035
r120 12 50 66.8787 $w=5e-07 $l=6.25e-07 $layer=POLY_cond $X=4.425 $Y=1.08
+ $X2=4.425 $Y2=1.705
r121 7 53 74.1538 $w=5.07e-07 $l=9.65453e-07 $layer=POLY_cond $X=3.985 $Y=5.995
+ $X2=4.765 $Y2=5.58
r122 7 9 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.985 $Y=5.995 $X2=3.985
+ $Y2=6.855
r123 2 34 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.345 $X2=3.255 $Y2=2.49
r124 1 29 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.705 $X2=3.255 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A_847_1221# 1 2 3 11 15 17 20 24 25
+ 28 32 37 38 42
r61 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.88
+ $Y=3.77 $X2=7.88 $Y2=3.77
r62 39 42 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=7.765 $Y=3.77
+ $X2=7.88 $Y2=3.77
r63 35 37 38.2402 $w=3.28e-07 $l=1.095e-06 $layer=LI1_cond $X=7.765 $Y=5.665
+ $X2=7.765 $Y2=4.57
r64 34 39 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.765 $Y=3.935
+ $X2=7.765 $Y2=3.77
r65 34 37 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=7.765 $Y=3.935
+ $X2=7.765 $Y2=4.57
r66 33 38 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.1 $Y=5.83
+ $X2=5.935 $Y2=5.83
r67 32 35 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=7.6 $Y=5.83
+ $X2=7.765 $Y2=5.665
r68 32 33 52.3838 $w=3.28e-07 $l=1.5e-06 $layer=LI1_cond $X=7.6 $Y=5.83 $X2=6.1
+ $Y2=5.83
r69 28 30 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=5.935 $Y=6.25
+ $X2=5.935 $Y2=7.46
r70 26 38 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.935 $Y=5.995
+ $X2=5.935 $Y2=5.83
r71 26 28 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.935 $Y=5.995
+ $X2=5.935 $Y2=6.25
r72 24 38 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.77 $Y=5.83
+ $X2=5.935 $Y2=5.83
r73 24 25 42.9547 $w=3.28e-07 $l=1.23e-06 $layer=LI1_cond $X=5.77 $Y=5.83
+ $X2=4.54 $Y2=5.83
r74 20 22 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=4.375 $Y=6.25
+ $X2=4.375 $Y2=7.46
r75 18 25 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=4.375 $Y=5.995
+ $X2=4.54 $Y2=5.83
r76 18 20 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.375 $Y=5.995
+ $X2=4.375 $Y2=6.25
r77 17 43 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=7.965 $Y=3.77
+ $X2=7.88 $Y2=3.77
r78 12 15 26.3581 $w=6.8e-07 $l=3.35e-07 $layer=POLY_cond $X=8.13 $Y=3.025
+ $X2=8.465 $Y2=3.025
r79 11 17 26.9307 $w=3.3e-07 $l=2.33345e-07 $layer=POLY_cond $X=8.13 $Y=3.605
+ $X2=7.965 $Y2=3.77
r80 10 12 19.6718 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.13 $Y=3.365
+ $X2=8.13 $Y2=3.025
r81 10 11 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=8.13 $Y=3.365
+ $X2=8.13 $Y2=3.605
r82 3 37 300 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=2 $X=7.6
+ $Y=4.425 $X2=7.825 $Y2=4.57
r83 2 30 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=5.795
+ $Y=6.105 $X2=5.935 $Y2=7.46
r84 2 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.795
+ $Y=6.105 $X2=5.935 $Y2=6.25
r85 1 22 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=4.235
+ $Y=6.105 $X2=4.375 $Y2=7.46
r86 1 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.235
+ $Y=6.105 $X2=4.375 $Y2=6.25
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A_935_141# 1 2 7 9 10 12 13 15 16
+ 18 21 25 27 28 29 30 32 38 41 42
r77 39 42 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=6.405 $Y=2.31
+ $X2=6.265 $Y2=2.31
r78 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.405
+ $Y=2.31 $X2=6.405 $Y2=2.31
r79 36 42 94.4251 $w=3.3e-07 $l=5.4e-07 $layer=POLY_cond $X=5.725 $Y=2.31
+ $X2=6.265 $Y2=2.31
r80 35 38 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.725 $Y=2.31
+ $X2=6.405 $Y2=2.31
r81 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.725
+ $Y=2.31 $X2=5.725 $Y2=2.31
r82 33 41 5.29963 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.66 $Y=2.31
+ $X2=5.495 $Y2=2.31
r83 33 35 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=5.66 $Y=2.31
+ $X2=5.725 $Y2=2.31
r84 32 41 1.23199 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=5.495 $Y=2.145
+ $X2=5.495 $Y2=2.31
r85 31 32 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=5.495 $Y=1.475
+ $X2=5.495 $Y2=2.145
r86 29 41 5.29963 $w=3.2e-07 $l=1.69926e-07 $layer=LI1_cond $X=5.33 $Y=2.32
+ $X2=5.495 $Y2=2.31
r87 29 30 13.0115 $w=3.08e-07 $l=3.5e-07 $layer=LI1_cond $X=5.33 $Y=2.32
+ $X2=4.98 $Y2=2.32
r88 27 31 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=5.33 $Y=1.31
+ $X2=5.495 $Y2=1.475
r89 27 28 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=5.33 $Y=1.31
+ $X2=4.98 $Y2=1.31
r90 23 30 6.82515 $w=3.1e-07 $l=2.29783e-07 $layer=LI1_cond $X=4.815 $Y=2.475
+ $X2=4.98 $Y2=2.32
r91 23 25 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.815 $Y=2.475
+ $X2=4.815 $Y2=2.49
r92 19 28 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=4.815 $Y=1.145
+ $X2=4.98 $Y2=1.31
r93 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.815 $Y=1.145
+ $X2=4.815 $Y2=0.85
r94 16 18 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.855 $Y=2.145
+ $X2=8.855 $Y2=1.285
r95 13 16 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=8.075 $Y=2.31
+ $X2=8.855 $Y2=2.31
r96 13 15 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.075 $Y=2.145
+ $X2=8.075 $Y2=1.285
r97 10 13 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=7.295 $Y=2.31
+ $X2=8.075 $Y2=2.31
r98 10 12 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.295 $Y=2.145
+ $X2=7.295 $Y2=1.285
r99 7 10 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=6.515 $Y=2.31
+ $X2=7.295 $Y2=2.31
r100 7 39 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=6.515 $Y=2.31
+ $X2=6.405 $Y2=2.31
r101 7 9 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.515 $Y=2.145 $X2=6.515
+ $Y2=1.285
r102 2 25 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.675
+ $Y=2.345 $X2=4.815 $Y2=2.49
r103 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.675
+ $Y=0.705 $X2=4.815 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%A_1353_107# 1 2 3 10 14 18 21 23 26
+ 29 33 34 36 37 38 41 47 53 57 58 60
r88 58 60 149.506 $w=3.3e-07 $l=8.55e-07 $layer=POLY_cond $X=8.8 $Y=5.37 $X2=8.8
+ $Y2=6.225
r89 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.8 $Y=5.37
+ $X2=8.8 $Y2=5.37
r90 54 57 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=8.38 $Y=5.37 $X2=8.8
+ $Y2=5.37
r91 48 60 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.8 $Y=6.39 $X2=8.8
+ $Y2=6.225
r92 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.8 $Y=6.39
+ $X2=8.8 $Y2=6.39
r93 45 57 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.8 $Y=5.535
+ $X2=8.8 $Y2=5.37
r94 45 47 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=8.8 $Y=5.535
+ $X2=8.8 $Y2=6.39
r95 41 44 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=8.465 $Y=0.68
+ $X2=8.465 $Y2=1.89
r96 39 53 5.16603 $w=3.3e-07 $l=1.85257e-07 $layer=LI1_cond $X=8.465 $Y=2.145
+ $X2=8.422 $Y2=2.31
r97 39 44 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=8.465 $Y=2.145
+ $X2=8.465 $Y2=1.89
r98 38 54 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.38 $Y=5.205
+ $X2=8.38 $Y2=5.37
r99 37 51 15.4589 $w=4.38e-07 $l=5.55e-07 $layer=LI1_cond $X=8.38 $Y=3.115
+ $X2=7.825 $Y2=3.115
r100 37 38 72.6388 $w=3.28e-07 $l=2.08e-06 $layer=LI1_cond $X=8.38 $Y=3.125
+ $X2=8.38 $Y2=5.205
r101 36 37 2.3974 $w=3.3e-07 $l=3.2e-07 $layer=LI1_cond $X=8.38 $Y=2.795
+ $X2=8.38 $Y2=3.115
r102 35 53 5.16603 $w=3.3e-07 $l=1.84811e-07 $layer=LI1_cond $X=8.38 $Y=2.475
+ $X2=8.422 $Y2=2.31
r103 35 36 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=8.38 $Y=2.475
+ $X2=8.38 $Y2=2.795
r104 33 53 1.34256 $w=3.3e-07 $l=2.07e-07 $layer=LI1_cond $X=8.215 $Y=2.31
+ $X2=8.422 $Y2=2.31
r105 33 34 39.9863 $w=3.28e-07 $l=1.145e-06 $layer=LI1_cond $X=8.215 $Y=2.31
+ $X2=7.07 $Y2=2.31
r106 29 32 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=6.905 $Y=0.68
+ $X2=6.905 $Y2=1.89
r107 27 34 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=6.905 $Y=2.145
+ $X2=7.07 $Y2=2.31
r108 27 32 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.905 $Y=2.145
+ $X2=6.905 $Y2=1.89
r109 24 58 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=8.8 $Y=4.975
+ $X2=8.8 $Y2=5.37
r110 23 24 19.6718 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.8 $Y=4.635
+ $X2=8.8 $Y2=4.975
r111 21 23 26.3581 $w=6.8e-07 $l=3.35e-07 $layer=POLY_cond $X=8.465 $Y=4.635
+ $X2=8.8 $Y2=4.635
r112 16 26 14.2643 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.895 $Y=6.555
+ $X2=9.895 $Y2=6.39
r113 16 18 72.229 $w=5e-07 $l=6.75e-07 $layer=POLY_cond $X=9.895 $Y=6.555
+ $X2=9.895 $Y2=7.23
r114 12 26 14.2643 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.895 $Y=6.225
+ $X2=9.895 $Y2=6.39
r115 12 14 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=9.895 $Y=6.225
+ $X2=9.895 $Y2=5.175
r116 11 48 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.965 $Y=6.39
+ $X2=8.8 $Y2=6.39
r117 10 26 11.3528 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=9.645 $Y=6.39
+ $X2=9.895 $Y2=6.39
r118 10 11 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=9.645 $Y=6.39
+ $X2=8.965 $Y2=6.39
r119 3 51 300 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=2 $X=7.6
+ $Y=2.815 $X2=7.825 $Y2=2.96
r120 2 44 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=8.325
+ $Y=0.535 $X2=8.465 $Y2=1.89
r121 2 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.325
+ $Y=0.535 $X2=8.465 $Y2=0.68
r122 1 32 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.535 $X2=6.905 $Y2=1.89
r123 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.535 $X2=6.905 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%VPWR 1 2 7 9 13 14 17 23 27 31 34
+ 40
r67 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.685 $Y=4.58
+ $X2=9.685 $Y2=4.58
r68 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.415 $Y=3.56
+ $X2=9.415 $Y2=3.56
r69 23 26 12.1635 $w=5.88e-07 $l=6e-07 $layer=LI1_cond $X=9.235 $Y=2.96
+ $X2=9.235 $Y2=3.56
r70 20 31 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.965 $Y=4.51
+ $X2=9.685 $Y2=4.51
r71 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.965 $Y=4.58
+ $X2=8.965 $Y2=4.58
r72 17 30 4.29026 $w=3.95e-07 $l=2.95e-07 $layer=LI1_cond $X=9.21 $Y=4.602
+ $X2=9.505 $Y2=4.602
r73 17 19 7.14806 $w=3.93e-07 $l=2.45e-07 $layer=LI1_cond $X=9.21 $Y=4.602
+ $X2=8.965 $Y2=4.602
r74 14 20 1.41469 $w=3.7e-07 $l=3.685e-06 $layer=MET1_cond $X=5.28 $Y=4.51
+ $X2=8.965 $Y2=4.51
r75 14 40 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=4.51
+ $X2=4.8 $Y2=4.51
r76 13 27 1.58745 $w=3.7e-07 $l=4.135e-06 $layer=MET1_cond $X=5.28 $Y=3.63
+ $X2=9.415 $Y2=3.63
r77 13 34 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=3.63
+ $X2=4.8 $Y2=3.63
r78 9 11 16.4207 $w=5.88e-07 $l=8.1e-07 $layer=LI1_cond $X=9.505 $Y=4.97
+ $X2=9.505 $Y2=5.78
r79 7 30 2.87956 $w=5.9e-07 $l=1.98e-07 $layer=LI1_cond $X=9.505 $Y=4.8
+ $X2=9.505 $Y2=4.602
r80 7 9 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=9.505 $Y=4.8 $X2=9.505
+ $Y2=4.97
r81 2 30 300 $w=1.7e-07 $l=6.08194e-07 $layer=licon1_PDIFF $count=2 $X=8.965
+ $Y=4.425 $X2=9.505 $Y2=4.57
r82 2 11 400 $w=1.7e-07 $l=1.60241e-06 $layer=licon1_PDIFF $count=1 $X=8.965
+ $Y=4.425 $X2=9.505 $Y2=5.78
r83 2 9 400 $w=1.7e-07 $l=7.68977e-07 $layer=licon1_PDIFF $count=1 $X=8.965
+ $Y=4.425 $X2=9.505 $Y2=4.97
r84 1 23 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.965
+ $Y=2.815 $X2=9.105 $Y2=2.96
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%X 1 2 7 8 9 10 11 18
r13 11 32 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=10.285 $Y=6.845
+ $X2=10.285 $Y2=7
r14 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.285 $Y=6.475
+ $X2=10.285 $Y2=6.845
r15 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.285 $Y=6.105
+ $X2=10.285 $Y2=6.475
r16 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.285 $Y=5.735
+ $X2=10.285 $Y2=6.105
r17 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.285 $Y=5.365
+ $X2=10.285 $Y2=5.735
r18 7 18 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=10.285 $Y=5.365
+ $X2=10.285 $Y2=4.57
r19 2 8 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=10.145
+ $Y=4.425 $X2=10.285 $Y2=5.78
r20 2 18 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=10.145
+ $Y=4.425 $X2=10.285 $Y2=4.57
r21 1 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.145
+ $Y=6.855 $X2=10.285 $Y2=7
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2HV_LH_1%VGND 1 2 3 4 5 6 7 8 25 26 27 28 29
+ 31 33 38 40 43 45 46 50 58 64 72 80 88 96 97 104 108 113 122
r113 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.685 $Y=7.63
+ $X2=9.685 $Y2=7.63
r114 104 107 12.7717 $w=5.88e-07 $l=6.3e-07 $layer=LI1_cond $X=9.505 $Y=7
+ $X2=9.505 $Y2=7.63
r115 99 101 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=9.245 $Y=0.68
+ $X2=9.245 $Y2=1.89
r116 96 99 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=9.245 $Y=0.51
+ $X2=9.245 $Y2=0.68
r117 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.425 $Y=0.51
+ $X2=9.425 $Y2=0.51
r118 91 93 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=7.685 $Y=0.68
+ $X2=7.685 $Y2=1.89
r119 89 97 0.598892 $w=3.7e-07 $l=1.56e-06 $layer=MET1_cond $X=7.865 $Y=0.44
+ $X2=9.425 $Y2=0.44
r120 88 91 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=7.685 $Y=0.51
+ $X2=7.685 $Y2=0.68
r121 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.865 $Y=0.51
+ $X2=7.865 $Y2=0.51
r122 86 108 1.0711 $w=3.7e-07 $l=2.79e-06 $layer=MET1_cond $X=6.895 $Y=7.7
+ $X2=9.685 $Y2=7.7
r123 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.895 $Y=7.63
+ $X2=6.895 $Y2=7.63
r124 83 85 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=6.715 $Y=7.46
+ $X2=6.715 $Y2=7.63
r125 80 83 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=6.715 $Y=6.25
+ $X2=6.715 $Y2=7.46
r126 75 77 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=6.125 $Y=0.68
+ $X2=6.125 $Y2=1.89
r127 73 89 0.598892 $w=3.7e-07 $l=1.56e-06 $layer=MET1_cond $X=6.305 $Y=0.44
+ $X2=7.865 $Y2=0.44
r128 72 75 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=6.125 $Y=0.51
+ $X2=6.125 $Y2=0.68
r129 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.305 $Y=0.51
+ $X2=6.305 $Y2=0.51
r130 67 69 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=5.155 $Y=7.46
+ $X2=5.155 $Y2=7.63
r131 64 67 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=5.155 $Y=6.25
+ $X2=5.155 $Y2=7.46
r132 59 113 0.224585 $w=3.7e-07 $l=5.85e-07 $layer=MET1_cond $X=4.215 $Y=0.44
+ $X2=4.8 $Y2=0.44
r133 58 61 6.89266 $w=5.88e-07 $l=3.4e-07 $layer=LI1_cond $X=4.035 $Y=0.51
+ $X2=4.035 $Y2=0.85
r134 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.215 $Y=0.51
+ $X2=4.215 $Y2=0.51
r135 56 122 0.355112 $w=3.7e-07 $l=9.25e-07 $layer=MET1_cond $X=3.775 $Y=7.7
+ $X2=4.7 $Y2=7.7
r136 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.775 $Y=7.63
+ $X2=3.775 $Y2=7.63
r137 53 55 3.44633 $w=5.88e-07 $l=1.7e-07 $layer=LI1_cond $X=3.595 $Y=7.46
+ $X2=3.595 $Y2=7.63
r138 50 53 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=3.595 $Y=6.25
+ $X2=3.595 $Y2=7.46
r139 46 86 0.620007 $w=3.7e-07 $l=1.615e-06 $layer=MET1_cond $X=5.28 $Y=7.7
+ $X2=6.895 $Y2=7.7
r140 46 122 0.222665 $w=3.7e-07 $l=5.8e-07 $layer=MET1_cond $X=5.28 $Y=7.7
+ $X2=4.7 $Y2=7.7
r141 46 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.335 $Y=7.63
+ $X2=5.335 $Y2=7.63
r142 45 73 0.393503 $w=3.7e-07 $l=1.025e-06 $layer=MET1_cond $X=5.28 $Y=0.44
+ $X2=6.305 $Y2=0.44
r143 45 113 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=5.28 $Y=0.44
+ $X2=4.8 $Y2=0.44
r144 44 96 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=9.245 $Y=0.425
+ $X2=9.245 $Y2=0.51
r145 42 88 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=7.685 $Y=0.425
+ $X2=7.685 $Y2=0.51
r146 42 43 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.685 $Y=0.425
+ $X2=7.685 $Y2=0.34
r147 41 85 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=6.715 $Y=7.715
+ $X2=6.715 $Y2=7.63
r148 39 72 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=6.125 $Y=0.425
+ $X2=6.125 $Y2=0.51
r149 39 40 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.125 $Y=0.425
+ $X2=6.125 $Y2=0.34
r150 37 69 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=7.715
+ $X2=5.155 $Y2=7.63
r151 37 38 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=7.715
+ $X2=5.155 $Y2=7.8
r152 36 58 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=0.425
+ $X2=4.035 $Y2=0.51
r153 35 55 1.72316 $w=5.88e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=7.715
+ $X2=3.595 $Y2=7.63
r154 34 43 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=7.98 $Y=0.34
+ $X2=7.685 $Y2=0.34
r155 33 44 9.96617 $w=1.7e-07 $l=3.34813e-07 $layer=LI1_cond $X=8.95 $Y=0.34
+ $X2=9.245 $Y2=0.425
r156 33 34 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=8.95 $Y=0.34
+ $X2=7.98 $Y2=0.34
r157 32 40 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.42 $Y=0.34
+ $X2=6.125 $Y2=0.34
r158 31 43 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=7.39 $Y=0.34
+ $X2=7.685 $Y2=0.34
r159 31 32 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=7.39 $Y=0.34
+ $X2=6.42 $Y2=0.34
r160 30 38 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=5.45 $Y=7.8
+ $X2=5.155 $Y2=7.8
r161 29 41 9.96617 $w=1.7e-07 $l=3.34813e-07 $layer=LI1_cond $X=6.42 $Y=7.8
+ $X2=6.715 $Y2=7.715
r162 29 30 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=6.42 $Y=7.8
+ $X2=5.45 $Y2=7.8
r163 28 36 9.96617 $w=1.7e-07 $l=3.34813e-07 $layer=LI1_cond $X=4.33 $Y=0.34
+ $X2=4.035 $Y2=0.425
r164 27 40 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=5.83 $Y=0.34
+ $X2=6.125 $Y2=0.34
r165 27 28 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=5.83 $Y=0.34
+ $X2=4.33 $Y2=0.34
r166 26 35 9.96617 $w=1.7e-07 $l=3.34813e-07 $layer=LI1_cond $X=3.89 $Y=7.8
+ $X2=3.595 $Y2=7.715
r167 25 38 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=4.86 $Y=7.8
+ $X2=5.155 $Y2=7.8
r168 25 26 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=4.86 $Y=7.8
+ $X2=3.89 $Y2=7.8
r169 8 104 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=9.38
+ $Y=6.855 $X2=9.505 $Y2=7
r170 7 101 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=9.105
+ $Y=0.535 $X2=9.245 $Y2=1.89
r171 7 99 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.105
+ $Y=0.535 $X2=9.245 $Y2=0.68
r172 6 93 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=7.545
+ $Y=0.535 $X2=7.685 $Y2=1.89
r173 6 91 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.545
+ $Y=0.535 $X2=7.685 $Y2=0.68
r174 5 83 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=6.575
+ $Y=6.105 $X2=6.715 $Y2=7.46
r175 5 80 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.575
+ $Y=6.105 $X2=6.715 $Y2=6.25
r176 4 77 91 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_NDIFF $count=2 $X=6
+ $Y=0.535 $X2=6.125 $Y2=1.89
r177 4 75 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6
+ $Y=0.535 $X2=6.125 $Y2=0.68
r178 3 67 91 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_NDIFF $count=2 $X=5.015
+ $Y=6.105 $X2=5.155 $Y2=7.46
r179 3 64 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.015
+ $Y=6.105 $X2=5.155 $Y2=6.25
r180 2 61 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.895
+ $Y=0.705 $X2=4.035 $Y2=0.85
r181 1 53 91 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_NDIFF $count=2 $X=3.47
+ $Y=6.105 $X2=3.595 $Y2=7.46
r182 1 50 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=3.47
+ $Y=6.105 $X2=3.595 $Y2=6.25
.ends

