* NGSPICE file created from sky130_fd_sc_hvl__nor3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__nor3_1 A B C VGND VNB VPB VPWR Y
M1000 a_205_443# A VPWR VPB phv w=1.5e+06u l=500000u
+  ad=3.15e+11p pd=3.42e+06u as=4.275e+11p ps=3.57e+06u
M1001 a_347_443# B a_205_443# VPB phv w=1.5e+06u l=500000u
+  ad=3.15e+11p pd=3.42e+06u as=0p ps=0u
M1002 Y C a_347_443# VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=0p ps=0u
M1003 Y A VGND VNB nhv w=750000u l=500000u
+  ad=4.0875e+11p pd=4.09e+06u as=4.0875e+11p ps=4.09e+06u
M1004 Y C VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B Y VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends

