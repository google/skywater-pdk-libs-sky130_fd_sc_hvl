# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__sdlxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdlxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.040000 2.185000 2.370000 3.260000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.060000 0.515000 11.400000 3.755000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515000 1.525000 3.860000 2.495000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  1.005000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 1.835000 2.770000 2.005000 ;
        RECT 0.585000 2.005000 1.795000 2.775000 ;
        RECT 2.600000 1.445000 2.985000 1.695000 ;
        RECT 2.600000 1.695000 2.770000 1.835000 ;
    END
  END SCE
  PIN GATE
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.370000 1.145000 4.665000 2.495000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 11.520000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 11.520000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 11.520000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 11.520000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 11.850000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 11.520000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.520000 0.085000 ;
      RECT  0.000000  3.985000 11.520000 4.155000 ;
      RECT  0.130000  0.495000  0.480000 1.175000 ;
      RECT  0.130000  1.175000  3.335000 1.265000 ;
      RECT  0.130000  1.265000  2.295000 1.345000 ;
      RECT  0.130000  1.345000  0.380000 3.395000 ;
      RECT  0.560000  2.995000  1.510000 3.705000 ;
      RECT  0.660000  0.365000  1.610000 0.995000 ;
      RECT  1.965000  1.095000  3.335000 1.175000 ;
      RECT  1.965000  1.345000  2.295000 1.655000 ;
      RECT  2.420000  0.495000  2.750000 0.745000 ;
      RECT  2.420000  0.745000  3.685000 0.915000 ;
      RECT  2.575000  2.675000  4.665000 2.845000 ;
      RECT  2.575000  2.845000  2.825000 3.725000 ;
      RECT  2.950000  1.905000  3.335000 2.495000 ;
      RECT  3.165000  1.265000  3.335000 1.905000 ;
      RECT  3.365000  3.025000  4.315000 3.725000 ;
      RECT  3.515000  0.915000  3.685000 1.175000 ;
      RECT  3.515000  1.175000  4.200000 1.345000 ;
      RECT  3.865000  0.365000  4.455000 0.975000 ;
      RECT  4.030000  1.345000  4.200000 2.675000 ;
      RECT  4.495000  2.845000  4.665000 3.635000 ;
      RECT  4.495000  3.635000  5.365000 3.805000 ;
      RECT  4.695000  0.515000  5.025000 0.975000 ;
      RECT  4.845000  0.975000  5.015000 1.175000 ;
      RECT  4.845000  1.175000  5.920000 1.345000 ;
      RECT  4.845000  1.345000  5.015000 3.455000 ;
      RECT  5.195000  2.235000  6.065000 2.405000 ;
      RECT  5.195000  2.405000  5.365000 3.635000 ;
      RECT  5.205000  0.365000  5.795000 0.995000 ;
      RECT  5.545000  2.585000  5.715000 3.705000 ;
      RECT  5.590000  1.345000  5.920000 1.845000 ;
      RECT  5.895000  2.405000  6.065000 3.595000 ;
      RECT  5.895000  3.595000  7.250000 3.765000 ;
      RECT  6.045000  0.265000  7.275000 0.435000 ;
      RECT  6.045000  0.435000  6.415000 0.975000 ;
      RECT  6.245000  0.975000  6.415000 2.585000 ;
      RECT  6.245000  2.585000  6.575000 3.415000 ;
      RECT  6.595000  0.615000  6.925000 0.975000 ;
      RECT  6.755000  0.975000  6.925000 2.925000 ;
      RECT  6.755000  2.925000  7.250000 3.595000 ;
      RECT  7.105000  0.435000  7.275000 1.585000 ;
      RECT  7.105000  1.585000  8.010000 1.755000 ;
      RECT  7.455000  0.495000  7.705000 1.075000 ;
      RECT  7.455000  1.075000  8.360000 1.245000 ;
      RECT  7.700000  2.925000  8.030000 3.755000 ;
      RECT  7.840000  1.755000  8.010000 2.215000 ;
      RECT  7.840000  2.215000  8.570000 2.475000 ;
      RECT  7.860000  2.655000  8.920000 2.825000 ;
      RECT  7.860000  2.825000  8.030000 2.925000 ;
      RECT  8.190000  1.245000  8.360000 1.835000 ;
      RECT  8.190000  1.835000 10.200000 2.005000 ;
      RECT  8.245000  0.365000  9.195000 0.895000 ;
      RECT  8.540000  1.075000  8.870000 1.405000 ;
      RECT  8.540000  1.405000 10.550000 1.575000 ;
      RECT  8.540000  1.575000  8.870000 1.655000 ;
      RECT  8.685000  3.005000  9.635000 3.705000 ;
      RECT  8.750000  2.005000  8.920000 2.655000 ;
      RECT  9.385000  2.185000 10.550000 2.355000 ;
      RECT  9.385000  2.355000  9.715000 2.675000 ;
      RECT  9.415000  0.845000  9.745000 1.405000 ;
      RECT  9.870000  1.755000 10.200000 1.835000 ;
      RECT  9.895000  2.535000 10.845000 3.755000 ;
      RECT  9.925000  0.365000 10.875000 1.225000 ;
      RECT 10.380000  1.575000 10.550000 2.185000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.590000  3.505000  0.760000 3.675000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.690000  0.395000  0.860000 0.565000 ;
      RECT  0.950000  3.505000  1.120000 3.675000 ;
      RECT  1.050000  0.395000  1.220000 0.565000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.310000  3.505000  1.480000 3.675000 ;
      RECT  1.410000  0.395000  1.580000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.395000  3.505000  3.565000 3.675000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.755000  3.505000  3.925000 3.675000 ;
      RECT  3.895000  0.395000  4.065000 0.565000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.115000  3.505000  4.285000 3.675000 ;
      RECT  4.255000  0.395000  4.425000 0.565000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.235000  0.395000  5.405000 0.565000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.545000  3.505000  5.715000 3.675000 ;
      RECT  5.595000  0.395000  5.765000 0.565000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.275000  0.395000  8.445000 0.565000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.635000  0.395000  8.805000 0.565000 ;
      RECT  8.715000  3.505000  8.885000 3.675000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.995000  0.395000  9.165000 0.565000 ;
      RECT  9.075000  3.505000  9.245000 3.675000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.435000  3.505000  9.605000 3.675000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.925000  3.505000 10.095000 3.675000 ;
      RECT  9.955000  0.395000 10.125000 0.565000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.285000  3.505000 10.455000 3.675000 ;
      RECT 10.315000  0.395000 10.485000 0.565000 ;
      RECT 10.645000  3.505000 10.815000 3.675000 ;
      RECT 10.675000  0.395000 10.845000 0.565000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
  END
END sky130_fd_sc_hvl__sdlxtp_1
END LIBRARY
