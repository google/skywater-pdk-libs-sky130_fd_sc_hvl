* NGSPICE file created from sky130_fd_sc_hvl__and2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__and2_1 A B VGND VNB VPB VPWR X
M1000 X a_30_107# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=7.509e+11p ps=5.41e+06u
M1001 a_30_107# A VPWR VPB phv w=420000u l=500000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1002 X a_30_107# VGND VNB nhv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=4.3845e+11p ps=3.14e+06u
M1003 VPWR B a_30_107# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND B a_183_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1005 a_183_107# A a_30_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends

