* File: sky130_fd_sc_hvl__and2_1.pex.spice
* Created: Wed Sep  2 09:03:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__AND2_1%VNB 5 7 11 25
r23 7 25 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0.058
r24 7 11 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0
r25 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r26 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__AND2_1%VPB 4 6 14 21
r23 10 21 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=4.07
+ $X2=1.68 $Y2=4.013
r24 10 14 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=4.07
+ $X2=3.12 $Y2=4.07
r25 9 14 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=3.12 $Y2=4.07
r26 9 10 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r27 6 21 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=4.012
+ $X2=1.68 $Y2=4.013
r28 4 14 52 $w=1.7e-07 $l=3.16221e-06 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=3.12 $Y2=4.07
r29 4 9 52 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__AND2_1%A 5 9 10 11 12 13 17
r34 17 19 23.0439 $w=7.15e-07 $l=2.55e-07 $layer=POLY_cond $X=0.557 $Y=1.34
+ $X2=0.557 $Y2=1.085
r35 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.34 $X2=0.385 $Y2=1.34
r36 13 18 9.13522 $w=4.08e-07 $l=3.25e-07 $layer=LI1_cond $X=0.33 $Y=1.665
+ $X2=0.33 $Y2=1.34
r37 12 18 1.26488 $w=4.08e-07 $l=4.5e-08 $layer=LI1_cond $X=0.33 $Y=1.295
+ $X2=0.33 $Y2=1.34
r38 10 11 15.8527 $w=7.15e-07 $l=1.55e-07 $layer=POLY_cond $X=0.672 $Y=1.95
+ $X2=0.672 $Y2=2.105
r39 9 11 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.895 $Y=2.425 $X2=0.895
+ $Y2=2.105
r40 5 19 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.665 $Y=0.745 $X2=0.665
+ $Y2=1.085
r41 1 17 7.33504 $w=7.15e-07 $l=1.02e-07 $layer=POLY_cond $X=0.557 $Y=1.442
+ $X2=0.557 $Y2=1.34
r42 1 10 36.5314 $w=7.15e-07 $l=5.08e-07 $layer=POLY_cond $X=0.557 $Y=1.442
+ $X2=0.557 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HVL__AND2_1%B 1 3 6 8 9 17
c38 17 0 1.08281e-19 $X=1.675 $Y=1.402
c39 6 0 9.31747e-20 $X=1.675 $Y=2.425
c40 1 0 1.77546e-19 $X=1.375 $Y=1.065
r41 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.29
+ $Y=1.23 $X2=1.29 $Y2=1.23
r42 9 14 1.92074 $w=3.88e-07 $l=6.5e-08 $layer=LI1_cond $X=1.26 $Y=1.295
+ $X2=1.26 $Y2=1.23
r43 8 14 9.0127 $w=3.88e-07 $l=3.05e-07 $layer=LI1_cond $X=1.26 $Y=0.925
+ $X2=1.26 $Y2=1.23
r44 4 17 9.86319 $w=5e-07 $l=3.38e-07 $layer=POLY_cond $X=1.675 $Y=1.74
+ $X2=1.675 $Y2=1.402
r45 4 6 73.299 $w=5e-07 $l=6.85e-07 $layer=POLY_cond $X=1.675 $Y=1.74 $X2=1.675
+ $Y2=2.425
r46 1 17 23.7791 $w=6.75e-07 $l=3e-07 $layer=POLY_cond $X=1.375 $Y=1.402
+ $X2=1.675 $Y2=1.402
r47 1 13 6.73741 $w=6.75e-07 $l=8.5e-08 $layer=POLY_cond $X=1.375 $Y=1.402
+ $X2=1.29 $Y2=1.402
r48 1 3 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.375 $Y=1.065 $X2=1.375
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__AND2_1%A_30_107# 1 2 9 13 17 19 20 22 23 24 27 29
+ 31 33 34
c65 33 0 9.31747e-20 $X=2.61 $Y=1.89
c66 22 0 1.08281e-19 $X=0.8 $Y=1.905
c67 19 0 1.77546e-19 $X=0.715 $Y=0.91
r68 34 40 20.0636 $w=5.2e-07 $l=1.95e-07 $layer=POLY_cond $X=2.685 $Y=1.89
+ $X2=2.685 $Y2=2.085
r69 34 39 48.8729 $w=5.2e-07 $l=4.75e-07 $layer=POLY_cond $X=2.685 $Y=1.89
+ $X2=2.685 $Y2=1.415
r70 33 36 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.61 $Y=1.89 $X2=2.61
+ $Y2=1.99
r71 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.89 $X2=2.61 $Y2=1.89
r72 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=1.99
+ $X2=1.285 $Y2=1.99
r73 29 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=1.99
+ $X2=2.61 $Y2=1.99
r74 29 30 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=2.445 $Y=1.99
+ $X2=1.37 $Y2=1.99
r75 25 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.075
+ $X2=1.285 $Y2=1.99
r76 25 27 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.285 $Y=2.075
+ $X2=1.285 $Y2=2.425
r77 23 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.99 $X2=1.285
+ $Y2=1.99
r78 23 24 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.2 $Y=1.99
+ $X2=0.885 $Y2=1.99
r79 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.8 $Y=1.905
+ $X2=0.885 $Y2=1.99
r80 21 22 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.8 $Y=0.995 $X2=0.8
+ $Y2=1.905
r81 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.715 $Y=0.91
+ $X2=0.8 $Y2=0.995
r82 19 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.715 $Y=0.91
+ $X2=0.38 $Y2=0.91
r83 15 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.255 $Y=0.825
+ $X2=0.38 $Y2=0.91
r84 15 17 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=0.255 $Y=0.825
+ $X2=0.255 $Y2=0.745
r85 13 39 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.695 $Y=0.91
+ $X2=2.695 $Y2=1.415
r86 9 40 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.675 $Y=2.965
+ $X2=2.675 $Y2=2.085
r87 2 27 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=2.215 $X2=1.285 $Y2=2.425
r88 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.535 $X2=0.275 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__AND2_1%VPWR 1 2 7 10 19 28
r25 24 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.715 $Y=3.59
+ $X2=2.715 $Y2=3.59
r26 22 24 8.1496 $w=1.248e-06 $l=8.35e-07 $layer=LI1_cond $X=2.175 $Y=2.755
+ $X2=2.175 $Y2=3.59
r27 19 22 4.0504 $w=1.248e-06 $l=4.15e-07 $layer=LI1_cond $X=2.175 $Y=2.34
+ $X2=2.175 $Y2=2.755
r28 14 16 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.195 $Y=3.63
+ $X2=0.915 $Y2=3.63
r29 13 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.915 $Y=3.59
+ $X2=0.915 $Y2=3.59
r30 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.195 $Y=3.59
+ $X2=0.195 $Y2=3.59
r31 10 13 15.2828 $w=9.28e-07 $l=1.165e-06 $layer=LI1_cond $X=0.555 $Y=2.425
+ $X2=0.555 $Y2=3.59
r32 7 28 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=1.635 $Y=3.63
+ $X2=2.715 $Y2=3.63
r33 7 16 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.635 $Y=3.63
+ $X2=0.915 $Y2=3.63
r34 7 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.635 $Y=3.59
+ $X2=1.635 $Y2=3.59
r35 2 24 400 $w=1.7e-07 $l=1.49708e-06 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=2.215 $X2=2.18 $Y2=3.59
r36 2 22 400 $w=1.7e-07 $l=6.5521e-07 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=2.215 $X2=2.18 $Y2=2.755
r37 2 19 600 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=2.215 $X2=2.18 $Y2=2.34
r38 1 10 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.36
+ $Y=2.215 $X2=0.505 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_HVL__AND2_1%X 1 2 7 8 9 10 11 12 13 22
r14 13 40 18.6486 $w=2.73e-07 $l=4.45e-07 $layer=LI1_cond $X=3.117 $Y=3.145
+ $X2=3.117 $Y2=3.59
r15 12 13 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.117 $Y=2.775
+ $X2=3.117 $Y2=3.145
r16 11 12 18.2296 $w=2.73e-07 $l=4.35e-07 $layer=LI1_cond $X=3.117 $Y=2.34
+ $X2=3.117 $Y2=2.775
r17 10 11 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=3.117 $Y=2.035
+ $X2=3.117 $Y2=2.34
r18 9 10 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.117 $Y=1.665
+ $X2=3.117 $Y2=2.035
r19 8 9 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.117 $Y=1.295
+ $X2=3.117 $Y2=1.665
r20 7 8 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.117 $Y=0.925
+ $X2=3.117 $Y2=1.295
r21 7 22 10.2672 $w=2.73e-07 $l=2.45e-07 $layer=LI1_cond $X=3.117 $Y=0.925
+ $X2=3.117 $Y2=0.68
r22 2 40 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.925
+ $Y=2.215 $X2=3.065 $Y2=3.59
r23 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.925
+ $Y=2.215 $X2=3.065 $Y2=2.34
r24 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.535 $X2=3.085 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__AND2_1%VGND 1 4 7 11
r24 15 17 5.11414 $w=9.88e-07 $l=4.15e-07 $layer=LI1_cond $X=2.13 $Y=0.745
+ $X2=2.13 $Y2=1.16
r25 13 15 1.04747 $w=9.88e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=0.66
+ $X2=2.13 $Y2=0.745
r26 8 11 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.77 $Y=0.44
+ $X2=2.49 $Y2=0.44
r27 7 13 2.21818 $w=9.88e-07 $l=1.8e-07 $layer=LI1_cond $X=2.13 $Y=0.48 $X2=2.13
+ $Y2=0.66
r28 7 11 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.49 $Y=0.48
+ $X2=2.49 $Y2=0.48
r29 7 8 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.77 $Y=0.48 $X2=1.77
+ $Y2=0.48
r30 4 8 0.0345515 $w=3.7e-07 $l=9e-08 $layer=MET1_cond $X=1.68 $Y=0.44 $X2=1.77
+ $Y2=0.44
r31 1 17 182 $w=1.7e-07 $l=9.42019e-07 $layer=licon1_NDIFF $count=1 $X=1.625
+ $Y=0.535 $X2=2.305 $Y2=1.16
r32 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.625
+ $Y=0.535 $X2=1.765 $Y2=0.745
r33 1 13 182 $w=1.7e-07 $l=7.39865e-07 $layer=licon1_NDIFF $count=1 $X=1.625
+ $Y=0.535 $X2=2.305 $Y2=0.66
.ends

