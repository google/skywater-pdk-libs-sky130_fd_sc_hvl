# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hvl__dfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.545000 3.350000 2.125000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.455000 0.675000 10.890000 1.465000 ;
        RECT 10.455000 2.195000 10.890000 3.735000 ;
        RECT 10.685000 1.465000 10.890000 2.195000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.460000 2.175000 13.810000 3.755000 ;
        RECT 13.480000 0.675000 13.810000 2.175000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.550000 0.890000 2.220000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 13.920000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 13.920000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 13.920000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 13.920000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.985000 13.920000 4.155000 ;
      RECT  0.110000  0.540000  0.440000 1.200000 ;
      RECT  0.110000  1.200000  1.545000 1.370000 ;
      RECT  0.110000  1.370000  0.380000 3.230000 ;
      RECT  0.570000  2.400000  1.160000 3.705000 ;
      RECT  0.620000  0.365000  1.570000 1.020000 ;
      RECT  1.215000  1.370000  1.545000 1.870000 ;
      RECT  1.340000  1.870000  1.510000 3.410000 ;
      RECT  1.340000  3.410000  2.290000 3.580000 ;
      RECT  1.690000  2.400000  1.940000 3.230000 ;
      RECT  1.750000  0.520000  1.920000 1.195000 ;
      RECT  1.750000  1.195000  3.340000 1.365000 ;
      RECT  1.750000  1.365000  1.940000 2.400000 ;
      RECT  2.100000  0.365000  2.990000 1.015000 ;
      RECT  2.120000  2.305000  3.350000 2.475000 ;
      RECT  2.120000  2.475000  2.290000 3.410000 ;
      RECT  2.470000  2.655000  3.000000 3.705000 ;
      RECT  3.170000  0.265000  4.980000 0.435000 ;
      RECT  3.170000  0.435000  3.340000 1.195000 ;
      RECT  3.180000  2.475000  3.350000 3.335000 ;
      RECT  3.180000  3.335000  5.085000 3.505000 ;
      RECT  3.520000  0.615000  3.850000 0.935000 ;
      RECT  3.530000  0.935000  3.700000 2.655000 ;
      RECT  3.530000  2.655000  3.770000 3.155000 ;
      RECT  3.880000  1.115000  4.120000 1.785000 ;
      RECT  3.950000  1.785000  4.120000 3.335000 ;
      RECT  4.300000  0.615000  4.630000 1.015000 ;
      RECT  4.300000  1.015000  4.470000 1.905000 ;
      RECT  4.300000  1.905000  6.540000 2.075000 ;
      RECT  4.300000  2.075000  4.550000 3.155000 ;
      RECT  4.650000  1.195000  4.980000 1.245000 ;
      RECT  4.650000  1.245000  6.485000 1.415000 ;
      RECT  4.650000  1.415000  4.980000 1.725000 ;
      RECT  4.755000  2.255000  5.085000 2.635000 ;
      RECT  4.755000  2.635000  6.565000 2.805000 ;
      RECT  4.755000  2.805000  5.085000 3.335000 ;
      RECT  4.810000  0.435000  4.980000 1.195000 ;
      RECT  5.185000  0.365000  6.135000 1.065000 ;
      RECT  5.265000  2.985000  6.215000 3.715000 ;
      RECT  5.435000  2.255000  5.765000 2.285000 ;
      RECT  5.435000  2.285000  6.915000 2.455000 ;
      RECT  6.210000  1.595000  6.540000 1.905000 ;
      RECT  6.210000  2.075000  6.540000 2.105000 ;
      RECT  6.315000  0.265000  7.345000 0.435000 ;
      RECT  6.315000  0.435000  6.485000 1.245000 ;
      RECT  6.395000  2.805000  6.565000 3.635000 ;
      RECT  6.395000  3.635000  8.245000 3.805000 ;
      RECT  6.665000  0.615000  6.995000 1.325000 ;
      RECT  6.745000  1.325000  6.915000 2.285000 ;
      RECT  6.745000  2.455000  6.915000 3.455000 ;
      RECT  7.095000  2.205000  7.425000 2.495000 ;
      RECT  7.095000  2.495000  7.265000 3.635000 ;
      RECT  7.175000  0.435000  7.345000 1.195000 ;
      RECT  7.175000  1.195000  7.445000 1.865000 ;
      RECT  7.445000  2.675000  7.795000 3.455000 ;
      RECT  7.540000  0.515000  8.595000 0.685000 ;
      RECT  7.540000  0.685000  7.795000 1.015000 ;
      RECT  7.625000  1.015000  7.795000 2.675000 ;
      RECT  7.975000  1.105000  8.245000 3.635000 ;
      RECT  8.425000  0.685000  8.595000 2.325000 ;
      RECT  8.425000  2.325000  9.725000 2.495000 ;
      RECT  8.505000  2.675000  9.455000 3.715000 ;
      RECT  8.775000  0.365000  9.725000 1.325000 ;
      RECT  8.775000  1.505000 10.235000 1.645000 ;
      RECT  8.775000  1.645000 10.505000 1.675000 ;
      RECT  8.775000  1.675000  9.105000 2.145000 ;
      RECT  9.395000  1.855000  9.725000 2.325000 ;
      RECT  9.905000  0.535000 10.235000 1.505000 ;
      RECT  9.905000  1.675000 10.505000 1.975000 ;
      RECT  9.905000  1.975000 10.235000 3.715000 ;
      RECT 11.070000  0.365000 11.625000 1.485000 ;
      RECT 11.070000  2.195000 11.605000 3.735000 ;
      RECT 11.785000  2.195000 12.115000 2.985000 ;
      RECT 11.805000  1.005000 12.135000 1.665000 ;
      RECT 11.805000  1.665000 13.300000 1.995000 ;
      RECT 11.805000  1.995000 12.115000 2.195000 ;
      RECT 12.295000  2.175000 13.245000 3.755000 ;
      RECT 12.315000  0.365000 13.265000 1.485000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.600000  3.505000  0.770000 3.675000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.650000  0.395000  0.820000 0.565000 ;
      RECT  0.960000  3.505000  1.130000 3.675000 ;
      RECT  1.010000  0.395000  1.180000 0.565000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.370000  0.395000  1.540000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.100000  0.395000  2.270000 0.565000 ;
      RECT  2.460000  0.395000  2.630000 0.565000 ;
      RECT  2.470000  3.505000  2.640000 3.675000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.820000  0.395000  2.990000 0.565000 ;
      RECT  2.830000  3.505000  3.000000 3.675000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.215000  0.395000  5.385000 0.565000 ;
      RECT  5.295000  3.505000  5.465000 3.675000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.575000  0.395000  5.745000 0.565000 ;
      RECT  5.655000  3.505000  5.825000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  5.935000  0.395000  6.105000 0.565000 ;
      RECT  6.015000  3.505000  6.185000 3.675000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.535000  3.515000  8.705000 3.685000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.805000  0.395000  8.975000 0.565000 ;
      RECT  8.895000  3.515000  9.065000 3.685000 ;
      RECT  9.165000  0.395000  9.335000 0.565000 ;
      RECT  9.255000  3.515000  9.425000 3.685000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.525000  0.395000  9.695000 0.565000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 11.070000  3.505000 11.240000 3.675000 ;
      RECT 11.080000  0.395000 11.250000 0.565000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.430000  3.505000 11.600000 3.675000 ;
      RECT 11.440000  0.395000 11.610000 0.565000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.325000  3.505000 12.495000 3.675000 ;
      RECT 12.345000  0.395000 12.515000 0.565000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 12.685000  3.505000 12.855000 3.675000 ;
      RECT 12.705000  0.395000 12.875000 0.565000 ;
      RECT 13.045000  3.505000 13.215000 3.675000 ;
      RECT 13.065000  0.395000 13.235000 0.565000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
  END
END sky130_fd_sc_hvl__dfxbp_1
