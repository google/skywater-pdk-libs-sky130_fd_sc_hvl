* File: sky130_fd_sc_hvl__nand3_1.pxi.spice
* Created: Wed Sep  2 09:08:31 2020
* 
x_PM_SKY130_FD_SC_HVL__NAND3_1%VNB N_VNB_M1002_b VNB N_VNB_c_7_p VNB
+ PM_SKY130_FD_SC_HVL__NAND3_1%VNB
x_PM_SKY130_FD_SC_HVL__NAND3_1%VPB N_VPB_M1001_b VPB N_VPB_c_20_p VPB
+ PM_SKY130_FD_SC_HVL__NAND3_1%VPB
x_PM_SKY130_FD_SC_HVL__NAND3_1%C N_C_M1001_g N_C_M1002_g C C N_C_c_49_n
+ N_C_c_50_n PM_SKY130_FD_SC_HVL__NAND3_1%C
x_PM_SKY130_FD_SC_HVL__NAND3_1%B N_B_M1003_g N_B_M1004_g B B N_B_c_70_n
+ N_B_c_71_n PM_SKY130_FD_SC_HVL__NAND3_1%B
x_PM_SKY130_FD_SC_HVL__NAND3_1%A N_A_M1005_g N_A_M1000_g A A N_A_c_100_n
+ N_A_c_101_n PM_SKY130_FD_SC_HVL__NAND3_1%A
x_PM_SKY130_FD_SC_HVL__NAND3_1%VPWR N_VPWR_M1001_s N_VPWR_M1004_d VPWR
+ N_VPWR_c_128_n N_VPWR_c_131_n N_VPWR_c_134_n PM_SKY130_FD_SC_HVL__NAND3_1%VPWR
x_PM_SKY130_FD_SC_HVL__NAND3_1%Y N_Y_M1005_d N_Y_M1001_d N_Y_M1000_d N_Y_c_155_n
+ N_Y_c_158_n N_Y_c_159_n Y Y Y Y Y Y Y N_Y_c_153_n Y
+ PM_SKY130_FD_SC_HVL__NAND3_1%Y
x_PM_SKY130_FD_SC_HVL__NAND3_1%VGND N_VGND_M1002_s VGND N_VGND_c_194_n
+ PM_SKY130_FD_SC_HVL__NAND3_1%VGND
cc_1 N_VNB_M1002_b N_C_M1002_g 0.043166f $X=-0.33 $Y=-0.265 $X2=0.965 $Y2=0.91
cc_2 N_VNB_M1002_b N_C_c_49_n 0.0552106f $X=-0.33 $Y=-0.265 $X2=0.83 $Y2=1.67
cc_3 N_VNB_M1002_b N_C_c_50_n 0.0287494f $X=-0.33 $Y=-0.265 $X2=0.83 $Y2=1.67
cc_4 N_VNB_M1002_b B 0.00396701f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_5 N_VNB_M1002_b N_B_c_70_n 0.0573719f $X=-0.33 $Y=-0.265 $X2=0.93 $Y2=1.67
cc_6 N_VNB_M1002_b N_B_c_71_n 0.0418452f $X=-0.33 $Y=-0.265 $X2=0.83 $Y2=1.67
cc_7 N_VNB_c_7_p N_B_c_71_n 0.00102867f $X=0.24 $Y=0 $X2=0.83 $Y2=1.67
cc_8 N_VNB_M1002_b N_A_c_100_n 0.0542405f $X=-0.33 $Y=-0.265 $X2=0.93 $Y2=1.67
cc_9 N_VNB_M1002_b N_A_c_101_n 0.0533149f $X=-0.33 $Y=-0.265 $X2=0.83 $Y2=1.67
cc_10 N_VNB_c_7_p N_A_c_101_n 0.0023273f $X=0.24 $Y=0 $X2=0.83 $Y2=1.67
cc_11 N_VNB_M1002_b Y 0.0371209f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_12 N_VNB_M1002_b N_Y_c_153_n 0.0363671f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_13 N_VNB_c_7_p N_Y_c_153_n 7.68678e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_14 N_VNB_M1002_b VGND 0.0707978f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_15 N_VNB_c_7_p VGND 0.359386f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_16 N_VNB_M1002_b N_VGND_c_194_n 0.133639f $X=-0.33 $Y=-0.265 $X2=0.965
+ $Y2=0.91
cc_17 N_VNB_c_7_p N_VGND_c_194_n 0.00457781f $X=0.24 $Y=0 $X2=0.965 $Y2=0.91
cc_18 N_VPB_M1001_b N_C_M1001_g 0.041634f $X=-0.33 $Y=1.885 $X2=0.895 $Y2=2.965
cc_19 VPB N_C_M1001_g 0.00970178f $X=0 $Y=3.955 $X2=0.895 $Y2=2.965
cc_20 N_VPB_c_20_p N_C_M1001_g 0.0152133f $X=3.12 $Y=4.07 $X2=0.895 $Y2=2.965
cc_21 N_VPB_M1001_b N_C_c_49_n 0.0285452f $X=-0.33 $Y=1.885 $X2=0.83 $Y2=1.67
cc_22 N_VPB_M1001_b N_B_M1004_g 0.0536223f $X=-0.33 $Y=1.885 $X2=0.965 $Y2=0.91
cc_23 VPB N_B_M1004_g 0.00970178f $X=0 $Y=3.955 $X2=0.965 $Y2=0.91
cc_24 N_VPB_c_20_p N_B_M1004_g 0.0152133f $X=3.12 $Y=4.07 $X2=0.965 $Y2=0.91
cc_25 N_VPB_M1001_b N_B_c_70_n 0.00611819f $X=-0.33 $Y=1.885 $X2=0.93 $Y2=1.67
cc_26 N_VPB_M1001_b N_A_M1000_g 0.060447f $X=-0.33 $Y=1.885 $X2=0.965 $Y2=0.91
cc_27 VPB N_A_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.965 $Y2=0.91
cc_28 N_VPB_c_20_p N_A_M1000_g 0.0152133f $X=3.12 $Y=4.07 $X2=0.965 $Y2=0.91
cc_29 N_VPB_M1001_b N_A_c_100_n 0.00301588f $X=-0.33 $Y=1.885 $X2=0.93 $Y2=1.67
cc_30 N_VPB_M1001_b N_VPWR_c_128_n 0.0820659f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_31 VPB N_VPWR_c_128_n 0.00349285f $X=0 $Y=3.955 $X2=0.635 $Y2=1.58
cc_32 N_VPB_c_20_p N_VPWR_c_128_n 0.0475576f $X=3.12 $Y=4.07 $X2=0.635 $Y2=1.58
cc_33 N_VPB_M1001_b N_VPWR_c_131_n 0.00243985f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_131_n 0.00512219f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_35 N_VPB_c_20_p N_VPWR_c_131_n 0.0629871f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_36 N_VPB_M1001_b N_VPWR_c_134_n 0.0451682f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_134_n 0.35668f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_38 N_VPB_c_20_p N_VPWR_c_134_n 0.0146238f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_39 N_VPB_M1001_b N_Y_c_155_n 0.00357947f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_40 VPB N_Y_c_155_n 5.14916e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_41 N_VPB_c_20_p N_Y_c_155_n 0.00887752f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_42 N_VPB_M1001_b N_Y_c_158_n 0.0165324f $X=-0.33 $Y=1.885 $X2=0.93 $Y2=1.415
cc_43 N_VPB_M1001_b N_Y_c_159_n 0.00249256f $X=-0.33 $Y=1.885 $X2=0.93 $Y2=2.085
cc_44 N_VPB_M1001_b Y 9.581e-19 $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_45 N_VPB_M1001_b Y 0.0661133f $X=-0.33 $Y=1.885 $X2=0.72 $Y2=1.67
cc_46 VPB Y 7.75439e-19 $X=0 $Y=3.955 $X2=0.72 $Y2=1.67
cc_47 N_VPB_c_20_p Y 0.0133691f $X=3.12 $Y=4.07 $X2=0.72 $Y2=1.67
cc_48 N_C_M1001_g N_B_M1004_g 0.0158348f $X=0.895 $Y=2.965 $X2=0 $Y2=0
cc_49 N_C_M1002_g B 0.00143007f $X=0.965 $Y=0.91 $X2=0 $Y2=0
cc_50 N_C_c_49_n N_B_c_70_n 0.0582313f $X=0.83 $Y=1.67 $X2=0 $Y2=0
cc_51 N_C_c_50_n N_B_c_70_n 0.00157627f $X=0.83 $Y=1.67 $X2=0 $Y2=0
cc_52 N_C_M1002_g N_B_c_71_n 0.0582313f $X=0.965 $Y=0.91 $X2=0 $Y2=0
cc_53 N_C_M1001_g N_VPWR_c_128_n 0.0813808f $X=0.895 $Y=2.965 $X2=0.24 $Y2=0
cc_54 N_C_c_50_n N_VPWR_c_128_n 0.0444099f $X=0.83 $Y=1.67 $X2=0.24 $Y2=0
cc_55 N_C_M1001_g N_VPWR_c_134_n 0.00832188f $X=0.895 $Y=2.965 $X2=0 $Y2=0
cc_56 N_C_M1001_g N_Y_c_155_n 0.00364307f $X=0.895 $Y=2.965 $X2=0 $Y2=0
cc_57 N_C_c_49_n N_Y_c_155_n 7.832e-19 $X=0.83 $Y=1.67 $X2=0 $Y2=0
cc_58 N_C_c_49_n N_Y_c_159_n 0.0105913f $X=0.83 $Y=1.67 $X2=3.12 $Y2=0
cc_59 N_C_M1002_g N_VGND_c_194_n 0.0807993f $X=0.965 $Y=0.91 $X2=0 $Y2=0
cc_60 N_C_c_49_n N_VGND_c_194_n 0.00211209f $X=0.83 $Y=1.67 $X2=0 $Y2=0
cc_61 N_C_c_50_n N_VGND_c_194_n 0.0711702f $X=0.83 $Y=1.67 $X2=0 $Y2=0
cc_62 N_B_M1004_g N_A_M1000_g 0.0278157f $X=1.675 $Y=2.965 $X2=0 $Y2=0
cc_63 B A 0.0685158f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_64 N_B_c_70_n A 2.66978e-19 $X=1.97 $Y=1.56 $X2=0 $Y2=0
cc_65 N_B_c_71_n A 3.98781e-19 $X=1.78 $Y=1.395 $X2=0 $Y2=0
cc_66 N_B_c_70_n N_A_c_100_n 0.0353097f $X=1.97 $Y=1.56 $X2=0 $Y2=0
cc_67 B N_A_c_101_n 0.00899683f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_68 N_B_c_71_n N_A_c_101_n 0.0282938f $X=1.78 $Y=1.395 $X2=0 $Y2=0
cc_69 N_B_M1004_g N_VPWR_c_131_n 0.0733167f $X=1.675 $Y=2.965 $X2=0 $Y2=0
cc_70 N_B_M1004_g N_VPWR_c_134_n 0.00803924f $X=1.675 $Y=2.965 $X2=0 $Y2=0
cc_71 N_B_M1004_g N_Y_c_155_n 0.00452076f $X=1.675 $Y=2.965 $X2=0 $Y2=0
cc_72 N_B_M1004_g N_Y_c_158_n 0.039355f $X=1.675 $Y=2.965 $X2=3.12 $Y2=0
cc_73 B N_Y_c_158_n 0.0301759f $X=2.075 $Y=0.84 $X2=3.12 $Y2=0
cc_74 N_B_c_70_n N_Y_c_158_n 0.00623726f $X=1.97 $Y=1.56 $X2=3.12 $Y2=0
cc_75 B VGND 0.0215992f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_76 N_B_c_71_n VGND 0.0140251f $X=1.78 $Y=1.395 $X2=0 $Y2=0
cc_77 B N_VGND_c_194_n 0.0395603f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_78 N_B_c_71_n N_VGND_c_194_n 0.0607659f $X=1.78 $Y=1.395 $X2=0 $Y2=0
cc_79 B A_385_107# 0.0123854f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_80 N_A_M1000_g N_VPWR_c_131_n 0.0988904f $X=2.675 $Y=2.965 $X2=0 $Y2=0
cc_81 N_A_M1000_g N_VPWR_c_134_n 0.00875302f $X=2.675 $Y=2.965 $X2=0 $Y2=0
cc_82 N_A_M1000_g N_Y_c_158_n 0.0386613f $X=2.675 $Y=2.965 $X2=3.12 $Y2=0
cc_83 A N_Y_c_158_n 0.019495f $X=2.555 $Y=0.84 $X2=3.12 $Y2=0
cc_84 N_A_c_100_n N_Y_c_158_n 0.00395599f $X=2.59 $Y=1.56 $X2=3.12 $Y2=0
cc_85 A Y 0.0225269f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_86 N_A_c_100_n Y 0.0192954f $X=2.59 $Y=1.56 $X2=0 $Y2=0
cc_87 N_A_c_101_n Y 0.00185135f $X=2.635 $Y=1.395 $X2=0 $Y2=0
cc_88 N_A_M1000_g Y 0.00974516f $X=2.675 $Y=2.965 $X2=1.68 $Y2=0
cc_89 A N_Y_c_153_n 0.0377151f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_90 N_A_c_101_n N_Y_c_153_n 0.0128032f $X=2.635 $Y=1.395 $X2=0 $Y2=0
cc_91 A VGND 0.0129858f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_92 N_A_c_101_n VGND 0.0266259f $X=2.635 $Y=1.395 $X2=0 $Y2=0
cc_93 N_A_c_101_n N_VGND_c_194_n 0.00220948f $X=2.635 $Y=1.395 $X2=0 $Y2=0
cc_94 N_VPWR_c_134_n N_Y_M1001_d 0.00442064f $X=2.715 $Y=3.59 $X2=0 $Y2=0
cc_95 N_VPWR_c_134_n N_Y_M1000_d 0.00221032f $X=2.715 $Y=3.59 $X2=0 $Y2=0
cc_96 N_VPWR_c_128_n N_Y_c_155_n 0.0676307f $X=0.505 $Y=2.34 $X2=0.24 $Y2=4.07
cc_97 N_VPWR_c_131_n N_Y_c_155_n 0.0630176f $X=2.065 $Y=2.34 $X2=0.24 $Y2=4.07
cc_98 N_VPWR_c_134_n N_Y_c_155_n 0.0229352f $X=2.715 $Y=3.59 $X2=0.24 $Y2=4.07
cc_99 N_VPWR_c_131_n N_Y_c_158_n 0.0891234f $X=2.065 $Y=2.34 $X2=3.12 $Y2=4.07
cc_100 N_VPWR_c_131_n Y 0.0630924f $X=2.065 $Y=2.34 $X2=1.68 $Y2=4.013
cc_101 N_VPWR_c_134_n Y 0.035852f $X=2.715 $Y=3.59 $X2=1.68 $Y2=4.013
cc_102 N_Y_M1005_d VGND 0.00250225f $X=2.845 $Y=0.535 $X2=0 $Y2=0
cc_103 N_Y_c_153_n VGND 0.0361585f $X=2.99 $Y=0.66 $X2=0 $Y2=0
cc_104 N_Y_c_158_n N_VGND_c_194_n 0.00966027f $X=2.98 $Y=1.99 $X2=0 $Y2=0
cc_105 N_Y_c_159_n N_VGND_c_194_n 0.00661618f $X=1.37 $Y=1.99 $X2=0 $Y2=0
cc_106 VGND A_385_107# 0.00620972f $X=0 $Y=0.255 $X2=0 $Y2=0
