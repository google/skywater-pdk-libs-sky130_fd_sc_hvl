* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__nor3_1 A B C VGND VNB VPB VPWR Y
M1000 a_205_443# A VPWR VPB phv w=1.5e+06u l=500000u
+  ad=3.15e+11p pd=3.42e+06u as=4.275e+11p ps=3.57e+06u
M1001 a_347_443# B a_205_443# VPB phv w=1.5e+06u l=500000u
+  ad=3.15e+11p pd=3.42e+06u as=0p ps=0u
M1002 Y C a_347_443# VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=0p ps=0u
M1003 Y A VGND VNB nhv w=750000u l=500000u
+  ad=4.0875e+11p pd=4.09e+06u as=4.0875e+11p ps=4.09e+06u
M1004 Y C VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B Y VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
