* File: sky130_fd_sc_hvl__a22o_1.pex.spice
* Created: Wed Sep  2 09:03:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__A22O_1%VNB 5 7 11 25
r30 7 25 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=0.057
+ $X2=2.64 $Y2=0.058
r31 7 11 0.00134943 $w=5.28e-06 $l=5.7e-08 $layer=MET1_cond $X=2.64 $Y=0.057
+ $X2=2.64 $Y2=0
r32 5 11 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r33 5 11 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__A22O_1%VPB 4 6 14 21
r45 10 21 0.00134943 $w=5.28e-06 $l=5.7e-08 $layer=MET1_cond $X=2.64 $Y=4.07
+ $X2=2.64 $Y2=4.013
r46 10 14 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=4.07
+ $X2=5.04 $Y2=4.07
r47 9 14 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=5.04
+ $Y2=4.07
r48 9 10 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r49 6 21 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=4.012
+ $X2=2.64 $Y2=4.013
r50 4 14 33.0909 $w=1.7e-07 $l=5.08232e-06 $layer=licon1_NTAP_notbjt $count=5
+ $X=0 $Y=3.985 $X2=5.04 $Y2=4.07
r51 4 9 33.0909 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=5
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__A22O_1%A_83_81# 1 2 9 12 13 17 22 23 24 27 29 33 35
+ 37 38
c65 23 0 9.16194e-20 $X=3.385 $Y=0.545
r66 33 38 52.9885 $w=5.2e-07 $l=5.15e-07 $layer=POLY_cond $X=0.675 $Y=1.59
+ $X2=0.675 $Y2=2.105
r67 33 37 20.0636 $w=5.2e-07 $l=1.95e-07 $layer=POLY_cond $X=0.675 $Y=1.59
+ $X2=0.675 $Y2=1.395
r68 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.59 $X2=0.75 $Y2=1.59
r69 29 32 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.75 $Y=1.51 $X2=0.75
+ $Y2=1.59
r70 25 27 1.38293 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=3.51 $Y=0.63 $X2=3.51
+ $Y2=0.66
r71 23 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.385 $Y=0.545
+ $X2=3.51 $Y2=0.63
r72 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.385 $Y=0.545
+ $X2=2.855 $Y2=0.545
r73 22 35 3.70735 $w=2.5e-07 $l=1.28662e-07 $layer=LI1_cond $X=2.77 $Y=1.425
+ $X2=2.677 $Y2=1.51
r74 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=0.63
+ $X2=2.855 $Y2=0.545
r75 21 22 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=2.77 $Y=0.63
+ $X2=2.77 $Y2=1.425
r76 17 19 35.9702 $w=3.28e-07 $l=1.03e-06 $layer=LI1_cond $X=2.665 $Y=2.34
+ $X2=2.665 $Y2=3.37
r77 15 35 3.70735 $w=2.5e-07 $l=9.0802e-08 $layer=LI1_cond $X=2.665 $Y=1.595
+ $X2=2.677 $Y2=1.51
r78 15 17 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=2.665 $Y=1.595
+ $X2=2.665 $Y2=2.34
r79 14 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=1.51
+ $X2=0.75 $Y2=1.51
r80 13 35 2.76166 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=2.5 $Y=1.51
+ $X2=2.677 $Y2=1.51
r81 13 14 103.406 $w=1.68e-07 $l=1.585e-06 $layer=LI1_cond $X=2.5 $Y=1.51
+ $X2=0.915 $Y2=1.51
r82 12 38 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.685 $Y=2.965
+ $X2=0.685 $Y2=2.105
r83 9 37 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.665 $Y=0.91 $X2=0.665
+ $Y2=1.395
r84 2 19 300 $w=1.7e-07 $l=1.223e-06 $layer=licon1_PDIFF $count=2 $X=2.525
+ $Y=2.215 $X2=2.665 $Y2=3.37
r85 2 17 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.525
+ $Y=2.215 $X2=2.665 $Y2=2.34
r86 1 27 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=3.305
+ $Y=0.535 $X2=3.47 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__A22O_1%B2 3 7 9 10 11 12 18 19
c29 18 0 2.77455e-19 $X=2.155 $Y=1.89
r30 18 21 18.987 $w=6.25e-07 $l=1.95e-07 $layer=POLY_cond $X=2.282 $Y=1.89
+ $X2=2.282 $Y2=2.085
r31 18 20 42.9564 $w=6.25e-07 $l=4.75e-07 $layer=POLY_cond $X=2.282 $Y=1.89
+ $X2=2.282 $Y2=1.415
r32 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.155
+ $Y=1.89 $X2=2.155 $Y2=1.89
r33 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.155 $Y=2.775
+ $X2=2.155 $Y2=3.145
r34 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.155 $Y=2.405
+ $X2=2.155 $Y2=2.775
r35 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.155 $Y=2.035
+ $X2=2.155 $Y2=2.405
r36 9 19 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.155 $Y=2.035
+ $X2=2.155 $Y2=1.89
r37 7 20 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.345 $Y=0.91 $X2=2.345
+ $Y2=1.415
r38 3 21 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.275 $Y=2.965
+ $X2=2.275 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_HVL__A22O_1%B1 1 2 3 8 14
c34 1 0 1.96526e-19 $X=3.12 $Y=0.925
r35 11 14 147.668 $w=5e-07 $l=1.38e-06 $layer=POLY_cond $X=3.055 $Y=1.585
+ $X2=3.055 $Y2=2.965
r36 8 11 72.229 $w=5e-07 $l=6.75e-07 $layer=POLY_cond $X=3.055 $Y=0.91 $X2=3.055
+ $Y2=1.585
r37 3 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.12
+ $Y=1.585 $X2=3.12 $Y2=1.585
r38 2 3 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.12 $Y=1.295 $X2=3.12
+ $Y2=1.585
r39 1 2 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=0.925 $X2=3.12
+ $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_HVL__A22O_1%A1 3 7 9 10 11 16
r34 16 19 46.5401 $w=5.25e-07 $l=4.55e-07 $layer=POLY_cond $X=3.847 $Y=1.63
+ $X2=3.847 $Y2=2.085
r35 16 18 22.0816 $w=5.25e-07 $l=2.15e-07 $layer=POLY_cond $X=3.847 $Y=1.63
+ $X2=3.847 $Y2=1.415
r36 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.77
+ $Y=1.63 $X2=3.77 $Y2=1.63
r37 10 11 22.5785 $w=2.43e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.627
+ $X2=4.56 $Y2=1.627
r38 10 17 14.5819 $w=2.43e-07 $l=3.1e-07 $layer=LI1_cond $X=4.08 $Y=1.627
+ $X2=3.77 $Y2=1.627
r39 9 17 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=3.6 $Y=1.627 $X2=3.77
+ $Y2=1.627
r40 7 18 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.86 $Y=0.91 $X2=3.86
+ $Y2=1.415
r41 3 19 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.835 $Y=2.965
+ $X2=3.835 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_HVL__A22O_1%A2 3 7 9 15
c21 3 0 9.16194e-20 $X=4.57 $Y=0.91
r22 13 15 29.9457 $w=6.7e-07 $l=3.75e-07 $layer=POLY_cond $X=4.615 $Y=1.75
+ $X2=4.99 $Y2=1.75
r23 11 13 3.59348 $w=6.7e-07 $l=4.5e-08 $layer=POLY_cond $X=4.57 $Y=1.75
+ $X2=4.615 $Y2=1.75
r24 9 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.63 $X2=4.99 $Y2=1.63
r25 5 13 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.615 $Y=2.085
+ $X2=4.615 $Y2=1.75
r26 5 7 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=4.615 $Y=2.085 $X2=4.615
+ $Y2=2.965
r27 1 11 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.57 $Y=1.415 $X2=4.57
+ $Y2=1.75
r28 1 3 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.57 $Y=1.415 $X2=4.57
+ $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HVL__A22O_1%X 1 2 7 8 9 10 11 12 13 22
r14 13 40 18.6486 $w=2.73e-07 $l=4.45e-07 $layer=LI1_cond $X=0.242 $Y=3.145
+ $X2=0.242 $Y2=3.59
r15 12 13 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.242 $Y=2.775
+ $X2=0.242 $Y2=3.145
r16 11 12 18.2296 $w=2.73e-07 $l=4.35e-07 $layer=LI1_cond $X=0.242 $Y=2.34
+ $X2=0.242 $Y2=2.775
r17 10 11 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.242 $Y=2.035
+ $X2=0.242 $Y2=2.34
r18 9 10 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.242 $Y=1.665
+ $X2=0.242 $Y2=2.035
r19 8 9 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.242 $Y=1.295
+ $X2=0.242 $Y2=1.665
r20 7 8 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.242 $Y=0.925
+ $X2=0.242 $Y2=1.295
r21 7 22 10.2672 $w=2.73e-07 $l=2.45e-07 $layer=LI1_cond $X=0.242 $Y=0.925
+ $X2=0.242 $Y2=0.68
r22 2 40 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.215 $X2=0.295 $Y2=3.59
r23 2 11 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.215 $X2=0.295 $Y2=2.34
r24 1 22 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.535 $X2=0.275 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__A22O_1%VPWR 1 2 7 10 20 27
r39 24 27 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.825 $Y=3.63
+ $X2=4.545 $Y2=3.63
r40 23 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.545 $Y=3.59
+ $X2=4.545 $Y2=3.59
r41 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.825 $Y=3.59
+ $X2=3.825 $Y2=3.59
r42 20 23 15.7316 $w=9.48e-07 $l=1.225e-06 $layer=LI1_cond $X=4.185 $Y=2.365
+ $X2=4.185 $Y2=3.59
r43 14 17 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.65 $Y=3.63
+ $X2=1.37 $Y2=3.63
r44 13 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.37 $Y=3.59
+ $X2=1.37 $Y2=3.59
r45 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.65 $Y=3.59
+ $X2=0.65 $Y2=3.59
r46 10 13 16.9444 $w=8.98e-07 $l=1.25e-06 $layer=LI1_cond $X=1.01 $Y=2.34
+ $X2=1.01 $Y2=3.59
r47 7 24 0.454928 $w=3.7e-07 $l=1.185e-06 $layer=MET1_cond $X=2.64 $Y=3.63
+ $X2=3.825 $Y2=3.63
r48 7 17 0.48756 $w=3.7e-07 $l=1.27e-06 $layer=MET1_cond $X=2.64 $Y=3.63
+ $X2=1.37 $Y2=3.63
r49 2 23 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=4.085
+ $Y=2.215 $X2=4.225 $Y2=3.59
r50 2 20 300 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=2 $X=4.085
+ $Y=2.215 $X2=4.225 $Y2=2.365
r51 1 13 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=0.935
+ $Y=2.215 $X2=1.075 $Y2=3.59
r52 1 10 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.935
+ $Y=2.215 $X2=1.075 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__A22O_1%A_316_443# 1 2 3 12 16 17 21 24 25 28
c50 25 0 8.09284e-20 $X=3.53 $Y=2.015
r51 28 30 42.2562 $w=3.28e-07 $l=1.21e-06 $layer=LI1_cond $X=5.005 $Y=2.36
+ $X2=5.005 $Y2=3.57
r52 26 28 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=5.005 $Y=2.1
+ $X2=5.005 $Y2=2.36
r53 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.84 $Y=2.015
+ $X2=5.005 $Y2=2.1
r54 24 25 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=4.84 $Y=2.015
+ $X2=3.53 $Y2=2.015
r55 21 23 57.6222 $w=2.48e-07 $l=1.25e-06 $layer=LI1_cond $X=3.405 $Y=2.34
+ $X2=3.405 $Y2=3.59
r56 19 23 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=3.405 $Y=3.635
+ $X2=3.405 $Y2=3.59
r57 18 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.405 $Y=2.1
+ $X2=3.53 $Y2=2.015
r58 18 21 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=3.405 $Y=2.1
+ $X2=3.405 $Y2=2.34
r59 16 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.28 $Y=3.72
+ $X2=3.405 $Y2=3.635
r60 16 17 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=3.28 $Y=3.72
+ $X2=1.81 $Y2=3.72
r61 12 15 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=1.725 $Y=2.34
+ $X2=1.725 $Y2=3.59
r62 10 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.725 $Y=3.635
+ $X2=1.81 $Y2=3.72
r63 10 15 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.725 $Y=3.635
+ $X2=1.725 $Y2=3.59
r64 3 30 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=2.215 $X2=5.005 $Y2=3.57
r65 3 28 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=2.215 $X2=5.005 $Y2=2.36
r66 2 23 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=3.305
+ $Y=2.215 $X2=3.445 $Y2=3.59
r67 2 21 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=3.305
+ $Y=2.215 $X2=3.445 $Y2=2.34
r68 1 15 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=1.58
+ $Y=2.215 $X2=1.725 $Y2=3.59
r69 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.58
+ $Y=2.215 $X2=1.725 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__A22O_1%VGND 1 2 7 10 26 27
r34 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.01 $Y=0.48
+ $X2=5.01 $Y2=0.48
r35 24 26 0.635417 $w=9.58e-07 $l=5e-08 $layer=LI1_cond $X=4.96 $Y=0.845
+ $X2=5.01 $Y2=0.845
r36 21 27 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=3.93 $Y=0.44
+ $X2=5.01 $Y2=0.44
r37 20 24 13.0896 $w=9.58e-07 $l=1.03e-06 $layer=LI1_cond $X=3.93 $Y=0.845
+ $X2=4.96 $Y2=0.845
r38 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.93 $Y=0.48
+ $X2=3.93 $Y2=0.48
r39 11 14 0.552824 $w=3.7e-07 $l=1.44e-06 $layer=MET1_cond $X=0.685 $Y=0.44
+ $X2=2.125 $Y2=0.44
r40 10 16 1.28421 $w=1.708e-06 $l=1.8e-07 $layer=LI1_cond $X=1.405 $Y=0.48
+ $X2=1.405 $Y2=0.66
r41 10 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.125 $Y=0.48
+ $X2=2.125 $Y2=0.48
r42 10 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.685 $Y=0.48
+ $X2=0.685 $Y2=0.48
r43 7 21 0.495238 $w=3.7e-07 $l=1.29e-06 $layer=MET1_cond $X=2.64 $Y=0.44
+ $X2=3.93 $Y2=0.44
r44 7 14 0.197711 $w=3.7e-07 $l=5.15e-07 $layer=MET1_cond $X=2.64 $Y=0.44
+ $X2=2.125 $Y2=0.44
r45 2 24 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.82
+ $Y=0.535 $X2=4.96 $Y2=0.66
r46 1 16 60.6667 $w=1.7e-07 $l=1.10073e-06 $layer=licon1_NDIFF $count=3 $X=0.915
+ $Y=0.535 $X2=1.955 $Y2=0.66
r47 1 16 60.6667 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=3 $X=0.915
+ $Y=0.535 $X2=1.055 $Y2=0.66
.ends

