* File: sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1.pxi.spice
* Created: Fri Aug 28 09:37:27 2020
* 
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%VNB N_VNB_M1009_b VNB VNB
+ N_VNB_c_8_p N_VNB_c_50_p VNB VNB
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%VNB
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%VPB N_VPB_M1014_b N_VPB_c_114_p
+ VPB N_VPB_c_171_p N_VPB_c_116_p VPB
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%VPB
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%LVPWR N_LVPWR_M1013_s
+ N_LVPWR_M1002_d N_LVPWR_M1002_b N_LVPWR_c_223_p N_LVPWR_c_211_p
+ N_LVPWR_c_201_p N_LVPWR_c_189_n LVPWR N_LVPWR_c_208_p N_LVPWR_c_187_n LVPWR
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%LVPWR
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_229_967# N_A_229_967#_M1004_s
+ N_A_229_967#_M1006_d N_A_229_967#_M1010_g N_A_229_967#_M1007_g
+ N_A_229_967#_c_256_n N_A_229_967#_M1014_g N_A_229_967#_c_257_n
+ N_A_229_967#_c_251_n N_A_229_967#_c_259_n N_A_229_967#_c_260_n
+ N_A_229_967#_c_272_p N_A_229_967#_c_261_n N_A_229_967#_c_262_n
+ N_A_229_967#_c_263_n PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_229_967#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_507_107# N_A_507_107#_M1011_d
+ N_A_507_107#_M1015_d N_A_507_107#_c_321_n N_A_507_107#_c_322_n
+ N_A_507_107#_c_326_n N_A_507_107#_c_332_p N_A_507_107#_c_342_p
+ N_A_507_107#_c_339_p N_A_507_107#_M1008_g
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_507_107#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_176_993# N_A_176_993#_M1001_s
+ N_A_176_993#_M1008_s N_A_176_993#_M1014_s N_A_176_993#_M1006_g
+ N_A_176_993#_c_364_n N_A_176_993#_c_358_n N_A_176_993#_c_368_n
+ N_A_176_993#_c_359_n N_A_176_993#_c_360_n N_A_176_993#_c_361_n
+ N_A_176_993#_c_362_n N_A_176_993#_c_372_n N_A_176_993#_c_374_n
+ N_A_176_993#_c_376_n N_A_176_993#_c_378_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_176_993#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%SLEEP_B N_SLEEP_B_M1011_g
+ N_SLEEP_B_M1015_g N_SLEEP_B_c_447_n N_SLEEP_B_c_448_n N_SLEEP_B_c_449_n
+ N_SLEEP_B_c_450_n N_SLEEP_B_M1003_g N_SLEEP_B_c_452_n N_SLEEP_B_M1016_g
+ N_SLEEP_B_c_454_n SLEEP_B N_SLEEP_B_c_455_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%SLEEP_B
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_553_1225#
+ N_A_553_1225#_M1009_s N_A_553_1225#_M1002_s N_A_553_1225#_M1004_g
+ N_A_553_1225#_c_504_n N_A_553_1225#_c_505_n N_A_553_1225#_M1012_g
+ N_A_553_1225#_c_507_n N_A_553_1225#_c_508_n N_A_553_1225#_c_509_n
+ N_A_553_1225#_c_510_n N_A_553_1225#_c_511_n N_A_553_1225#_c_512_n
+ N_A_553_1225#_c_513_n N_A_553_1225#_c_514_n N_A_553_1225#_c_515_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_553_1225#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_241_1225#
+ N_A_241_1225#_M1000_d N_A_241_1225#_M1013_d N_A_241_1225#_M1001_g
+ N_A_241_1225#_c_560_n N_A_241_1225#_c_561_n N_A_241_1225#_M1005_g
+ N_A_241_1225#_c_563_n N_A_241_1225#_c_578_n N_A_241_1225#_c_579_n
+ N_A_241_1225#_c_564_n N_A_241_1225#_c_565_n N_A_241_1225#_c_566_n
+ N_A_241_1225#_c_567_n N_A_241_1225#_c_568_n N_A_241_1225#_c_569_n
+ N_A_241_1225#_M1009_g N_A_241_1225#_c_582_n N_A_241_1225#_M1002_g
+ N_A_241_1225#_c_572_n N_A_241_1225#_c_573_n N_A_241_1225#_c_574_n
+ N_A_241_1225#_c_575_n N_A_241_1225#_c_593_n N_A_241_1225#_c_595_n
+ N_A_241_1225#_c_576_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_241_1225#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A N_A_c_675_n N_A_M1013_g
+ N_A_M1000_g N_A_c_672_n N_A_c_673_n A N_A_c_674_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%X N_X_M1010_s N_X_M1007_s
+ N_X_c_694_n N_X_c_700_n N_X_c_695_n N_X_c_697_n X
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%X
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%VPWR N_VPWR_M1007_d
+ N_VPWR_M1014_d N_VPWR_M1015_s N_VPWR_c_712_n N_VPWR_c_713_n N_VPWR_c_714_n
+ N_VPWR_c_715_n N_VPWR_c_717_n N_VPWR_c_719_n VPWR VPWR N_VPWR_c_729_n
+ N_VPWR_c_731_n N_VPWR_c_760_n VPWR VPWR
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%VPWR
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_188_1293#
+ N_A_188_1293#_M1001_d N_A_188_1293#_M1005_d N_A_188_1293#_M1012_d
+ N_A_188_1293#_M1003_d N_A_188_1293#_M1016_d N_A_188_1293#_c_819_n
+ N_A_188_1293#_c_820_n N_A_188_1293#_c_822_n N_A_188_1293#_c_824_n
+ N_A_188_1293#_c_825_n N_A_188_1293#_c_827_n N_A_188_1293#_c_828_n
+ N_A_188_1293#_c_830_n N_A_188_1293#_c_831_n N_A_188_1293#_c_832_n
+ N_A_188_1293#_c_833_n N_A_188_1293#_c_834_n N_A_188_1293#_c_835_n
+ N_A_188_1293#_c_836_n N_A_188_1293#_c_838_n N_A_188_1293#_c_840_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%A_188_1293#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%VGND N_VGND_M1010_d
+ N_VGND_M1008_d N_VGND_M1003_s N_VGND_M1000_s N_VGND_M1009_d N_VGND_c_915_n
+ N_VGND_c_917_n N_VGND_c_918_n N_VGND_c_919_n N_VGND_c_920_n N_VGND_c_921_n
+ VGND VGND N_VGND_c_922_n N_VGND_c_924_n N_VGND_c_926_n N_VGND_c_928_n
+ N_VGND_c_930_n N_VGND_c_932_n N_VGND_c_934_n VGND VGND
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_ISOSRCHVAON_1%VGND
cc_1 N_VNB_M1009_b VPB 0.0940884f $X=-0.33 $Y=-0.265 $X2=0 $Y2=3.955
cc_2 N_VNB_M1009_b N_LVPWR_c_187_n 0.221985f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_3 N_VNB_M1009_b N_A_229_967#_M1010_g 0.080251f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_4 N_VNB_M1009_b N_A_229_967#_c_251_n 0.0114605f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_5 N_VNB_M1009_b N_A_507_107#_c_321_n 0.00652742f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_6 N_VNB_M1009_b N_A_507_107#_c_322_n 0.0188413f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_7 N_VNB_M1009_b N_A_507_107#_M1008_g 0.112035f $X=-0.33 $Y=-0.265 $X2=6.72
+ $Y2=4.07
cc_8 N_VNB_c_8_p N_A_507_107#_M1008_g 0.00257434f $X=13.68 $Y=0 $X2=6.72
+ $Y2=4.07
cc_9 N_VNB_M1009_b N_A_176_993#_c_358_n 0.00370893f $X=-0.33 $Y=-0.265 $X2=0.445
+ $Y2=4.07
cc_10 N_VNB_M1009_b N_A_176_993#_c_359_n 0.00934456f $X=-0.33 $Y=-0.265 $X2=0.6
+ $Y2=4.07
cc_11 N_VNB_M1009_b N_A_176_993#_c_360_n 0.0139924f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1009_b N_A_176_993#_c_361_n 0.00294992f $X=-0.33 $Y=-0.265 $X2=0.6
+ $Y2=4.07
cc_13 N_VNB_M1009_b N_A_176_993#_c_362_n 0.0285726f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_M1009_b N_SLEEP_B_M1011_g 0.0790536f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_15 N_VNB_c_8_p N_SLEEP_B_M1011_g 0.00164919f $X=13.68 $Y=0 $X2=0 $Y2=0
cc_16 N_VNB_M1009_b N_SLEEP_B_c_447_n 0.058037f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_17 N_VNB_M1009_b N_SLEEP_B_c_448_n 0.0925818f $X=-0.33 $Y=-0.265 $X2=0.36
+ $Y2=4.07
cc_18 N_VNB_M1009_b N_SLEEP_B_c_449_n 0.147901f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_19 N_VNB_M1009_b N_SLEEP_B_c_450_n 0.0365987f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_20 N_VNB_M1009_b N_SLEEP_B_M1003_g 0.0365298f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_21 N_VNB_M1009_b N_SLEEP_B_c_452_n 0.124466f $X=-0.33 $Y=-0.265 $X2=0.6
+ $Y2=4.07
cc_22 N_VNB_M1009_b N_SLEEP_B_M1016_g 0.0355997f $X=-0.33 $Y=-0.265 $X2=0.6
+ $Y2=4.07
cc_23 N_VNB_M1009_b N_SLEEP_B_c_454_n 0.0188805f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_24 N_VNB_M1009_b N_SLEEP_B_c_455_n 0.0107327f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_25 N_VNB_M1009_b N_A_553_1225#_M1004_g 0.0422442f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_26 N_VNB_M1009_b N_A_553_1225#_c_504_n 0.0113759f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_27 N_VNB_M1009_b N_A_553_1225#_c_505_n 0.0216544f $X=-0.33 $Y=-0.265 $X2=0.36
+ $Y2=4.07
cc_28 N_VNB_M1009_b N_A_553_1225#_M1012_g 0.0462583f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_29 N_VNB_M1009_b N_A_553_1225#_c_507_n 0.0848416f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_30 N_VNB_M1009_b N_A_553_1225#_c_508_n 0.0668213f $X=-0.33 $Y=-0.265 $X2=0.6
+ $Y2=4.07
cc_31 N_VNB_M1009_b N_A_553_1225#_c_509_n 0.0675514f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_32 N_VNB_M1009_b N_A_553_1225#_c_510_n 0.0180451f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_33 N_VNB_M1009_b N_A_553_1225#_c_511_n 0.0184961f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_M1009_b N_A_553_1225#_c_512_n 0.179745f $X=-0.33 $Y=-0.265 $X2=0.6
+ $Y2=4.07
cc_35 N_VNB_M1009_b N_A_553_1225#_c_513_n 0.0587081f $X=-0.33 $Y=-0.265 $X2=6.72
+ $Y2=4.07
cc_36 N_VNB_M1009_b N_A_553_1225#_c_514_n 0.0528677f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_37 N_VNB_M1009_b N_A_553_1225#_c_515_n 0.0200025f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_38 N_VNB_M1009_b N_A_241_1225#_M1001_g 0.0488142f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_39 N_VNB_M1009_b N_A_241_1225#_c_560_n 0.0115773f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_M1009_b N_A_241_1225#_c_561_n 0.0213036f $X=-0.33 $Y=-0.265 $X2=0.36
+ $Y2=4.07
cc_41 N_VNB_M1009_b N_A_241_1225#_M1005_g 0.0422442f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_42 N_VNB_M1009_b N_A_241_1225#_c_563_n 0.012156f $X=-0.33 $Y=-0.265 $X2=0.445
+ $Y2=4.07
cc_43 N_VNB_M1009_b N_A_241_1225#_c_564_n 0.048705f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_44 N_VNB_M1009_b N_A_241_1225#_c_565_n 0.195832f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_45 N_VNB_M1009_b N_A_241_1225#_c_566_n 0.0108066f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_M1009_b N_A_241_1225#_c_567_n 0.0181728f $X=-0.33 $Y=-0.265 $X2=6.72
+ $Y2=4.07
cc_47 N_VNB_M1009_b N_A_241_1225#_c_568_n 0.0451987f $X=-0.33 $Y=-0.265 $X2=6.72
+ $Y2=4.07
cc_48 N_VNB_M1009_b N_A_241_1225#_c_569_n 0.0183097f $X=-0.33 $Y=-0.265 $X2=6.96
+ $Y2=4.07
cc_49 N_VNB_M1009_b N_A_241_1225#_M1009_g 0.0338135f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_c_50_p N_A_241_1225#_M1009_g 5.5155e-19 $X=13.68 $Y=8.14 $X2=0 $Y2=0
cc_51 N_VNB_M1009_b N_A_241_1225#_c_572_n 0.0221004f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_52 N_VNB_M1009_b N_A_241_1225#_c_573_n 0.0142375f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_53 N_VNB_M1009_b N_A_241_1225#_c_574_n 0.059575f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_54 N_VNB_M1009_b N_A_241_1225#_c_575_n 0.0283209f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_55 N_VNB_M1009_b N_A_241_1225#_c_576_n 0.0794649f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_56 N_VNB_M1009_b N_A_M1000_g 0.0346504f $X=-0.33 $Y=-0.265 $X2=0.445
+ $Y2=4.155
cc_57 N_VNB_c_8_p N_A_M1000_g 5.48702e-19 $X=13.68 $Y=0 $X2=0.445 $Y2=4.155
cc_58 N_VNB_M1009_b N_A_c_672_n 0.0870401f $X=-0.33 $Y=-0.265 $X2=0.445
+ $Y2=4.935
cc_59 N_VNB_M1009_b N_A_c_673_n 0.0200814f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_60 N_VNB_M1009_b N_A_c_674_n 0.0148731f $X=-0.33 $Y=-0.265 $X2=0.24 $Y2=4.07
cc_61 N_VNB_M1009_b N_X_c_694_n 0.00402584f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_62 N_VNB_M1009_b N_X_c_695_n 0.0203437f $X=-0.33 $Y=-0.265 $X2=0.6 $Y2=4.07
cc_63 N_VNB_M1009_b X 0.0262322f $X=-0.33 $Y=-0.265 $X2=6.72 $Y2=4.07
cc_64 N_VNB_M1009_b VPWR 0.116044f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_65 N_VNB_M1009_b VPWR 0.241646f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_66 N_VNB_M1009_b N_A_188_1293#_c_819_n 0.00928749f $X=-0.33 $Y=-0.265
+ $X2=0.445 $Y2=4.07
cc_67 N_VNB_M1009_b N_A_188_1293#_c_820_n 0.107167f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_68 N_VNB_c_50_p N_A_188_1293#_c_820_n 0.00430188f $X=13.68 $Y=8.14 $X2=0
+ $Y2=0
cc_69 N_VNB_M1009_b N_A_188_1293#_c_822_n 0.0182742f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_70 N_VNB_c_50_p N_A_188_1293#_c_822_n 7.03553e-19 $X=13.68 $Y=8.14 $X2=0.24
+ $Y2=4.07
cc_71 N_VNB_M1009_b N_A_188_1293#_c_824_n 0.00829083f $X=-0.33 $Y=-0.265
+ $X2=6.72 $Y2=4.07
cc_72 N_VNB_M1009_b N_A_188_1293#_c_825_n 0.107167f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_73 N_VNB_c_50_p N_A_188_1293#_c_825_n 0.00430188f $X=13.68 $Y=8.14 $X2=0
+ $Y2=0
cc_74 N_VNB_M1009_b N_A_188_1293#_c_827_n 0.00711152f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_75 N_VNB_M1009_b N_A_188_1293#_c_828_n 0.0495784f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_76 N_VNB_c_50_p N_A_188_1293#_c_828_n 0.00193854f $X=13.68 $Y=8.14 $X2=0
+ $Y2=0
cc_77 N_VNB_M1009_b N_A_188_1293#_c_830_n 0.0332819f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_78 N_VNB_M1009_b N_A_188_1293#_c_831_n 0.0578198f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_79 N_VNB_M1009_b N_A_188_1293#_c_832_n 0.00323136f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_80 N_VNB_M1009_b N_A_188_1293#_c_833_n 0.00519817f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_81 N_VNB_M1009_b N_A_188_1293#_c_834_n 0.0197499f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_82 N_VNB_M1009_b N_A_188_1293#_c_835_n 0.00992757f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_83 N_VNB_M1009_b N_A_188_1293#_c_836_n 0.0154258f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_84 N_VNB_c_50_p N_A_188_1293#_c_836_n 7.03553e-19 $X=13.68 $Y=8.14 $X2=0
+ $Y2=0
cc_85 N_VNB_M1009_b N_A_188_1293#_c_838_n 0.0154258f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_86 N_VNB_c_50_p N_A_188_1293#_c_838_n 7.03553e-19 $X=13.68 $Y=8.14 $X2=0
+ $Y2=0
cc_87 N_VNB_M1009_b N_A_188_1293#_c_840_n 0.00296153f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_88 N_VNB_M1009_b N_VGND_c_915_n 0.015144f $X=-0.33 $Y=-0.265 $X2=0.445
+ $Y2=4.07
cc_89 N_VNB_c_8_p N_VGND_c_915_n 6.23864e-19 $X=13.68 $Y=0 $X2=0.445 $Y2=4.07
cc_90 N_VNB_M1009_b N_VGND_c_917_n 0.0187375f $X=-0.33 $Y=-0.265 $X2=0.6
+ $Y2=4.07
cc_91 N_VNB_M1009_b N_VGND_c_918_n 7.42527e-19 $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_92 N_VNB_M1009_b N_VGND_c_919_n 0.0200414f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_93 N_VNB_M1009_b N_VGND_c_920_n 0.0386749f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_94 N_VNB_M1009_b N_VGND_c_921_n 0.0388573f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_95 N_VNB_M1009_b N_VGND_c_922_n 0.0262848f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_96 N_VNB_c_8_p N_VGND_c_922_n 9.92366e-19 $X=13.68 $Y=0 $X2=0 $Y2=0
cc_97 N_VNB_M1009_b N_VGND_c_924_n 0.0308064f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_98 N_VNB_c_8_p N_VGND_c_924_n 0.00162748f $X=13.68 $Y=0 $X2=0 $Y2=0
cc_99 N_VNB_M1009_b N_VGND_c_926_n 0.0412926f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_100 N_VNB_c_8_p N_VGND_c_926_n 0.00162748f $X=13.68 $Y=0 $X2=0 $Y2=0
cc_101 N_VNB_M1009_b N_VGND_c_928_n 0.0399733f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_102 N_VNB_c_8_p N_VGND_c_928_n 0.00162748f $X=13.68 $Y=0 $X2=0 $Y2=0
cc_103 N_VNB_M1009_b N_VGND_c_930_n 0.607661f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_104 N_VNB_c_8_p N_VGND_c_930_n 1.48992f $X=13.68 $Y=0 $X2=0 $Y2=0
cc_105 N_VNB_M1009_b N_VGND_c_932_n 0.0403177f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_106 N_VNB_c_50_p N_VGND_c_932_n 0.00164324f $X=13.68 $Y=8.14 $X2=0 $Y2=0
cc_107 N_VNB_M1009_b N_VGND_c_934_n 0.527793f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_108 N_VNB_c_50_p N_VGND_c_934_n 1.48892f $X=13.68 $Y=8.14 $X2=0 $Y2=0
cc_109 VPB N_LVPWR_M1002_b 0.00912905f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_110 VPB N_LVPWR_c_189_n 0.0480172f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_111 N_VPB_M1014_b N_LVPWR_c_187_n 0.184034f $X=-0.33 $Y=1.885 $X2=13.68
+ $Y2=8.14
cc_112 N_VPB_M1014_b N_A_229_967#_M1010_g 0.239808f $X=-0.33 $Y=1.885 $X2=-0.33
+ $Y2=-0.265
cc_113 N_VPB_c_114_p N_A_229_967#_M1010_g 0.007418f $X=0.445 $Y=4.935 $X2=-0.33
+ $Y2=-0.265
cc_114 VPB N_A_229_967#_M1010_g 0.0203353f $X=0 $Y=3.955 $X2=-0.33 $Y2=-0.265
cc_115 N_VPB_c_116_p N_A_229_967#_M1010_g 0.00289032f $X=0.6 $Y=4.07 $X2=-0.33
+ $Y2=-0.265
cc_116 N_VPB_M1014_b N_A_229_967#_c_256_n 0.0775521f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_117 N_VPB_M1014_b N_A_229_967#_c_257_n 0.0160285f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_118 N_VPB_M1014_b N_A_229_967#_c_251_n 0.0063829f $X=-0.33 $Y=1.885 $X2=13.68
+ $Y2=0
cc_119 N_VPB_M1014_b N_A_229_967#_c_259_n 0.022549f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_120 N_VPB_M1014_b N_A_229_967#_c_260_n 0.0218907f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_121 N_VPB_M1014_b N_A_229_967#_c_261_n 0.0044313f $X=-0.33 $Y=1.885 $X2=13.68
+ $Y2=8.14
cc_122 N_VPB_M1014_b N_A_229_967#_c_262_n 0.00336157f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_123 N_VPB_M1014_b N_A_229_967#_c_263_n 0.110867f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_124 N_VPB_M1014_b N_A_507_107#_c_321_n 0.00662204f $X=-0.33 $Y=1.885
+ $X2=-0.33 $Y2=-0.265
cc_125 N_VPB_M1014_b N_A_507_107#_c_326_n 0.0124911f $X=-0.33 $Y=1.885 $X2=0.24
+ $Y2=0
cc_126 VPB N_A_507_107#_c_326_n 0.00139266f $X=0 $Y=3.955 $X2=0.24 $Y2=0
cc_127 N_VPB_M1014_b N_A_507_107#_M1008_g 0.0523563f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_128 N_VPB_M1014_b N_A_176_993#_M1006_g 0.311338f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=8.025
cc_129 N_VPB_M1014_b N_A_176_993#_c_364_n 0.113863f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_130 VPB N_A_176_993#_c_364_n 0.0442545f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_131 N_VPB_M1014_b N_A_176_993#_c_358_n 0.0392726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_132 N_VPB_c_114_p N_A_176_993#_c_358_n 0.0207253f $X=0.445 $Y=4.935 $X2=0
+ $Y2=0
cc_133 N_VPB_M1014_b N_A_176_993#_c_368_n 0.00595729f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_134 N_VPB_c_114_p N_A_176_993#_c_368_n 0.00870039f $X=0.445 $Y=4.935 $X2=0
+ $Y2=0
cc_135 VPB N_A_176_993#_c_368_n 9.22053e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_136 N_VPB_M1014_b N_A_176_993#_c_362_n 0.0403661f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_137 N_VPB_M1014_b N_A_176_993#_c_372_n 0.039445f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_138 VPB N_A_176_993#_c_372_n 0.023715f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_139 N_VPB_M1014_b N_A_176_993#_c_374_n 0.012052f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_140 VPB N_A_176_993#_c_374_n 0.00752576f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_141 N_VPB_M1014_b N_A_176_993#_c_376_n 0.012063f $X=-0.33 $Y=1.885 $X2=6.72
+ $Y2=0
cc_142 VPB N_A_176_993#_c_376_n 0.00937877f $X=0 $Y=3.955 $X2=6.72 $Y2=0
cc_143 N_VPB_M1014_b N_A_176_993#_c_378_n 0.0240518f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_144 N_VPB_M1014_b N_SLEEP_B_M1015_g 0.0558834f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_145 VPB N_SLEEP_B_M1015_g 0.0101591f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_146 N_VPB_M1014_b N_SLEEP_B_c_447_n 0.0472943f $X=-0.33 $Y=1.885 $X2=-0.33
+ $Y2=-0.265
cc_147 N_VPB_M1014_b N_SLEEP_B_c_448_n 0.0223426f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=8.025
cc_148 VPB N_SLEEP_B_M1003_g 0.0152278f $X=0 $Y=3.955 $X2=0.24 $Y2=0
cc_149 VPB N_SLEEP_B_M1016_g 0.0152278f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_150 N_VPB_M1014_b N_SLEEP_B_c_454_n 0.00444617f $X=-0.33 $Y=1.885 $X2=13.68
+ $Y2=0
cc_151 N_VPB_M1014_b N_SLEEP_B_c_455_n 0.00260186f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_152 N_VPB_M1014_b N_A_241_1225#_c_563_n 0.0102392f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_153 N_VPB_M1014_b N_A_241_1225#_c_578_n 0.169102f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_154 N_VPB_M1014_b N_A_241_1225#_c_579_n 0.00893153f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_155 N_VPB_M1014_b N_A_241_1225#_c_564_n 0.00886596f $X=-0.33 $Y=1.885
+ $X2=13.68 $Y2=0
cc_156 VPB N_A_241_1225#_c_575_n 0.0273935f $X=0 $Y=3.955 $X2=6.96 $Y2=8.14
cc_157 N_VPB_M1014_b N_X_c_697_n 0.0239225f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_158 N_VPB_M1014_b X 0.0173065f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_159 N_VPB_M1014_b N_VPWR_c_712_n 0.0153873f $X=-0.33 $Y=1.885 $X2=0 $Y2=8.025
cc_160 N_VPB_M1014_b N_VPWR_c_713_n 0.0111837f $X=-0.33 $Y=1.885 $X2=0.24 $Y2=0
cc_161 N_VPB_M1014_b N_VPWR_c_714_n 0.00338215f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_162 N_VPB_M1014_b N_VPWR_c_715_n 0.0130763f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_715_n 0.0248012f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_164 N_VPB_M1014_b N_VPWR_c_717_n 0.00774898f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_717_n 0.00102873f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_166 N_VPB_M1014_b N_VPWR_c_719_n 3.9775e-19 $X=-0.33 $Y=1.885 $X2=0.24
+ $Y2=8.14
cc_167 VPB N_VPWR_c_719_n 0.00181684f $X=0 $Y=3.955 $X2=0.24 $Y2=8.14
cc_168 N_VPB_M1014_b VPWR 0.0969117f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_169 VPB VPWR 1.45987f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_170 N_VPB_c_171_p VPWR 0.00524668f $X=0.36 $Y=4.07 $X2=0 $Y2=0
cc_171 N_VPB_M1014_b VPWR 0.0895597f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_172 N_VPB_c_114_p VPWR 0.0392895f $X=0.445 $Y=4.935 $X2=0 $Y2=0
cc_173 VPB VPWR 1.45232f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_174 N_VPB_c_171_p VPWR 0.00275993f $X=0.36 $Y=4.07 $X2=0 $Y2=0
cc_175 N_VPB_c_116_p VPWR 0.00127427f $X=0.6 $Y=4.07 $X2=0 $Y2=0
cc_176 N_VPB_M1014_b N_VPWR_c_729_n 0.014783f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_729_n 0.00200815f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_178 N_VPB_M1014_b N_VPWR_c_731_n 0.013412f $X=-0.33 $Y=1.885 $X2=0.24 $Y2=0
cc_179 VPB N_VPWR_c_731_n 0.00169334f $X=0 $Y=3.955 $X2=0.24 $Y2=0
cc_180 VPB N_A_188_1293#_M1003_d 7.10164e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_181 VPB N_A_188_1293#_M1016_d 7.10164e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_182 VPB N_A_188_1293#_c_833_n 0.0243768f $X=0 $Y=3.955 $X2=0.24 $Y2=8.14
cc_183 VPB N_A_188_1293#_c_835_n 0.02289f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_184 VPB N_VGND_M1003_s 7.42444e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_185 VPB N_VGND_c_919_n 0.0236427f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_186 N_LVPWR_c_187_n N_A_229_967#_M1010_g 0.0382341f $X=9.78 $Y=3.165
+ $X2=-0.33 $Y2=-0.265
cc_187 N_LVPWR_c_187_n N_A_507_107#_M1015_d 0.00214577f $X=9.78 $Y=3.165 $X2=0
+ $Y2=0
cc_188 N_LVPWR_c_187_n N_A_507_107#_c_326_n 0.0377559f $X=9.78 $Y=3.165 $X2=0.24
+ $Y2=0
cc_189 N_LVPWR_c_187_n N_A_176_993#_c_362_n 0.00107082f $X=9.78 $Y=3.165 $X2=0
+ $Y2=0
cc_190 N_LVPWR_c_187_n N_A_176_993#_c_372_n 0.0193689f $X=9.78 $Y=3.165 $X2=0
+ $Y2=0
cc_191 N_LVPWR_c_187_n N_A_176_993#_c_378_n 0.0305351f $X=9.78 $Y=3.165 $X2=0
+ $Y2=0
cc_192 N_LVPWR_c_187_n N_SLEEP_B_M1015_g 0.0308731f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_193 N_LVPWR_c_187_n N_SLEEP_B_M1003_g 0.0373574f $X=9.78 $Y=3.165 $X2=0.24
+ $Y2=0
cc_194 N_LVPWR_c_187_n N_SLEEP_B_M1016_g 0.0373574f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_195 N_LVPWR_M1002_b N_A_553_1225#_c_515_n 0.0543708f $X=8.89 $Y=2.045 $X2=0
+ $Y2=0
cc_196 N_LVPWR_c_201_p N_A_553_1225#_c_515_n 0.0394385f $X=9.87 $Y=4.94 $X2=0
+ $Y2=0
cc_197 N_LVPWR_c_189_n N_A_553_1225#_c_515_n 0.0049861f $X=9.695 $Y=4.07 $X2=0
+ $Y2=0
cc_198 N_LVPWR_M1002_b N_A_241_1225#_c_582_n 0.0210363f $X=8.89 $Y=2.045 $X2=0
+ $Y2=0
cc_199 N_LVPWR_c_201_p N_A_241_1225#_c_582_n 0.0247487f $X=9.87 $Y=4.94 $X2=0
+ $Y2=0
cc_200 N_LVPWR_c_189_n N_A_241_1225#_c_582_n 0.0040027f $X=9.695 $Y=4.07 $X2=0
+ $Y2=0
cc_201 N_LVPWR_M1002_b N_A_241_1225#_c_573_n 0.00929544f $X=8.89 $Y=2.045 $X2=0
+ $Y2=0
cc_202 N_LVPWR_M1002_b N_A_241_1225#_c_574_n 0.0378778f $X=8.89 $Y=2.045 $X2=0
+ $Y2=0
cc_203 N_LVPWR_c_208_p N_A_241_1225#_c_574_n 0.0177293f $X=9.78 $Y=3.165 $X2=0
+ $Y2=0
cc_204 N_LVPWR_c_187_n N_A_241_1225#_c_574_n 0.019656f $X=9.78 $Y=3.165 $X2=0
+ $Y2=0
cc_205 N_LVPWR_M1002_b N_A_241_1225#_c_575_n 0.128322f $X=8.89 $Y=2.045 $X2=6.96
+ $Y2=8.14
cc_206 N_LVPWR_c_211_p N_A_241_1225#_c_575_n 0.0240019f $X=9.73 $Y=3.905
+ $X2=6.96 $Y2=8.14
cc_207 N_LVPWR_c_201_p N_A_241_1225#_c_575_n 0.126534f $X=9.87 $Y=4.94 $X2=6.96
+ $Y2=8.14
cc_208 N_LVPWR_c_189_n N_A_241_1225#_c_575_n 0.0257037f $X=9.695 $Y=4.07
+ $X2=6.96 $Y2=8.14
cc_209 N_LVPWR_M1002_b N_A_241_1225#_c_593_n 0.0111655f $X=8.89 $Y=2.045 $X2=0
+ $Y2=0
cc_210 N_LVPWR_c_187_n N_A_241_1225#_c_593_n 0.0338983f $X=9.78 $Y=3.165 $X2=0
+ $Y2=0
cc_211 N_LVPWR_c_201_p N_A_241_1225#_c_595_n 0.0161088f $X=9.87 $Y=4.94 $X2=0
+ $Y2=0
cc_212 N_LVPWR_c_201_p N_A_241_1225#_c_576_n 0.00691125f $X=9.87 $Y=4.94 $X2=0
+ $Y2=0
cc_213 N_LVPWR_M1002_b N_A_c_675_n 0.020335f $X=8.89 $Y=2.045 $X2=0 $Y2=0
cc_214 N_LVPWR_c_211_p N_A_c_675_n 0.00267857f $X=9.73 $Y=3.905 $X2=0 $Y2=0
cc_215 N_LVPWR_c_189_n N_A_c_675_n 0.00301595f $X=9.695 $Y=4.07 $X2=0 $Y2=0
cc_216 N_LVPWR_c_208_p N_A_c_675_n 0.00649494f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_217 N_LVPWR_c_187_n N_A_c_675_n 0.0115796f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_218 N_LVPWR_c_223_p N_A_c_672_n 0.0068971f $X=9.73 $Y=2.5 $X2=0 $Y2=0
cc_219 N_LVPWR_M1002_b N_A_c_673_n 0.0112699f $X=8.89 $Y=2.045 $X2=-0.33
+ $Y2=-0.265
cc_220 N_LVPWR_c_223_p N_A_c_674_n 0.0161182f $X=9.73 $Y=2.5 $X2=0 $Y2=0
cc_221 N_LVPWR_c_187_n N_X_M1007_s 0.00130208f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_222 N_LVPWR_c_187_n N_X_c_700_n 0.0136661f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_223 N_LVPWR_c_187_n N_X_c_697_n 0.00948348f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_224 N_LVPWR_c_187_n N_VPWR_M1007_d 0.00382442f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_225 N_LVPWR_c_187_n N_VPWR_M1015_s 0.00208078f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_226 N_LVPWR_c_187_n N_VPWR_c_712_n 0.0327037f $X=9.78 $Y=3.165 $X2=0
+ $Y2=8.025
cc_227 N_LVPWR_c_187_n N_VPWR_c_714_n 0.0358445f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_228 N_LVPWR_M1002_b VPWR 0.0188783f $X=8.89 $Y=2.045 $X2=0 $Y2=0
cc_229 N_LVPWR_c_211_p VPWR 0.0388194f $X=9.73 $Y=3.905 $X2=0 $Y2=0
cc_230 N_LVPWR_c_189_n VPWR 0.0151963f $X=9.695 $Y=4.07 $X2=0 $Y2=0
cc_231 N_LVPWR_c_208_p VPWR 0.00401479f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_232 N_LVPWR_c_187_n VPWR 1.45918f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_233 N_LVPWR_M1002_b VPWR 0.0417867f $X=8.89 $Y=2.045 $X2=0 $Y2=0
cc_234 N_LVPWR_c_201_p VPWR 0.0535389f $X=9.87 $Y=4.94 $X2=0 $Y2=0
cc_235 N_LVPWR_c_189_n VPWR 0.0139504f $X=9.695 $Y=4.07 $X2=0 $Y2=0
cc_236 N_LVPWR_c_187_n N_VPWR_c_729_n 0.0030545f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_237 N_LVPWR_c_187_n N_VPWR_c_731_n 0.00296306f $X=9.78 $Y=3.165 $X2=0.24
+ $Y2=0
cc_238 N_LVPWR_c_187_n N_A_188_1293#_M1003_d 0.00214577f $X=9.78 $Y=3.165 $X2=0
+ $Y2=0
cc_239 N_LVPWR_c_187_n N_A_188_1293#_M1016_d 0.00214577f $X=9.78 $Y=3.165 $X2=0
+ $Y2=0
cc_240 N_LVPWR_c_187_n N_A_188_1293#_c_833_n 0.0383201f $X=9.78 $Y=3.165
+ $X2=0.24 $Y2=8.14
cc_241 N_LVPWR_c_189_n N_A_188_1293#_c_835_n 0.0060929f $X=9.695 $Y=4.07 $X2=0
+ $Y2=0
cc_242 N_LVPWR_c_187_n N_A_188_1293#_c_835_n 0.0383201f $X=9.78 $Y=3.165 $X2=0
+ $Y2=0
cc_243 N_LVPWR_c_187_n N_VGND_M1003_s 0.0022433f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_244 N_LVPWR_c_187_n N_VGND_c_919_n 0.0377827f $X=9.78 $Y=3.165 $X2=0 $Y2=0
cc_245 N_A_229_967#_c_256_n N_A_176_993#_M1006_g 0.0172438f $X=2.035 $Y=5.175
+ $X2=0 $Y2=8.025
cc_246 N_A_229_967#_c_259_n N_A_176_993#_M1006_g 0.0435278f $X=5.455 $Y=5.775
+ $X2=0 $Y2=8.025
cc_247 N_A_229_967#_c_260_n N_A_176_993#_M1006_g 0.00965081f $X=5.565 $Y=5.11
+ $X2=0 $Y2=8.025
cc_248 N_A_229_967#_c_262_n N_A_176_993#_M1006_g 0.00258529f $X=3.405 $Y=5.775
+ $X2=0 $Y2=8.025
cc_249 N_A_229_967#_M1010_g N_A_176_993#_c_364_n 0.00997297f $X=1.455 $Y=1.29
+ $X2=0 $Y2=0
cc_250 N_A_229_967#_c_256_n N_A_176_993#_c_364_n 0.0710192f $X=2.035 $Y=5.175
+ $X2=0 $Y2=0
cc_251 N_A_229_967#_M1010_g N_A_176_993#_c_358_n 0.00172901f $X=1.455 $Y=1.29
+ $X2=0 $Y2=0
cc_252 N_A_229_967#_c_272_p N_A_176_993#_c_358_n 0.0199563f $X=1.87 $Y=5.72
+ $X2=0 $Y2=0
cc_253 N_A_229_967#_c_263_n N_A_176_993#_c_358_n 0.0278657f $X=1.59 $Y=5.175
+ $X2=0 $Y2=0
cc_254 N_A_229_967#_c_272_p N_A_176_993#_c_359_n 0.0468407f $X=1.87 $Y=5.72
+ $X2=0 $Y2=0
cc_255 N_A_229_967#_c_263_n N_A_176_993#_c_359_n 0.0101473f $X=1.59 $Y=5.175
+ $X2=0 $Y2=0
cc_256 N_A_229_967#_M1010_g N_A_176_993#_c_362_n 0.0247537f $X=1.455 $Y=1.29
+ $X2=0 $Y2=0
cc_257 N_A_229_967#_M1010_g N_A_176_993#_c_374_n 0.0544508f $X=1.455 $Y=1.29
+ $X2=0 $Y2=0
cc_258 N_A_229_967#_c_263_n N_A_176_993#_c_374_n 0.0230061f $X=1.59 $Y=5.175
+ $X2=0 $Y2=0
cc_259 N_A_229_967#_M1010_g N_A_176_993#_c_376_n 0.00245496f $X=1.455 $Y=1.29
+ $X2=6.72 $Y2=0
cc_260 N_A_229_967#_c_256_n N_A_176_993#_c_376_n 0.0200624f $X=2.035 $Y=5.175
+ $X2=6.72 $Y2=0
cc_261 N_A_229_967#_c_251_n N_A_553_1225#_M1004_g 0.00409313f $X=3.405 $Y=6.61
+ $X2=-0.33 $Y2=-0.265
cc_262 N_A_229_967#_c_251_n N_A_553_1225#_c_504_n 0.0240779f $X=3.405 $Y=6.61
+ $X2=0 $Y2=0
cc_263 N_A_229_967#_c_259_n N_A_553_1225#_c_504_n 0.00991893f $X=5.455 $Y=5.775
+ $X2=0 $Y2=0
cc_264 N_A_229_967#_c_257_n N_A_553_1225#_c_505_n 0.00380491f $X=3.295 $Y=5.775
+ $X2=0 $Y2=8.025
cc_265 N_A_229_967#_c_251_n N_A_553_1225#_M1012_g 0.00409313f $X=3.405 $Y=6.61
+ $X2=0 $Y2=0
cc_266 N_A_229_967#_c_261_n N_A_241_1225#_c_560_n 9.26782e-19 $X=2.035 $Y=5.72
+ $X2=0 $Y2=0
cc_267 N_A_229_967#_c_272_p N_A_241_1225#_c_561_n 3.24684e-19 $X=1.87 $Y=5.72
+ $X2=0 $Y2=8.025
cc_268 N_A_229_967#_c_263_n N_A_241_1225#_c_561_n 0.0472427f $X=1.59 $Y=5.175
+ $X2=0 $Y2=8.025
cc_269 N_A_229_967#_c_257_n N_A_241_1225#_c_578_n 0.0294474f $X=3.295 $Y=5.775
+ $X2=0 $Y2=0
cc_270 N_A_229_967#_c_251_n N_A_241_1225#_c_578_n 0.00519662f $X=3.405 $Y=6.61
+ $X2=0 $Y2=0
cc_271 N_A_229_967#_c_259_n N_A_241_1225#_c_578_n 0.0775093f $X=5.455 $Y=5.775
+ $X2=0 $Y2=0
cc_272 N_A_229_967#_c_262_n N_A_241_1225#_c_578_n 0.00546089f $X=3.405 $Y=5.775
+ $X2=0 $Y2=0
cc_273 N_A_229_967#_c_256_n N_A_241_1225#_c_579_n 0.051994f $X=2.035 $Y=5.175
+ $X2=0 $Y2=0
cc_274 N_A_229_967#_c_257_n N_A_241_1225#_c_579_n 0.0131201f $X=3.295 $Y=5.775
+ $X2=0 $Y2=0
cc_275 N_A_229_967#_c_263_n N_A_241_1225#_c_579_n 0.00720297f $X=1.59 $Y=5.175
+ $X2=0 $Y2=0
cc_276 N_A_229_967#_c_256_n N_A_241_1225#_c_572_n 0.00373733f $X=2.035 $Y=5.175
+ $X2=0 $Y2=0
cc_277 N_A_229_967#_c_257_n N_A_241_1225#_c_572_n 0.00678093f $X=3.295 $Y=5.775
+ $X2=0 $Y2=0
cc_278 N_A_229_967#_M1010_g N_X_c_694_n 6.87047e-19 $X=1.455 $Y=1.29 $X2=-0.33
+ $Y2=-0.265
cc_279 N_A_229_967#_M1010_g N_X_c_697_n 6.78719e-19 $X=1.455 $Y=1.29 $X2=0 $Y2=0
cc_280 N_A_229_967#_M1010_g X 0.0304805f $X=1.455 $Y=1.29 $X2=0 $Y2=0
cc_281 N_A_229_967#_M1010_g N_VPWR_c_712_n 0.0139357f $X=1.455 $Y=1.29 $X2=0
+ $Y2=8.025
cc_282 N_A_229_967#_c_256_n N_VPWR_c_713_n 0.00463212f $X=2.035 $Y=5.175
+ $X2=0.24 $Y2=0
cc_283 N_A_229_967#_c_257_n N_VPWR_c_713_n 0.00756962f $X=3.295 $Y=5.775
+ $X2=0.24 $Y2=0
cc_284 N_A_229_967#_c_262_n N_VPWR_c_713_n 0.00687946f $X=3.405 $Y=5.775
+ $X2=0.24 $Y2=0
cc_285 N_A_229_967#_M1010_g N_VPWR_c_717_n 0.0112163f $X=1.455 $Y=1.29 $X2=0
+ $Y2=0
cc_286 N_A_229_967#_M1010_g VPWR 0.0286549f $X=1.455 $Y=1.29 $X2=0 $Y2=0
cc_287 N_A_229_967#_M1010_g VPWR 0.0140984f $X=1.455 $Y=1.29 $X2=0 $Y2=0
cc_288 N_A_229_967#_c_256_n VPWR 0.00624975f $X=2.035 $Y=5.175 $X2=0 $Y2=0
cc_289 N_A_229_967#_c_260_n VPWR 0.0115415f $X=5.565 $Y=5.11 $X2=0 $Y2=0
cc_290 N_A_229_967#_c_257_n N_A_188_1293#_c_824_n 0.00732086f $X=3.295 $Y=5.775
+ $X2=0 $Y2=0
cc_291 N_A_229_967#_c_251_n N_A_188_1293#_c_824_n 6.41575e-19 $X=3.405 $Y=6.61
+ $X2=0 $Y2=0
cc_292 N_A_229_967#_c_251_n N_A_188_1293#_c_825_n 0.0136171f $X=3.405 $Y=6.61
+ $X2=0 $Y2=0
cc_293 N_A_229_967#_c_251_n N_A_188_1293#_c_827_n 6.41575e-19 $X=3.405 $Y=6.61
+ $X2=13.68 $Y2=8.14
cc_294 N_A_229_967#_c_259_n N_A_188_1293#_c_827_n 0.00728074f $X=5.455 $Y=5.775
+ $X2=13.68 $Y2=8.14
cc_295 N_A_229_967#_c_259_n N_A_188_1293#_c_831_n 0.0283631f $X=5.455 $Y=5.775
+ $X2=6.72 $Y2=0
cc_296 N_A_229_967#_c_259_n N_A_188_1293#_c_832_n 0.0083633f $X=5.455 $Y=5.775
+ $X2=6.96 $Y2=0
cc_297 N_A_229_967#_M1010_g N_VGND_c_917_n 0.00575784f $X=1.455 $Y=1.29 $X2=0
+ $Y2=0
cc_298 N_A_229_967#_M1010_g N_VGND_c_922_n 0.0118486f $X=1.455 $Y=1.29 $X2=0
+ $Y2=0
cc_299 N_A_229_967#_M1010_g N_VGND_c_930_n 0.015856f $X=1.455 $Y=1.29 $X2=0
+ $Y2=0
cc_300 N_A_229_967#_c_251_n N_VGND_c_934_n 0.00761805f $X=3.405 $Y=6.61 $X2=0
+ $Y2=0
cc_301 N_A_507_107#_c_326_n N_A_176_993#_M1006_g 0.00532931f $X=4.315 $Y=2.57
+ $X2=0 $Y2=8.025
cc_302 N_A_507_107#_c_332_p N_A_176_993#_c_362_n 0.0266938f $X=3.155 $Y=1.995
+ $X2=0 $Y2=0
cc_303 N_A_507_107#_M1008_g N_A_176_993#_c_362_n 0.0189301f $X=2.935 $Y=1.165
+ $X2=0 $Y2=0
cc_304 N_A_507_107#_c_322_n N_SLEEP_B_M1011_g 0.0191923f $X=4.315 $Y=0.81 $X2=0
+ $Y2=0
cc_305 N_A_507_107#_M1008_g N_SLEEP_B_M1011_g 0.0420548f $X=2.935 $Y=1.165 $X2=0
+ $Y2=0
cc_306 N_A_507_107#_c_326_n N_SLEEP_B_M1015_g 0.0143848f $X=4.315 $Y=2.57 $X2=0
+ $Y2=0
cc_307 N_A_507_107#_c_321_n N_SLEEP_B_c_447_n 0.00290251f $X=4.205 $Y=2.05
+ $X2=-0.33 $Y2=-0.265
cc_308 N_A_507_107#_c_322_n N_SLEEP_B_c_447_n 0.0129097f $X=4.315 $Y=0.81
+ $X2=-0.33 $Y2=-0.265
cc_309 N_A_507_107#_c_339_p N_SLEEP_B_c_447_n 0.014364f $X=4.315 $Y=2.05
+ $X2=-0.33 $Y2=-0.265
cc_310 N_A_507_107#_c_322_n N_SLEEP_B_c_450_n 0.0235901f $X=4.315 $Y=0.81 $X2=0
+ $Y2=0
cc_311 N_A_507_107#_c_321_n N_SLEEP_B_c_454_n 0.0588792f $X=4.205 $Y=2.05
+ $X2=13.68 $Y2=0
cc_312 N_A_507_107#_c_342_p N_SLEEP_B_c_454_n 7.61715e-19 $X=3.32 $Y=1.995
+ $X2=13.68 $Y2=0
cc_313 N_A_507_107#_c_322_n N_SLEEP_B_c_455_n 0.00525668f $X=4.315 $Y=0.81 $X2=0
+ $Y2=0
cc_314 N_A_507_107#_c_339_p N_SLEEP_B_c_455_n 0.0115536f $X=4.315 $Y=2.05 $X2=0
+ $Y2=0
cc_315 N_A_507_107#_c_321_n N_VPWR_c_714_n 0.0145072f $X=4.205 $Y=2.05 $X2=0
+ $Y2=0
cc_316 N_A_507_107#_c_326_n N_VPWR_c_714_n 0.0033803f $X=4.315 $Y=2.57 $X2=0
+ $Y2=0
cc_317 N_A_507_107#_M1015_d VPWR 0.00222341f $X=4.175 $Y=2.425 $X2=0 $Y2=0
cc_318 N_A_507_107#_c_326_n VPWR 0.0317547f $X=4.315 $Y=2.57 $X2=0 $Y2=0
cc_319 N_A_507_107#_c_326_n N_VPWR_c_760_n 0.00283783f $X=4.315 $Y=2.57 $X2=0
+ $Y2=0
cc_320 N_A_507_107#_M1008_g N_VGND_c_915_n 0.00150144f $X=2.935 $Y=1.165 $X2=0
+ $Y2=0
cc_321 N_A_507_107#_M1008_g N_VGND_c_917_n 0.00224123f $X=2.935 $Y=1.165 $X2=0
+ $Y2=0
cc_322 N_A_507_107#_c_321_n N_VGND_c_918_n 0.0122869f $X=4.205 $Y=2.05 $X2=0
+ $Y2=0
cc_323 N_A_507_107#_c_322_n N_VGND_c_918_n 0.0186066f $X=4.315 $Y=0.81 $X2=0
+ $Y2=0
cc_324 N_A_507_107#_M1008_g N_VGND_c_918_n 0.00115279f $X=2.935 $Y=1.165 $X2=0
+ $Y2=0
cc_325 N_A_507_107#_M1008_g N_VGND_c_924_n 0.0112527f $X=2.935 $Y=1.165 $X2=0
+ $Y2=0
cc_326 N_A_507_107#_c_322_n N_VGND_c_930_n 0.00998275f $X=4.315 $Y=0.81 $X2=0
+ $Y2=0
cc_327 N_A_507_107#_M1008_g N_VGND_c_930_n 0.0474832f $X=2.935 $Y=1.165 $X2=0
+ $Y2=0
cc_328 N_A_176_993#_M1006_g N_SLEEP_B_M1015_g 0.0329689f $X=4.425 $Y=5.175 $X2=0
+ $Y2=0
cc_329 N_A_176_993#_c_361_n N_A_241_1225#_M1001_g 0.00409313f $X=1.845 $Y=6.61
+ $X2=-0.33 $Y2=-0.265
cc_330 N_A_176_993#_c_359_n N_A_241_1225#_c_560_n 0.0131832f $X=1.735 $Y=6.165
+ $X2=0 $Y2=0
cc_331 N_A_176_993#_c_361_n N_A_241_1225#_c_560_n 0.00552251f $X=1.845 $Y=6.61
+ $X2=0 $Y2=0
cc_332 N_A_176_993#_c_359_n N_A_241_1225#_c_561_n 0.0349265f $X=1.735 $Y=6.165
+ $X2=0 $Y2=8.025
cc_333 N_A_176_993#_c_361_n N_A_241_1225#_M1005_g 0.00409313f $X=1.845 $Y=6.61
+ $X2=0 $Y2=0
cc_334 N_A_176_993#_c_359_n N_A_241_1225#_c_563_n 0.00240307f $X=1.735 $Y=6.165
+ $X2=0 $Y2=0
cc_335 N_A_176_993#_M1006_g N_A_241_1225#_c_578_n 0.124133f $X=4.425 $Y=5.175
+ $X2=0 $Y2=0
cc_336 N_A_176_993#_c_362_n N_VPWR_c_712_n 0.0214345f $X=2.395 $Y=0.81 $X2=0
+ $Y2=8.025
cc_337 N_A_176_993#_c_372_n N_VPWR_c_712_n 0.0076976f $X=2.67 $Y=4.295 $X2=0
+ $Y2=8.025
cc_338 N_A_176_993#_c_378_n N_VPWR_c_712_n 0.010357f $X=2.67 $Y=2.972 $X2=0
+ $Y2=8.025
cc_339 N_A_176_993#_M1006_g N_VPWR_c_713_n 0.0141061f $X=4.425 $Y=5.175 $X2=0.24
+ $Y2=0
cc_340 N_A_176_993#_c_364_n N_VPWR_c_713_n 0.00573559f $X=3.425 $Y=4.905
+ $X2=0.24 $Y2=0
cc_341 N_A_176_993#_c_376_n N_VPWR_c_713_n 0.00674734f $X=2.67 $Y=4.545 $X2=0.24
+ $Y2=0
cc_342 N_A_176_993#_c_372_n N_VPWR_c_714_n 0.00718977f $X=2.67 $Y=4.295 $X2=0
+ $Y2=0
cc_343 N_A_176_993#_c_378_n N_VPWR_c_714_n 0.00592812f $X=2.67 $Y=2.972 $X2=0
+ $Y2=0
cc_344 N_A_176_993#_M1006_g N_VPWR_c_715_n 0.0137658f $X=4.425 $Y=5.175 $X2=0
+ $Y2=0
cc_345 N_A_176_993#_c_372_n N_VPWR_c_715_n 0.012223f $X=2.67 $Y=4.295 $X2=0
+ $Y2=0
cc_346 N_A_176_993#_c_376_n N_VPWR_c_715_n 0.00151856f $X=2.67 $Y=4.545 $X2=0
+ $Y2=0
cc_347 N_A_176_993#_M1006_g N_VPWR_c_719_n 0.0149572f $X=4.425 $Y=5.175 $X2=0.24
+ $Y2=8.14
cc_348 N_A_176_993#_c_364_n N_VPWR_c_719_n 0.0148868f $X=3.425 $Y=4.905 $X2=0.24
+ $Y2=8.14
cc_349 N_A_176_993#_c_376_n N_VPWR_c_719_n 0.00513693f $X=2.67 $Y=4.545 $X2=0.24
+ $Y2=8.14
cc_350 N_A_176_993#_c_372_n VPWR 0.0271968f $X=2.67 $Y=4.295 $X2=0 $Y2=0
cc_351 N_A_176_993#_c_378_n VPWR 0.00130244f $X=2.67 $Y=2.972 $X2=0 $Y2=0
cc_352 N_A_176_993#_M1006_g VPWR 0.131589f $X=4.425 $Y=5.175 $X2=0 $Y2=0
cc_353 N_A_176_993#_c_364_n VPWR 0.00727763f $X=3.425 $Y=4.905 $X2=0 $Y2=0
cc_354 N_A_176_993#_c_368_n VPWR 0.0243452f $X=1.115 $Y=4.685 $X2=0 $Y2=0
cc_355 N_A_176_993#_c_372_n VPWR 3.58021e-19 $X=2.67 $Y=4.295 $X2=0 $Y2=0
cc_356 N_A_176_993#_c_374_n VPWR 0.0731742f $X=2.11 $Y=4.545 $X2=0 $Y2=0
cc_357 N_A_176_993#_c_376_n VPWR 0.0606381f $X=2.67 $Y=4.545 $X2=0 $Y2=0
cc_358 N_A_176_993#_c_364_n N_VPWR_c_729_n 0.00371497f $X=3.425 $Y=4.905 $X2=0
+ $Y2=0
cc_359 N_A_176_993#_c_372_n N_VPWR_c_729_n 0.0169761f $X=2.67 $Y=4.295 $X2=0
+ $Y2=0
cc_360 N_A_176_993#_c_376_n N_VPWR_c_729_n 0.00369637f $X=2.67 $Y=4.545 $X2=0
+ $Y2=0
cc_361 N_A_176_993#_c_378_n N_VPWR_c_729_n 0.00303277f $X=2.67 $Y=2.972 $X2=0
+ $Y2=0
cc_362 N_A_176_993#_c_364_n N_VPWR_c_731_n 0.00633079f $X=3.425 $Y=4.905
+ $X2=0.24 $Y2=0
cc_363 N_A_176_993#_c_372_n N_VPWR_c_731_n 0.0127956f $X=2.67 $Y=4.295 $X2=0.24
+ $Y2=0
cc_364 N_A_176_993#_c_359_n N_A_188_1293#_c_819_n 0.00503295f $X=1.735 $Y=6.165
+ $X2=0 $Y2=0
cc_365 N_A_176_993#_c_360_n N_A_188_1293#_c_819_n 0.0148979f $X=1.115 $Y=6.165
+ $X2=0 $Y2=0
cc_366 N_A_176_993#_c_361_n N_A_188_1293#_c_819_n 6.41575e-19 $X=1.845 $Y=6.61
+ $X2=0 $Y2=0
cc_367 N_A_176_993#_c_361_n N_A_188_1293#_c_820_n 0.0136171f $X=1.845 $Y=6.61
+ $X2=13.68 $Y2=0
cc_368 N_A_176_993#_c_361_n N_A_188_1293#_c_824_n 6.41575e-19 $X=1.845 $Y=6.61
+ $X2=0 $Y2=0
cc_369 N_A_176_993#_c_362_n N_VGND_c_917_n 0.0524073f $X=2.395 $Y=0.81 $X2=0
+ $Y2=0
cc_370 N_A_176_993#_c_362_n N_VGND_c_930_n 0.00998275f $X=2.395 $Y=0.81 $X2=0
+ $Y2=0
cc_371 N_A_176_993#_c_361_n N_VGND_c_934_n 0.00761805f $X=1.845 $Y=6.61 $X2=0
+ $Y2=0
cc_372 N_SLEEP_B_M1003_g N_A_241_1225#_c_565_n 0.0359861f $X=7.015 $Y=3.825
+ $X2=13.68 $Y2=0
cc_373 N_SLEEP_B_M1016_g N_A_241_1225#_c_565_n 0.0359861f $X=7.895 $Y=3.825
+ $X2=13.68 $Y2=0
cc_374 N_SLEEP_B_M1016_g N_A_241_1225#_c_569_n 0.00302418f $X=7.895 $Y=3.825
+ $X2=0.24 $Y2=8.14
cc_375 N_SLEEP_B_M1015_g N_VPWR_c_714_n 0.00171116f $X=3.925 $Y=3.175 $X2=0
+ $Y2=0
cc_376 N_SLEEP_B_M1015_g N_VPWR_c_715_n 0.00925806f $X=3.925 $Y=3.175 $X2=0
+ $Y2=0
cc_377 N_SLEEP_B_M1015_g VPWR 0.0154473f $X=3.925 $Y=3.175 $X2=0 $Y2=0
cc_378 N_SLEEP_B_M1003_g VPWR 0.0181736f $X=7.015 $Y=3.825 $X2=0 $Y2=0
cc_379 N_SLEEP_B_M1016_g VPWR 0.0181736f $X=7.895 $Y=3.825 $X2=0 $Y2=0
cc_380 N_SLEEP_B_M1015_g VPWR 4.58359e-19 $X=3.925 $Y=3.175 $X2=0 $Y2=0
cc_381 N_SLEEP_B_M1003_g VPWR 0.0397626f $X=7.015 $Y=3.825 $X2=0 $Y2=0
cc_382 N_SLEEP_B_M1016_g VPWR 0.0397626f $X=7.895 $Y=3.825 $X2=0 $Y2=0
cc_383 N_SLEEP_B_c_449_n N_A_188_1293#_c_833_n 0.00754195f $X=6.715 $Y=1.03
+ $X2=0.24 $Y2=8.14
cc_384 N_SLEEP_B_M1003_g N_A_188_1293#_c_833_n 0.0114929f $X=7.015 $Y=3.825
+ $X2=0.24 $Y2=8.14
cc_385 N_SLEEP_B_M1003_g N_A_188_1293#_c_834_n 0.0440698f $X=7.015 $Y=3.825
+ $X2=6.96 $Y2=8.14
cc_386 N_SLEEP_B_M1016_g N_A_188_1293#_c_834_n 0.0423879f $X=7.895 $Y=3.825
+ $X2=6.96 $Y2=8.14
cc_387 N_SLEEP_B_M1016_g N_A_188_1293#_c_835_n 0.0111671f $X=7.895 $Y=3.825
+ $X2=0 $Y2=0
cc_388 N_SLEEP_B_M1011_g N_VGND_c_918_n 0.0152266f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_389 N_SLEEP_B_M1003_g N_VGND_c_919_n 0.00856748f $X=7.015 $Y=3.825 $X2=0
+ $Y2=0
cc_390 N_SLEEP_B_c_452_n N_VGND_c_919_n 0.0435632f $X=7.895 $Y=1.195 $X2=0 $Y2=0
cc_391 N_SLEEP_B_M1016_g N_VGND_c_919_n 0.00856748f $X=7.895 $Y=3.825 $X2=0
+ $Y2=0
cc_392 N_SLEEP_B_M1011_g N_VGND_c_924_n 0.00768888f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_393 N_SLEEP_B_c_452_n N_VGND_c_926_n 0.0135388f $X=7.895 $Y=1.195 $X2=0 $Y2=0
cc_394 N_SLEEP_B_M1011_g N_VGND_c_930_n 0.0302397f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_395 N_SLEEP_B_c_450_n N_VGND_c_930_n 0.0835489f $X=5.4 $Y=1.03 $X2=0 $Y2=0
cc_396 N_A_553_1225#_M1004_g N_A_241_1225#_M1005_g 0.0135837f $X=3.015 $Y=6.965
+ $X2=0 $Y2=0
cc_397 N_A_553_1225#_c_505_n N_A_241_1225#_c_578_n 0.168241f $X=3.265 $Y=6.215
+ $X2=0 $Y2=0
cc_398 N_A_553_1225#_c_507_n N_A_241_1225#_c_564_n 0.0250618f $X=5.2 $Y=6.215
+ $X2=13.68 $Y2=0
cc_399 N_A_553_1225#_c_511_n N_A_241_1225#_c_565_n 0.0372807f $X=7.915 $Y=7.24
+ $X2=13.68 $Y2=0
cc_400 N_A_553_1225#_c_513_n N_A_241_1225#_c_565_n 0.0218547f $X=9.205 $Y=7.24
+ $X2=13.68 $Y2=0
cc_401 N_A_553_1225#_c_508_n N_A_241_1225#_c_566_n 0.0250618f $X=5.29 $Y=7.225
+ $X2=0 $Y2=0
cc_402 N_A_553_1225#_c_512_n N_A_241_1225#_c_566_n 0.0867719f $X=7.75 $Y=7.24
+ $X2=0 $Y2=0
cc_403 N_A_553_1225#_c_515_n N_A_241_1225#_c_567_n 0.00946615f $X=9.37 $Y=4.94
+ $X2=0 $Y2=0
cc_404 N_A_553_1225#_c_513_n N_A_241_1225#_c_568_n 0.00437638f $X=9.205 $Y=7.24
+ $X2=0 $Y2=0
cc_405 N_A_553_1225#_c_515_n N_A_241_1225#_c_568_n 0.0255574f $X=9.37 $Y=4.94
+ $X2=0 $Y2=0
cc_406 N_A_553_1225#_c_513_n N_A_241_1225#_M1009_g 0.00439373f $X=9.205 $Y=7.24
+ $X2=0 $Y2=0
cc_407 N_A_553_1225#_c_515_n N_A_241_1225#_M1009_g 0.0162867f $X=9.37 $Y=4.94
+ $X2=0 $Y2=0
cc_408 N_A_553_1225#_c_515_n N_A_241_1225#_c_582_n 0.0173558f $X=9.37 $Y=4.94
+ $X2=0 $Y2=0
cc_409 N_A_553_1225#_c_505_n N_A_241_1225#_c_572_n 0.0135837f $X=3.265 $Y=6.215
+ $X2=0 $Y2=0
cc_410 N_A_553_1225#_c_515_n N_A_241_1225#_c_573_n 0.0147868f $X=9.37 $Y=4.94
+ $X2=0 $Y2=0
cc_411 N_A_553_1225#_c_515_n N_A_241_1225#_c_575_n 0.00888683f $X=9.37 $Y=4.94
+ $X2=6.96 $Y2=8.14
cc_412 N_A_553_1225#_c_515_n N_A_241_1225#_c_595_n 0.0261825f $X=9.37 $Y=4.94
+ $X2=0 $Y2=0
cc_413 N_A_553_1225#_c_515_n VPWR 0.0136949f $X=9.37 $Y=4.94 $X2=0 $Y2=0
cc_414 N_A_553_1225#_M1004_g N_A_188_1293#_c_824_n 0.00342455f $X=3.015 $Y=6.965
+ $X2=0 $Y2=0
cc_415 N_A_553_1225#_M1004_g N_A_188_1293#_c_825_n 0.0194561f $X=3.015 $Y=6.965
+ $X2=0 $Y2=0
cc_416 N_A_553_1225#_M1012_g N_A_188_1293#_c_825_n 0.0194561f $X=3.795 $Y=6.965
+ $X2=0 $Y2=0
cc_417 N_A_553_1225#_M1012_g N_A_188_1293#_c_827_n 0.00606773f $X=3.795 $Y=6.965
+ $X2=13.68 $Y2=8.14
cc_418 N_A_553_1225#_c_507_n N_A_188_1293#_c_827_n 0.00434898f $X=5.2 $Y=6.215
+ $X2=13.68 $Y2=8.14
cc_419 N_A_553_1225#_c_508_n N_A_188_1293#_c_830_n 0.0288925f $X=5.29 $Y=7.225
+ $X2=6.72 $Y2=0
cc_420 N_A_553_1225#_c_507_n N_A_188_1293#_c_831_n 0.0110516f $X=5.2 $Y=6.215
+ $X2=6.72 $Y2=0
cc_421 N_A_553_1225#_c_508_n N_A_188_1293#_c_831_n 0.0183164f $X=5.29 $Y=7.225
+ $X2=6.72 $Y2=0
cc_422 N_A_553_1225#_M1012_g N_A_188_1293#_c_832_n 0.00420376f $X=3.795 $Y=6.965
+ $X2=6.96 $Y2=0
cc_423 N_A_553_1225#_c_507_n N_A_188_1293#_c_832_n 0.00912f $X=5.2 $Y=6.215
+ $X2=6.96 $Y2=0
cc_424 N_A_553_1225#_c_513_n N_A_188_1293#_c_834_n 0.0223112f $X=9.205 $Y=7.24
+ $X2=6.96 $Y2=8.14
cc_425 N_A_553_1225#_c_513_n N_VGND_c_921_n 0.0146948f $X=9.205 $Y=7.24 $X2=0
+ $Y2=0
cc_426 N_A_553_1225#_c_515_n N_VGND_c_921_n 0.017638f $X=9.37 $Y=4.94 $X2=0
+ $Y2=0
cc_427 N_A_553_1225#_M1004_g N_VGND_c_934_n 0.0298664f $X=3.015 $Y=6.965 $X2=0
+ $Y2=0
cc_428 N_A_553_1225#_M1012_g N_VGND_c_934_n 0.0306791f $X=3.795 $Y=6.965 $X2=0
+ $Y2=0
cc_429 N_A_553_1225#_c_509_n N_VGND_c_934_n 0.0876966f $X=5.38 $Y=7.315 $X2=0
+ $Y2=0
cc_430 N_A_553_1225#_c_513_n N_VGND_c_934_n 0.0714146f $X=9.205 $Y=7.24 $X2=0
+ $Y2=0
cc_431 N_A_241_1225#_c_574_n N_A_c_675_n 0.0172459f $X=10.23 $Y=0.9 $X2=0 $Y2=0
cc_432 N_A_241_1225#_c_575_n N_A_c_675_n 0.00234456f $X=10.37 $Y=6.125 $X2=0
+ $Y2=0
cc_433 N_A_241_1225#_c_593_n N_A_c_675_n 0.00290158f $X=10.23 $Y=3.2 $X2=0 $Y2=0
cc_434 N_A_241_1225#_c_574_n N_A_M1000_g 0.0214512f $X=10.23 $Y=0.9 $X2=0 $Y2=0
cc_435 N_A_241_1225#_c_574_n N_A_c_673_n 0.0213303f $X=10.23 $Y=0.9 $X2=-0.33
+ $Y2=-0.265
cc_436 N_A_241_1225#_c_574_n N_A_c_674_n 0.0262132f $X=10.23 $Y=0.9 $X2=0 $Y2=0
cc_437 N_A_241_1225#_c_578_n N_VPWR_c_713_n 0.00143768f $X=5.59 $Y=5.825
+ $X2=0.24 $Y2=0
cc_438 N_A_241_1225#_c_575_n VPWR 0.0412306f $X=10.37 $Y=6.125 $X2=0 $Y2=0
cc_439 N_A_241_1225#_c_593_n VPWR 0.00503115f $X=10.23 $Y=3.2 $X2=0 $Y2=0
cc_440 N_A_241_1225#_c_582_n VPWR 0.00924659f $X=9.595 $Y=5.99 $X2=0 $Y2=0
cc_441 N_A_241_1225#_c_575_n VPWR 0.0535389f $X=10.37 $Y=6.125 $X2=0 $Y2=0
cc_442 N_A_241_1225#_M1001_g N_A_188_1293#_c_819_n 0.00606773f $X=1.455 $Y=6.965
+ $X2=0 $Y2=0
cc_443 N_A_241_1225#_M1001_g N_A_188_1293#_c_820_n 0.0194561f $X=1.455 $Y=6.965
+ $X2=13.68 $Y2=0
cc_444 N_A_241_1225#_M1005_g N_A_188_1293#_c_820_n 0.0194561f $X=2.235 $Y=6.965
+ $X2=13.68 $Y2=0
cc_445 N_A_241_1225#_M1005_g N_A_188_1293#_c_824_n 0.00342455f $X=2.235 $Y=6.965
+ $X2=0 $Y2=0
cc_446 N_A_241_1225#_c_578_n N_A_188_1293#_c_824_n 0.00265986f $X=5.59 $Y=5.825
+ $X2=0 $Y2=0
cc_447 N_A_241_1225#_c_578_n N_A_188_1293#_c_827_n 5.76597e-19 $X=5.59 $Y=5.825
+ $X2=13.68 $Y2=8.14
cc_448 N_A_241_1225#_c_578_n N_A_188_1293#_c_831_n 0.00329947f $X=5.59 $Y=5.825
+ $X2=6.72 $Y2=0
cc_449 N_A_241_1225#_c_564_n N_A_188_1293#_c_831_n 0.0244388f $X=5.68 $Y=6.665
+ $X2=6.72 $Y2=0
cc_450 N_A_241_1225#_c_565_n N_A_188_1293#_c_831_n 0.0222477f $X=8.75 $Y=6.755
+ $X2=6.72 $Y2=0
cc_451 N_A_241_1225#_c_578_n N_A_188_1293#_c_832_n 5.43119e-19 $X=5.59 $Y=5.825
+ $X2=6.96 $Y2=0
cc_452 N_A_241_1225#_c_578_n N_A_188_1293#_c_833_n 0.0124254f $X=5.59 $Y=5.825
+ $X2=0.24 $Y2=8.14
cc_453 N_A_241_1225#_c_565_n N_A_188_1293#_c_834_n 0.0386474f $X=8.75 $Y=6.755
+ $X2=6.96 $Y2=8.14
cc_454 N_A_241_1225#_c_569_n N_A_188_1293#_c_834_n 0.00658137f $X=8.93 $Y=6.365
+ $X2=6.96 $Y2=8.14
cc_455 N_A_241_1225#_c_569_n N_A_188_1293#_c_835_n 4.36573e-19 $X=8.93 $Y=6.365
+ $X2=0 $Y2=0
cc_456 N_A_241_1225#_c_565_n N_A_188_1293#_c_840_n 0.00940321f $X=8.75 $Y=6.755
+ $X2=0 $Y2=0
cc_457 N_A_241_1225#_c_574_n N_VGND_c_920_n 0.0308485f $X=10.23 $Y=0.9 $X2=0
+ $Y2=0
cc_458 N_A_241_1225#_M1009_g N_VGND_c_921_n 0.0200849f $X=9.585 $Y=7.015 $X2=0
+ $Y2=0
cc_459 N_A_241_1225#_c_595_n N_VGND_c_921_n 0.0276613f $X=10.21 $Y=6.29 $X2=0
+ $Y2=0
cc_460 N_A_241_1225#_c_576_n N_VGND_c_921_n 0.00764098f $X=10.21 $Y=6.29 $X2=0
+ $Y2=0
cc_461 N_A_241_1225#_c_574_n N_VGND_c_930_n 0.0137111f $X=10.23 $Y=0.9 $X2=0
+ $Y2=0
cc_462 N_A_241_1225#_M1001_g N_VGND_c_934_n 0.0306791f $X=1.455 $Y=6.965 $X2=0
+ $Y2=0
cc_463 N_A_241_1225#_M1005_g N_VGND_c_934_n 0.0298664f $X=2.235 $Y=6.965 $X2=0
+ $Y2=0
cc_464 N_A_241_1225#_M1009_g N_VGND_c_934_n 0.00798778f $X=9.585 $Y=7.015 $X2=0
+ $Y2=0
cc_465 N_A_c_675_n VPWR 0.00428181f $X=10.005 $Y=2.15 $X2=0 $Y2=0
cc_466 N_A_M1000_g N_VGND_c_920_n 0.0199091f $X=10.015 $Y=1.125 $X2=0 $Y2=0
cc_467 N_A_c_672_n N_VGND_c_920_n 0.00764098f $X=9.915 $Y=1.85 $X2=0 $Y2=0
cc_468 N_A_c_674_n N_VGND_c_920_n 0.0276613f $X=9.73 $Y=1.85 $X2=0 $Y2=0
cc_469 N_A_M1000_g N_VGND_c_930_n 0.00523016f $X=10.015 $Y=1.125 $X2=0 $Y2=0
cc_470 N_X_c_700_n N_VPWR_c_712_n 4.93218e-19 $X=1.065 $Y=2.91 $X2=0 $Y2=8.025
cc_471 N_X_c_697_n N_VPWR_c_712_n 6.08073e-19 $X=1.065 $Y=2.57 $X2=0 $Y2=8.025
cc_472 N_X_c_700_n VPWR 0.00100963f $X=1.065 $Y=2.91 $X2=0 $Y2=0
cc_473 N_X_c_694_n N_VGND_c_917_n 6.2289e-19 $X=1.065 $Y=1.06 $X2=0 $Y2=0
cc_474 N_X_c_694_n N_VGND_c_930_n 0.0107813f $X=1.065 $Y=1.06 $X2=0 $Y2=0
cc_475 VPWR N_A_188_1293#_M1003_d 7.12537e-19 $X=0 $Y=3.445 $X2=0 $Y2=0
cc_476 VPWR N_A_188_1293#_M1003_d 0.00219125f $X=0 $Y=4.325 $X2=0 $Y2=0
cc_477 VPWR N_A_188_1293#_M1016_d 7.12537e-19 $X=0 $Y=3.445 $X2=0 $Y2=0
cc_478 VPWR N_A_188_1293#_M1016_d 0.00219125f $X=0 $Y=4.325 $X2=0 $Y2=0
cc_479 VPWR N_A_188_1293#_c_833_n 0.0358238f $X=0 $Y=3.445 $X2=0.24 $Y2=8.14
cc_480 VPWR N_A_188_1293#_c_833_n 0.0454973f $X=0 $Y=4.325 $X2=0.24 $Y2=8.14
cc_481 VPWR N_A_188_1293#_c_835_n 0.0358238f $X=0 $Y=3.445 $X2=0 $Y2=0
cc_482 VPWR N_A_188_1293#_c_835_n 0.0454973f $X=0 $Y=4.325 $X2=0 $Y2=0
cc_483 VPWR N_VGND_M1003_s 7.44925e-19 $X=0 $Y=3.445 $X2=0 $Y2=0
cc_484 VPWR N_VGND_M1003_s 0.00229085f $X=0 $Y=4.325 $X2=0 $Y2=0
cc_485 VPWR N_VGND_c_919_n 0.0344873f $X=0 $Y=3.445 $X2=0 $Y2=0
cc_486 VPWR N_VGND_c_919_n 0.0446046f $X=0 $Y=4.325 $X2=0 $Y2=0
cc_487 N_A_188_1293#_c_834_n N_VGND_M1003_s 0.0020735f $X=8.225 $Y=6.405 $X2=0
+ $Y2=0
cc_488 N_A_188_1293#_c_833_n N_VGND_c_919_n 0.0100222f $X=6.575 $Y=1.47 $X2=0
+ $Y2=0
cc_489 N_A_188_1293#_c_834_n N_VGND_c_919_n 0.0106431f $X=8.225 $Y=6.405 $X2=0
+ $Y2=0
cc_490 N_A_188_1293#_c_835_n N_VGND_c_919_n 0.0100222f $X=8.335 $Y=1.47 $X2=0
+ $Y2=0
cc_491 N_A_188_1293#_c_819_n N_VGND_c_934_n 0.0227121f $X=1.065 $Y=6.61 $X2=0
+ $Y2=0
cc_492 N_A_188_1293#_c_820_n N_VGND_c_934_n 0.0667646f $X=2.515 $Y=7.735 $X2=0
+ $Y2=0
cc_493 N_A_188_1293#_c_822_n N_VGND_c_934_n 0.0139725f $X=1.175 $Y=7.735 $X2=0
+ $Y2=0
cc_494 N_A_188_1293#_c_824_n N_VGND_c_934_n 0.0227121f $X=2.625 $Y=6.61 $X2=0
+ $Y2=0
cc_495 N_A_188_1293#_c_825_n N_VGND_c_934_n 0.0667646f $X=4.075 $Y=7.735 $X2=0
+ $Y2=0
cc_496 N_A_188_1293#_c_827_n N_VGND_c_934_n 0.0210219f $X=4.185 $Y=6.61 $X2=0
+ $Y2=0
cc_497 N_A_188_1293#_c_828_n N_VGND_c_934_n 0.0342788f $X=4.68 $Y=7.735 $X2=0
+ $Y2=0
cc_498 N_A_188_1293#_c_830_n N_VGND_c_934_n 0.0210219f $X=4.79 $Y=7.625 $X2=0
+ $Y2=0
cc_499 N_A_188_1293#_c_836_n N_VGND_c_934_n 0.00632071f $X=2.625 $Y=7.735 $X2=0
+ $Y2=0
cc_500 N_A_188_1293#_c_838_n N_VGND_c_934_n 0.00632071f $X=4.185 $Y=7.735 $X2=0
+ $Y2=0
