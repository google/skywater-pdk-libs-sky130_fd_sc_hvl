* File: sky130_fd_sc_hvl__and2_1.pxi.spice
* Created: Wed Sep  2 09:03:37 2020
* 
x_PM_SKY130_FD_SC_HVL__AND2_1%VNB N_VNB_M1005_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__AND2_1%VNB
x_PM_SKY130_FD_SC_HVL__AND2_1%VPB N_VPB_M1001_b VPB N_VPB_c_29_p VPB
+ PM_SKY130_FD_SC_HVL__AND2_1%VPB
x_PM_SKY130_FD_SC_HVL__AND2_1%A N_A_M1005_g N_A_M1001_g N_A_c_49_n N_A_c_53_n A
+ A N_A_c_51_n PM_SKY130_FD_SC_HVL__AND2_1%A
x_PM_SKY130_FD_SC_HVL__AND2_1%B N_B_c_81_n N_B_M1004_g N_B_M1003_g B B
+ N_B_c_85_n PM_SKY130_FD_SC_HVL__AND2_1%B
x_PM_SKY130_FD_SC_HVL__AND2_1%A_30_107# N_A_30_107#_M1005_s N_A_30_107#_M1001_d
+ N_A_30_107#_M1000_g N_A_30_107#_M1002_g N_A_30_107#_c_121_n
+ N_A_30_107#_c_123_n N_A_30_107#_c_124_n N_A_30_107#_c_140_n
+ N_A_30_107#_c_129_n N_A_30_107#_c_146_n N_A_30_107#_c_130_n
+ N_A_30_107#_c_131_n N_A_30_107#_c_132_n N_A_30_107#_c_163_n
+ N_A_30_107#_c_125_n PM_SKY130_FD_SC_HVL__AND2_1%A_30_107#
x_PM_SKY130_FD_SC_HVL__AND2_1%VPWR N_VPWR_M1001_s N_VPWR_M1003_d VPWR
+ N_VPWR_c_184_n N_VPWR_c_187_n N_VPWR_c_190_n PM_SKY130_FD_SC_HVL__AND2_1%VPWR
x_PM_SKY130_FD_SC_HVL__AND2_1%X N_X_M1002_d N_X_M1000_d X X X X X X X
+ N_X_c_209_n PM_SKY130_FD_SC_HVL__AND2_1%X
x_PM_SKY130_FD_SC_HVL__AND2_1%VGND N_VGND_M1004_d VGND N_VGND_c_225_n
+ N_VGND_c_227_n PM_SKY130_FD_SC_HVL__AND2_1%VGND
cc_1 N_VNB_M1005_b N_A_M1005_g 0.0560659f $X=-0.33 $Y=-0.265 $X2=0.665 $Y2=0.745
cc_2 N_VNB_c_2_p N_A_M1005_g 0.0023273f $X=0.24 $Y=0 $X2=0.665 $Y2=0.745
cc_3 N_VNB_M1005_b N_A_c_49_n 0.0563243f $X=-0.33 $Y=-0.265 $X2=0.672 $Y2=1.95
cc_4 N_VNB_M1005_b A 0.0272617f $X=-0.33 $Y=-0.265 $X2=0.155 $Y2=1.21
cc_5 N_VNB_M1005_b N_A_c_51_n 0.0511455f $X=-0.33 $Y=-0.265 $X2=0.385 $Y2=1.34
cc_6 N_VNB_M1005_b N_B_c_81_n 0.050684f $X=-0.33 $Y=-0.265 $X2=0.557 $Y2=1.442
cc_7 N_VNB_c_2_p N_B_c_81_n 0.0023273f $X=0.24 $Y=0 $X2=0.557 $Y2=1.442
cc_8 N_VNB_M1005_b N_B_M1003_g 0.0155423f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_M1005_b B 0.00511152f $X=-0.33 $Y=-0.265 $X2=0.895 $Y2=2.425
cc_10 N_VNB_M1005_b N_B_c_85_n 0.097544f $X=-0.33 $Y=-0.265 $X2=0.385 $Y2=1.34
cc_11 N_VNB_M1005_b N_A_30_107#_M1002_g 0.0525102f $X=-0.33 $Y=-0.265 $X2=0.155
+ $Y2=1.58
cc_12 N_VNB_c_2_p N_A_30_107#_M1002_g 0.00149413f $X=0.24 $Y=0 $X2=0.155
+ $Y2=1.58
cc_13 N_VNB_M1005_b N_A_30_107#_c_121_n 0.0185704f $X=-0.33 $Y=-0.265 $X2=0.385
+ $Y2=1.34
cc_14 N_VNB_c_2_p N_A_30_107#_c_121_n 5.84425e-19 $X=0.24 $Y=0 $X2=0.385
+ $Y2=1.34
cc_15 N_VNB_M1005_b N_A_30_107#_c_123_n 2.01423e-19 $X=-0.33 $Y=-0.265 $X2=0.557
+ $Y2=1.085
cc_16 N_VNB_M1005_b N_A_30_107#_c_124_n 0.00890956f $X=-0.33 $Y=-0.265 $X2=0.33
+ $Y2=1.295
cc_17 N_VNB_M1005_b N_A_30_107#_c_125_n 0.0506835f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1005_b N_X_c_209_n 0.0702124f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_19 N_VNB_c_2_p N_X_c_209_n 6.39784e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_20 N_VNB_M1005_b N_VGND_c_225_n 0.0643722f $X=-0.33 $Y=-0.265 $X2=0.895
+ $Y2=2.105
cc_21 N_VNB_c_2_p N_VGND_c_225_n 0.00280401f $X=0.24 $Y=0 $X2=0.895 $Y2=2.105
cc_22 N_VNB_M1005_b N_VGND_c_227_n 0.0734326f $X=-0.33 $Y=-0.265 $X2=0.672
+ $Y2=2.105
cc_23 N_VNB_c_2_p N_VGND_c_227_n 0.359498f $X=0.24 $Y=0 $X2=0.672 $Y2=2.105
cc_24 N_VPB_M1001_b N_A_c_49_n 0.00985739f $X=-0.33 $Y=1.885 $X2=0.672 $Y2=1.95
cc_25 N_VPB_M1001_b N_A_c_53_n 0.0885133f $X=-0.33 $Y=1.885 $X2=0.672 $Y2=2.105
cc_26 N_VPB_M1001_b N_B_M1003_g 0.0608308f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_27 N_VPB_M1001_b N_A_30_107#_M1000_g 0.0429733f $X=-0.33 $Y=1.885 $X2=0.895
+ $Y2=2.425
cc_28 VPB N_A_30_107#_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.895 $Y2=2.425
cc_29 N_VPB_c_29_p N_A_30_107#_M1000_g 0.0152133f $X=3.12 $Y=4.07 $X2=0.895
+ $Y2=2.425
cc_30 N_VPB_M1001_b N_A_30_107#_c_129_n 0.00804448f $X=-0.33 $Y=1.885 $X2=0.33
+ $Y2=1.34
cc_31 N_VPB_M1001_b N_A_30_107#_c_130_n 0.0100565f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_32 N_VPB_M1001_b N_A_30_107#_c_131_n 0.015526f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_33 N_VPB_M1001_b N_A_30_107#_c_132_n 0.00105788f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_34 N_VPB_M1001_b N_A_30_107#_c_125_n 0.0212253f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_35 N_VPB_M1001_b N_VPWR_c_184_n 0.105628f $X=-0.33 $Y=1.885 $X2=0.672
+ $Y2=1.95
cc_36 VPB N_VPWR_c_184_n 0.00263373f $X=0 $Y=3.955 $X2=0.672 $Y2=1.95
cc_37 N_VPB_c_29_p N_VPWR_c_184_n 0.0401319f $X=3.12 $Y=4.07 $X2=0.672 $Y2=1.95
cc_38 N_VPB_M1001_b N_VPWR_c_187_n 0.0303717f $X=-0.33 $Y=1.885 $X2=0.557
+ $Y2=1.085
cc_39 VPB N_VPWR_c_187_n 0.00447364f $X=0 $Y=3.955 $X2=0.557 $Y2=1.085
cc_40 N_VPB_c_29_p N_VPWR_c_187_n 0.0644672f $X=3.12 $Y=4.07 $X2=0.557 $Y2=1.085
cc_41 N_VPB_M1001_b N_VPWR_c_190_n 0.07185f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_190_n 0.35834f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_43 N_VPB_c_29_p N_VPWR_c_190_n 0.0157795f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_44 N_VPB_M1001_b N_X_c_209_n 0.0708798f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_45 VPB N_X_c_209_n 8.36738e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_46 N_VPB_c_29_p N_X_c_209_n 0.014426f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_47 N_A_M1005_g N_B_c_81_n 0.0458183f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_48 N_A_c_49_n N_B_M1003_g 0.00577517f $X=0.672 $Y=1.95 $X2=0 $Y2=0
cc_49 N_A_c_53_n N_B_M1003_g 0.0189105f $X=0.672 $Y=2.105 $X2=0 $Y2=0
cc_50 N_A_M1005_g B 0.00634892f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_51 N_A_c_53_n B 4.30373e-19 $X=0.672 $Y=2.105 $X2=0 $Y2=0
cc_52 N_A_c_53_n N_B_c_85_n 0.00132975f $X=0.672 $Y=2.105 $X2=3.12 $Y2=0
cc_53 N_A_c_51_n N_B_c_85_n 0.0458183f $X=0.385 $Y=1.34 $X2=3.12 $Y2=0
cc_54 N_A_M1005_g N_A_30_107#_c_121_n 0.00262285f $X=0.665 $Y=0.745 $X2=3.12
+ $Y2=0
cc_55 N_A_M1005_g N_A_30_107#_c_123_n 0.0264878f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_56 A N_A_30_107#_c_123_n 0.0108632f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_57 N_A_c_51_n N_A_30_107#_c_123_n 0.00101475f $X=0.385 $Y=1.34 $X2=0 $Y2=0
cc_58 A N_A_30_107#_c_124_n 0.0204357f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_59 N_A_c_51_n N_A_30_107#_c_124_n 0.00537387f $X=0.385 $Y=1.34 $X2=0 $Y2=0
cc_60 N_A_M1005_g N_A_30_107#_c_140_n 0.00539106f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_61 N_A_c_49_n N_A_30_107#_c_140_n 0.0197992f $X=0.672 $Y=1.95 $X2=0 $Y2=0
cc_62 A N_A_30_107#_c_140_n 0.0464444f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_63 N_A_c_51_n N_A_30_107#_c_140_n 0.0151074f $X=0.385 $Y=1.34 $X2=0 $Y2=0
cc_64 N_A_c_49_n N_A_30_107#_c_129_n 0.00218365f $X=0.672 $Y=1.95 $X2=1.68
+ $Y2=0.057
cc_65 N_A_c_53_n N_A_30_107#_c_129_n 0.0151257f $X=0.672 $Y=2.105 $X2=1.68
+ $Y2=0.057
cc_66 N_A_c_49_n N_A_30_107#_c_146_n 0.00285714f $X=0.672 $Y=1.95 $X2=1.68
+ $Y2=0.058
cc_67 N_A_c_53_n N_A_30_107#_c_146_n 0.010648f $X=0.672 $Y=2.105 $X2=1.68
+ $Y2=0.058
cc_68 N_A_c_53_n N_A_30_107#_c_130_n 0.00399883f $X=0.672 $Y=2.105 $X2=0 $Y2=0
cc_69 N_A_c_53_n N_VPWR_c_184_n 0.0582298f $X=0.672 $Y=2.105 $X2=0.24 $Y2=0
cc_70 A N_VPWR_c_184_n 0.0187637f $X=0.155 $Y=1.21 $X2=0.24 $Y2=0
cc_71 N_A_c_53_n N_VPWR_c_187_n 4.47923e-19 $X=0.672 $Y=2.105 $X2=0 $Y2=0
cc_72 N_A_M1005_g N_VGND_c_227_n 0.018715f $X=0.665 $Y=0.745 $X2=0.24 $Y2=0
cc_73 A N_VGND_c_227_n 0.00111256f $X=0.155 $Y=1.21 $X2=0.24 $Y2=0
cc_74 N_B_M1003_g N_A_30_107#_M1000_g 0.0182556f $X=1.675 $Y=2.425 $X2=0 $Y2=0
cc_75 N_B_c_85_n N_A_30_107#_M1002_g 0.00591666f $X=1.675 $Y=1.402 $X2=0 $Y2=0
cc_76 B N_A_30_107#_c_123_n 0.0136282f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_77 N_B_c_81_n N_A_30_107#_c_140_n 7.69232e-19 $X=1.375 $Y=1.065 $X2=0 $Y2=0
cc_78 N_B_M1003_g N_A_30_107#_c_140_n 9.87195e-19 $X=1.675 $Y=2.425 $X2=0 $Y2=0
cc_79 B N_A_30_107#_c_140_n 0.0534579f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_80 B N_A_30_107#_c_129_n 0.0104865f $X=1.115 $Y=0.84 $X2=1.68 $Y2=0.057
cc_81 N_B_c_85_n N_A_30_107#_c_129_n 0.00158264f $X=1.675 $Y=1.402 $X2=1.68
+ $Y2=0.057
cc_82 N_B_M1003_g N_A_30_107#_c_130_n 0.00398996f $X=1.675 $Y=2.425 $X2=0 $Y2=0
cc_83 N_B_M1003_g N_A_30_107#_c_131_n 0.0402205f $X=1.675 $Y=2.425 $X2=0 $Y2=0
cc_84 B N_A_30_107#_c_131_n 0.00628149f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_85 N_B_c_85_n N_A_30_107#_c_131_n 0.00146185f $X=1.675 $Y=1.402 $X2=0 $Y2=0
cc_86 B N_A_30_107#_c_132_n 0.0145113f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_87 N_B_c_85_n N_A_30_107#_c_132_n 0.00468389f $X=1.675 $Y=1.402 $X2=0 $Y2=0
cc_88 N_B_c_85_n N_A_30_107#_c_163_n 0.00110847f $X=1.675 $Y=1.402 $X2=0 $Y2=0
cc_89 N_B_c_85_n N_A_30_107#_c_125_n 0.0182556f $X=1.675 $Y=1.402 $X2=0 $Y2=0
cc_90 N_B_M1003_g N_VPWR_c_184_n 4.47923e-19 $X=1.675 $Y=2.425 $X2=0.24 $Y2=0
cc_91 N_B_M1003_g N_VPWR_c_187_n 0.0468908f $X=1.675 $Y=2.425 $X2=0 $Y2=0
cc_92 B A_183_107# 0.00132067f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_93 N_B_c_81_n N_VGND_c_225_n 0.0105486f $X=1.375 $Y=1.065 $X2=0 $Y2=0
cc_94 B N_VGND_c_225_n 0.0341716f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_95 N_B_c_85_n N_VGND_c_225_n 0.03089f $X=1.675 $Y=1.402 $X2=0 $Y2=0
cc_96 N_B_c_81_n N_VGND_c_227_n 0.0237489f $X=1.375 $Y=1.065 $X2=0.24 $Y2=0
cc_97 B N_VGND_c_227_n 0.0192137f $X=1.115 $Y=0.84 $X2=0.24 $Y2=0
cc_98 N_B_c_85_n N_VGND_c_227_n 2.59715e-19 $X=1.675 $Y=1.402 $X2=0.24 $Y2=0
cc_99 N_A_30_107#_c_129_n N_VPWR_c_184_n 0.00971499f $X=1.2 $Y=1.99 $X2=0.24
+ $Y2=0
cc_100 N_A_30_107#_c_146_n N_VPWR_c_184_n 0.0137383f $X=0.885 $Y=1.99 $X2=0.24
+ $Y2=0
cc_101 N_A_30_107#_c_130_n N_VPWR_c_184_n 0.0182289f $X=1.285 $Y=2.425 $X2=0.24
+ $Y2=0
cc_102 N_A_30_107#_M1000_g N_VPWR_c_187_n 0.10669f $X=2.675 $Y=2.965 $X2=0 $Y2=0
cc_103 N_A_30_107#_c_130_n N_VPWR_c_187_n 0.0182289f $X=1.285 $Y=2.425 $X2=0
+ $Y2=0
cc_104 N_A_30_107#_c_131_n N_VPWR_c_187_n 0.0634128f $X=2.445 $Y=1.99 $X2=0
+ $Y2=0
cc_105 N_A_30_107#_c_163_n N_VPWR_c_187_n 0.0252329f $X=2.61 $Y=1.89 $X2=0 $Y2=0
cc_106 N_A_30_107#_M1000_g N_VPWR_c_190_n 0.00915578f $X=2.675 $Y=2.965 $X2=0
+ $Y2=0
cc_107 N_A_30_107#_M1000_g N_X_c_209_n 0.00932666f $X=2.675 $Y=2.965 $X2=0 $Y2=0
cc_108 N_A_30_107#_M1002_g N_X_c_209_n 0.0345604f $X=2.695 $Y=0.91 $X2=0 $Y2=0
cc_109 N_A_30_107#_c_163_n N_X_c_209_n 0.0237234f $X=2.61 $Y=1.89 $X2=0 $Y2=0
cc_110 N_A_30_107#_M1002_g N_VGND_c_225_n 0.0445357f $X=2.695 $Y=0.91 $X2=0
+ $Y2=0
cc_111 N_A_30_107#_c_131_n N_VGND_c_225_n 0.0265726f $X=2.445 $Y=1.99 $X2=0
+ $Y2=0
cc_112 N_A_30_107#_c_163_n N_VGND_c_225_n 0.00716041f $X=2.61 $Y=1.89 $X2=0
+ $Y2=0
cc_113 N_A_30_107#_c_125_n N_VGND_c_225_n 7.34328e-19 $X=2.61 $Y=1.89 $X2=0
+ $Y2=0
cc_114 N_A_30_107#_M1005_s N_VGND_c_227_n 2.95251e-19 $X=0.15 $Y=0.535 $X2=0.24
+ $Y2=0
cc_115 N_A_30_107#_M1002_g N_VGND_c_227_n 0.0210736f $X=2.695 $Y=0.91 $X2=0.24
+ $Y2=0
cc_116 N_A_30_107#_c_121_n N_VGND_c_227_n 0.0200915f $X=0.275 $Y=0.745 $X2=0.24
+ $Y2=0
cc_117 N_A_30_107#_c_123_n N_VGND_c_227_n 0.0219126f $X=0.715 $Y=0.91 $X2=0.24
+ $Y2=0
cc_118 N_VPWR_c_190_n N_X_M1000_d 0.00221032f $X=2.715 $Y=3.59 $X2=0 $Y2=0
cc_119 N_VPWR_c_187_n N_X_c_209_n 0.0631064f $X=2.18 $Y=2.34 $X2=1.68 $Y2=4.07
cc_120 N_VPWR_c_190_n N_X_c_209_n 0.0375086f $X=2.715 $Y=3.59 $X2=1.68 $Y2=4.07
cc_121 N_X_c_209_n N_VGND_c_225_n 0.0204194f $X=3.085 $Y=0.68 $X2=0 $Y2=0
cc_122 N_X_M1002_d N_VGND_c_227_n 0.00137624f $X=2.945 $Y=0.535 $X2=0.24 $Y2=0
cc_123 N_X_c_209_n N_VGND_c_227_n 0.0293415f $X=3.085 $Y=0.68 $X2=0.24 $Y2=0
cc_124 A_183_107# N_VGND_c_227_n 0.00681585f $X=0.915 $Y=0.535 $X2=0 $Y2=0
