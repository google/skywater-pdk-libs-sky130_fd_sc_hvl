* File: sky130_fd_sc_hvl__probec_p_8.spice
* Created: Wed Sep  2 09:09:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__probec_p_8.pex.spice"
.subckt sky130_fd_sc_hvl__probec_p_8  VNB VPB A VPWR VGND X
* 
* X	X
* VGND	VGND
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_A_45_443#_M1003_d N_A_M1003_g N_VGND_M1003_s N_VNB_M1003_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.2025 PD=2.07 PS=1.29 NRD=3.0324 NRS=6.0762 M=1 R=1.5
+ SA=250000 SB=250008 A=0.375 P=2.5 MULT=1
MM1008 N_A_45_443#_M1008_d N_A_M1008_g N_VGND_M1003_s N_VNB_M1003_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.2025 PD=1.03 PS=1.29 NRD=0 NRS=33.4362 M=1 R=1.5
+ SA=250001 SB=250007 A=0.375 P=2.5 MULT=1
MM1015 N_A_45_443#_M1008_d N_A_M1015_g N_VGND_M1015_s N_VNB_M1003_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250002
+ SB=250006 A=0.375 P=2.5 MULT=1
MM1001 N_noxref_6_M1001_d N_A_45_443#_M1001_g N_VGND_M1015_s N_VNB_M1003_b NHV
+ L=0.5 W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250003
+ SB=250005 A=0.375 P=2.5 MULT=1
MM1002 N_noxref_6_M1001_d N_A_45_443#_M1002_g N_VGND_M1002_s N_VNB_M1003_b NHV
+ L=0.5 W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250003
+ SB=250005 A=0.375 P=2.5 MULT=1
MM1009 N_noxref_6_M1009_d N_A_45_443#_M1009_g N_VGND_M1002_s N_VNB_M1003_b NHV
+ L=0.5 W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250004
+ SB=250004 A=0.375 P=2.5 MULT=1
MM1013 N_noxref_6_M1009_d N_A_45_443#_M1013_g N_VGND_M1013_s N_VNB_M1003_b NHV
+ L=0.5 W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250005
+ SB=250003 A=0.375 P=2.5 MULT=1
MM1014 N_noxref_6_M1014_d N_A_45_443#_M1014_g N_VGND_M1013_s N_VNB_M1003_b NHV
+ L=0.5 W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250006
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1018 N_noxref_6_M1014_d N_A_45_443#_M1018_g N_VGND_M1018_s N_VNB_M1003_b NHV
+ L=0.5 W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250007
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1020 N_noxref_6_M1020_d N_A_45_443#_M1020_g N_VGND_M1018_s N_VNB_M1003_b NHV
+ L=0.5 W=0.75 AD=0.105 AS=0.105 PD=1.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250007
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1021 N_noxref_6_M1020_d N_A_45_443#_M1021_g N_VGND_M1021_s N_VNB_M1003_b NHV
+ L=0.5 W=0.75 AD=0.105 AS=0.21375 PD=1.03 PS=2.07 NRD=0 NRS=3.0324 M=1 R=1.5
+ SA=250008 SB=250000 A=0.375 P=2.5 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_45_443#_M1006_s N_VPB_M1006_b PHV L=0.5
+ W=1.5 AD=0.42 AS=0.4275 PD=2.06 PS=3.57 NRD=0 NRS=2.5403 M=1 R=3 SA=250000
+ SB=250008 A=0.75 P=4 MULT=1
MM1007 N_VPWR_M1006_d N_A_M1007_g N_A_45_443#_M1007_s N_VPB_M1006_b PHV L=0.5
+ W=1.5 AD=0.42 AS=0.21 PD=2.06 PS=1.78 NRD=35.6406 NRS=0 M=1 R=3 SA=250001
+ SB=250007 A=0.75 P=4 MULT=1
MM1019 N_VPWR_M1019_d N_A_M1019_g N_A_45_443#_M1007_s N_VPB_M1006_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002 SB=250006
+ A=0.75 P=4 MULT=1
MM1000 N_noxref_6_M1000_d N_A_45_443#_M1000_g N_VPWR_M1019_d N_VPB_M1006_b PHV
+ L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250003
+ SB=250005 A=0.75 P=4 MULT=1
MM1004 N_noxref_6_M1000_d N_A_45_443#_M1004_g N_VPWR_M1004_s N_VPB_M1006_b PHV
+ L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250003
+ SB=250005 A=0.75 P=4 MULT=1
MM1005 N_noxref_6_M1005_d N_A_45_443#_M1005_g N_VPWR_M1004_s N_VPB_M1006_b PHV
+ L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250004
+ SB=250004 A=0.75 P=4 MULT=1
MM1010 N_noxref_6_M1005_d N_A_45_443#_M1010_g N_VPWR_M1010_s N_VPB_M1006_b PHV
+ L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250005
+ SB=250003 A=0.75 P=4 MULT=1
MM1011 N_noxref_6_M1011_d N_A_45_443#_M1011_g N_VPWR_M1010_s N_VPB_M1006_b PHV
+ L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250006
+ SB=250002 A=0.75 P=4 MULT=1
MM1012 N_noxref_6_M1011_d N_A_45_443#_M1012_g N_VPWR_M1012_s N_VPB_M1006_b PHV
+ L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250007
+ SB=250002 A=0.75 P=4 MULT=1
MM1016 N_noxref_6_M1016_d N_A_45_443#_M1016_g N_VPWR_M1012_s N_VPB_M1006_b PHV
+ L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250007
+ SB=250001 A=0.75 P=4 MULT=1
MM1017 N_noxref_6_M1016_d N_A_45_443#_M1017_g N_VPWR_M1017_s N_VPB_M1006_b PHV
+ L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 M=1 R=3 SA=250008
+ SB=250000 A=0.75 P=4 MULT=1
DX22_noxref N_VNB_M1003_b N_VPB_M1006_b NWDIODE A=26.676 P=25.72
R23_noxref N_X_R23_noxref_pos N_noxref_6_R23_noxref_neg SHORT 0.01 M=1
*
.include "sky130_fd_sc_hvl__probec_p_8.pxi.spice"
*
.ends
*
*
