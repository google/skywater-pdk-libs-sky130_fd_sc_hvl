* File: sky130_fd_sc_hvl__inv_2.pxi.spice
* Created: Fri Aug 28 09:36:06 2020
* 
x_PM_SKY130_FD_SC_HVL__INV_2%VNB N_VNB_M1001_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__INV_2%VNB
x_PM_SKY130_FD_SC_HVL__INV_2%VPB N_VPB_M1000_b VPB N_VPB_c_17_p VPB
+ PM_SKY130_FD_SC_HVL__INV_2%VPB
x_PM_SKY130_FD_SC_HVL__INV_2%A N_A_M1001_g N_A_M1000_g N_A_M1003_g N_A_M1002_g A
+ A N_A_c_38_n N_A_c_39_n PM_SKY130_FD_SC_HVL__INV_2%A
x_PM_SKY130_FD_SC_HVL__INV_2%VPWR N_VPWR_M1000_d N_VPWR_M1002_d VPWR
+ N_VPWR_c_74_n N_VPWR_c_77_n N_VPWR_c_80_n PM_SKY130_FD_SC_HVL__INV_2%VPWR
x_PM_SKY130_FD_SC_HVL__INV_2%Y N_Y_M1001_d N_Y_M1000_s N_Y_c_97_n Y Y Y
+ N_Y_c_95_n Y PM_SKY130_FD_SC_HVL__INV_2%Y
x_PM_SKY130_FD_SC_HVL__INV_2%VGND N_VGND_M1001_s N_VGND_M1003_s VGND
+ N_VGND_c_122_n N_VGND_c_124_n N_VGND_c_126_n PM_SKY130_FD_SC_HVL__INV_2%VGND
cc_1 N_VNB_M1001_b N_A_M1001_g 0.0474057f $X=-0.33 $Y=-0.265 $X2=0.935 $Y2=0.955
cc_2 N_VNB_c_2_p N_A_M1001_g 7.33495e-19 $X=0.24 $Y=0 $X2=0.935 $Y2=0.955
cc_3 N_VNB_M1001_b N_A_M1003_g 0.0528627f $X=-0.33 $Y=-0.265 $X2=1.715 $Y2=0.955
cc_4 N_VNB_c_2_p N_A_M1003_g 0.00220932f $X=0.24 $Y=0 $X2=1.715 $Y2=0.955
cc_5 N_VNB_M1001_b N_A_c_38_n 0.0202641f $X=-0.33 $Y=-0.265 $X2=0.905 $Y2=1.715
cc_6 N_VNB_M1001_b N_A_c_39_n 0.122712f $X=-0.33 $Y=-0.265 $X2=1.715 $Y2=1.772
cc_7 N_VNB_M1001_b N_Y_c_95_n 0.0189319f $X=-0.33 $Y=-0.265 $X2=0.24 $Y2=1.715
cc_8 N_VNB_c_2_p N_Y_c_95_n 0.00201821f $X=0.24 $Y=0 $X2=0.24 $Y2=1.715
cc_9 N_VNB_M1001_b N_VGND_c_122_n 0.0980976f $X=-0.33 $Y=-0.265 $X2=1.715
+ $Y2=0.955
cc_10 N_VNB_c_2_p N_VGND_c_122_n 0.00263373f $X=0.24 $Y=0 $X2=1.715 $Y2=0.955
cc_11 N_VNB_M1001_b N_VGND_c_124_n 0.067735f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_12 N_VNB_c_2_p N_VGND_c_124_n 9.30887e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_13 N_VNB_M1001_b N_VGND_c_126_n 0.0609797f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_14 N_VNB_c_2_p N_VGND_c_126_n 0.256675f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_15 N_VPB_M1000_b N_A_M1000_g 0.0412236f $X=-0.33 $Y=1.885 $X2=0.935 $Y2=2.965
cc_16 VPB N_A_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.935 $Y2=2.965
cc_17 N_VPB_c_17_p N_A_M1000_g 0.0152133f $X=2.16 $Y=4.07 $X2=0.935 $Y2=2.965
cc_18 N_VPB_M1000_b N_A_M1002_g 0.0407066f $X=-0.33 $Y=1.885 $X2=1.715 $Y2=2.965
cc_19 VPB N_A_M1002_g 0.00970178f $X=0 $Y=3.955 $X2=1.715 $Y2=2.965
cc_20 N_VPB_c_17_p N_A_M1002_g 0.0160007f $X=2.16 $Y=4.07 $X2=1.715 $Y2=2.965
cc_21 N_VPB_M1000_b N_A_c_39_n 0.0521325f $X=-0.33 $Y=1.885 $X2=1.715 $Y2=1.772
cc_22 N_VPB_M1000_b N_VPWR_c_74_n 0.0815209f $X=-0.33 $Y=1.885 $X2=1.715
+ $Y2=0.955
cc_23 VPB N_VPWR_c_74_n 0.00355415f $X=0 $Y=3.955 $X2=1.715 $Y2=0.955
cc_24 N_VPB_c_17_p N_VPWR_c_74_n 0.0486145f $X=2.16 $Y=4.07 $X2=1.715 $Y2=0.955
cc_25 N_VPB_M1000_b N_VPWR_c_77_n 0.0699853f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_26 VPB N_VPWR_c_77_n 0.00229469f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_27 N_VPB_c_17_p N_VPWR_c_77_n 0.0299474f $X=2.16 $Y=4.07 $X2=0 $Y2=0
cc_28 N_VPB_M1000_b N_VPWR_c_80_n 0.0447014f $X=-0.33 $Y=1.885 $X2=1.715
+ $Y2=1.772
cc_29 VPB N_VPWR_c_80_n 0.254901f $X=0 $Y=3.955 $X2=1.715 $Y2=1.772
cc_30 N_VPB_c_17_p N_VPWR_c_80_n 0.0107625f $X=2.16 $Y=4.07 $X2=1.715 $Y2=1.772
cc_31 N_VPB_M1000_b N_Y_c_97_n 0.00229403f $X=-0.33 $Y=1.885 $X2=1.715 $Y2=1.46
cc_32 VPB N_Y_c_97_n 8.01732e-19 $X=0 $Y=3.955 $X2=1.715 $Y2=1.46
cc_33 N_VPB_c_17_p N_Y_c_97_n 0.0130099f $X=2.16 $Y=4.07 $X2=1.715 $Y2=1.46
cc_34 N_A_M1000_g N_VPWR_c_74_n 0.0800526f $X=0.935 $Y=2.965 $X2=0.24 $Y2=0
cc_35 N_A_M1002_g N_VPWR_c_74_n 6.71148e-19 $X=1.715 $Y=2.965 $X2=0.24 $Y2=0
cc_36 N_A_c_38_n N_VPWR_c_74_n 0.051693f $X=0.905 $Y=1.715 $X2=0.24 $Y2=0
cc_37 N_A_c_39_n N_VPWR_c_74_n 0.00618002f $X=1.715 $Y=1.772 $X2=0.24 $Y2=0
cc_38 N_A_M1002_g N_VPWR_c_77_n 0.0791104f $X=1.715 $Y=2.965 $X2=0 $Y2=0
cc_39 N_A_M1000_g N_VPWR_c_80_n 0.00830187f $X=0.935 $Y=2.965 $X2=1.2 $Y2=0.058
cc_40 N_A_M1002_g N_VPWR_c_80_n 0.0110007f $X=1.715 $Y=2.965 $X2=1.2 $Y2=0.058
cc_41 N_A_M1000_g N_Y_c_97_n 0.00383933f $X=0.935 $Y=2.965 $X2=0 $Y2=0
cc_42 N_A_M1002_g N_Y_c_97_n 0.0311988f $X=1.715 $Y=2.965 $X2=0 $Y2=0
cc_43 N_A_c_38_n N_Y_c_97_n 0.00774718f $X=0.905 $Y=1.715 $X2=0 $Y2=0
cc_44 N_A_c_39_n N_Y_c_97_n 0.0343483f $X=1.715 $Y=1.772 $X2=0 $Y2=0
cc_45 N_A_M1001_g Y 5.17969e-19 $X=0.935 $Y=0.955 $X2=0 $Y2=0
cc_46 N_A_M1003_g Y 0.00672922f $X=1.715 $Y=0.955 $X2=0 $Y2=0
cc_47 N_A_c_38_n Y 0.00191561f $X=0.905 $Y=1.715 $X2=0 $Y2=0
cc_48 N_A_c_39_n Y 0.0155831f $X=1.715 $Y=1.772 $X2=0 $Y2=0
cc_49 N_A_c_38_n Y 0.0140049f $X=0.905 $Y=1.715 $X2=0 $Y2=0
cc_50 N_A_c_39_n Y 0.0355066f $X=1.715 $Y=1.772 $X2=0 $Y2=0
cc_51 N_A_M1001_g N_Y_c_95_n 0.00145816f $X=0.935 $Y=0.955 $X2=0 $Y2=0
cc_52 N_A_M1003_g N_Y_c_95_n 0.0397835f $X=1.715 $Y=0.955 $X2=0 $Y2=0
cc_53 N_A_c_39_n N_Y_c_95_n 0.00304639f $X=1.715 $Y=1.772 $X2=0 $Y2=0
cc_54 N_A_M1001_g N_VGND_c_122_n 0.0547661f $X=0.935 $Y=0.955 $X2=0.24 $Y2=0
cc_55 N_A_M1003_g N_VGND_c_122_n 0.00102944f $X=1.715 $Y=0.955 $X2=0.24 $Y2=0
cc_56 N_A_c_38_n N_VGND_c_122_n 0.071843f $X=0.905 $Y=1.715 $X2=0.24 $Y2=0
cc_57 N_A_c_39_n N_VGND_c_122_n 0.00660654f $X=1.715 $Y=1.772 $X2=0.24 $Y2=0
cc_58 N_A_M1003_g N_VGND_c_124_n 0.00870988f $X=1.715 $Y=0.955 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_VGND_c_126_n 0.0100782f $X=0.935 $Y=0.955 $X2=0 $Y2=0
cc_60 N_A_M1003_g N_VGND_c_126_n 0.015568f $X=1.715 $Y=0.955 $X2=0 $Y2=0
cc_61 N_VPWR_c_80_n N_Y_M1000_s 0.00221032f $X=2.155 $Y=3.59 $X2=0 $Y2=0
cc_62 N_VPWR_c_74_n N_Y_c_97_n 0.0677867f $X=0.545 $Y=2.34 $X2=0.24 $Y2=4.07
cc_63 N_VPWR_c_77_n N_Y_c_97_n 0.107316f $X=2.105 $Y=2.34 $X2=0.24 $Y2=4.07
cc_64 N_VPWR_c_80_n N_Y_c_97_n 0.0306945f $X=2.155 $Y=3.59 $X2=0.24 $Y2=4.07
cc_65 N_VPWR_c_77_n Y 0.00437535f $X=2.105 $Y=2.34 $X2=2.16 $Y2=4.07
cc_66 N_Y_c_95_n N_VGND_c_122_n 0.0363049f $X=1.325 $Y=0.705 $X2=0.24 $Y2=0
cc_67 N_Y_c_95_n N_VGND_c_124_n 0.0347041f $X=1.325 $Y=0.705 $X2=0 $Y2=0
cc_68 N_Y_M1001_d N_VGND_c_126_n 5.42154e-19 $X=1.185 $Y=0.58 $X2=0 $Y2=0
cc_69 N_Y_c_95_n N_VGND_c_126_n 0.0515038f $X=1.325 $Y=0.705 $X2=0 $Y2=0
