* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_271_107# A2 VGND VNB nhv w=750000u l=500000u
+  ad=1.575e+11p pd=1.92e+06u as=4.125e+11p ps=4.1e+06u
M1001 Y B1 a_56_443# VPB phv w=1.5e+06u l=500000u
+  ad=5.475e+11p pd=3.73e+06u as=8.475e+11p ps=7.13e+06u
M1002 VGND B1 Y VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=2.85e+11p ps=2.26e+06u
M1003 VPWR A2 a_56_443# VPB phv w=1.5e+06u l=500000u
+  ad=7.5e+11p pd=4e+06u as=0p ps=0u
M1004 Y A1 a_271_107# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_56_443# A1 VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
