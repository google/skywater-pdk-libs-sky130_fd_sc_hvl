* File: sky130_fd_sc_hvl__sdfrtp_1.pxi.spice
* Created: Wed Sep  2 09:10:03 2020
* 
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%VNB N_VNB_M1002_b VNB N_VNB_c_8_p
+ PM_SKY130_FD_SC_HVL__SDFRTP_1%VNB
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%VPB N_VPB_M1008_b VPB N_VPB_c_134_p
+ PM_SKY130_FD_SC_HVL__SDFRTP_1%VPB
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%A_116_451# N_A_116_451#_M1012_d
+ N_A_116_451#_M1014_d N_A_116_451#_c_347_n N_A_116_451#_M1008_g
+ N_A_116_451#_c_339_n N_A_116_451#_M1038_g N_A_116_451#_c_351_n
+ N_A_116_451#_c_352_n N_A_116_451#_c_452_p N_A_116_451#_c_341_n
+ N_A_116_451#_c_342_n N_A_116_451#_c_343_n N_A_116_451#_c_354_n
+ N_A_116_451#_c_355_n N_A_116_451#_c_356_n N_A_116_451#_c_357_n
+ N_A_116_451#_c_344_n N_A_116_451#_c_358_n N_A_116_451#_c_359_n
+ N_A_116_451#_c_360_n N_A_116_451#_c_361_n N_A_116_451#_c_345_n
+ N_A_116_451#_c_372_p N_A_116_451#_c_393_p
+ PM_SKY130_FD_SC_HVL__SDFRTP_1%A_116_451#
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%SCD N_SCD_c_500_n N_SCD_M1002_g N_SCD_c_501_n
+ N_SCD_M1011_g N_SCD_c_502_n N_SCD_c_503_n SCD SCD N_SCD_c_504_n
+ PM_SKY130_FD_SC_HVL__SDFRTP_1%SCD
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%SCE N_SCE_M1016_g N_SCE_c_560_n N_SCE_M1035_g
+ N_SCE_M1014_g N_SCE_c_567_n N_SCE_c_552_n N_SCE_c_553_n N_SCE_c_568_n
+ N_SCE_c_554_n N_SCE_c_555_n SCE SCE SCE SCE SCE N_SCE_M1012_g N_SCE_c_559_n
+ PM_SKY130_FD_SC_HVL__SDFRTP_1%SCE
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%D N_D_c_681_n N_D_M1004_g D D N_D_c_683_n
+ N_D_M1037_g PM_SKY130_FD_SC_HVL__SDFRTP_1%D
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%A_1212_471# N_A_1212_471#_M1032_s
+ N_A_1212_471#_M1020_s N_A_1212_471#_c_737_n N_A_1212_471#_M1030_g
+ N_A_1212_471#_c_738_n N_A_1212_471#_c_750_n N_A_1212_471#_c_739_n
+ N_A_1212_471#_c_741_n N_A_1212_471#_c_753_n N_A_1212_471#_c_756_n
+ N_A_1212_471#_c_743_n N_A_1212_471#_c_744_n N_A_1212_471#_c_786_p
+ N_A_1212_471#_c_759_n N_A_1212_471#_c_788_p N_A_1212_471#_c_745_n
+ N_A_1212_471#_c_836_p N_A_1212_471#_c_760_n N_A_1212_471#_c_763_n
+ N_A_1212_471#_c_766_n N_A_1212_471#_c_767_n N_A_1212_471#_c_795_p
+ N_A_1212_471#_c_768_n N_A_1212_471#_c_798_p N_A_1212_471#_c_769_n
+ N_A_1212_471#_c_800_p N_A_1212_471#_c_770_n N_A_1212_471#_c_887_p
+ N_A_1212_471#_c_746_n N_A_1212_471#_c_771_n N_A_1212_471#_c_772_n
+ N_A_1212_471#_c_802_p N_A_1212_471#_M1026_g N_A_1212_471#_M1001_g
+ N_A_1212_471#_M1023_g PM_SKY130_FD_SC_HVL__SDFRTP_1%A_1212_471#
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%A_1212_100# N_A_1212_100#_M1033_s
+ N_A_1212_100#_M1018_d N_A_1212_100#_M1022_g N_A_1212_100#_c_1003_n
+ N_A_1212_100#_c_1004_n N_A_1212_100#_c_1005_n N_A_1212_100#_M1003_g
+ N_A_1212_100#_c_977_n N_A_1212_100#_M1032_g N_A_1212_100#_c_978_n
+ N_A_1212_100#_M1020_g N_A_1212_100#_c_1013_n N_A_1212_100#_M1036_g
+ N_A_1212_100#_c_979_n N_A_1212_100#_M1000_g N_A_1212_100#_c_1062_n
+ N_A_1212_100#_c_981_n N_A_1212_100#_c_982_n N_A_1212_100#_c_983_n
+ N_A_1212_100#_c_1070_n N_A_1212_100#_c_984_n N_A_1212_100#_c_986_n
+ N_A_1212_100#_c_988_n N_A_1212_100#_c_989_n N_A_1212_100#_c_990_n
+ N_A_1212_100#_c_991_n N_A_1212_100#_c_992_n N_A_1212_100#_c_994_n
+ N_A_1212_100#_c_996_n N_A_1212_100#_c_997_n N_A_1212_100#_c_998_n
+ N_A_1212_100#_c_1018_n N_A_1212_100#_c_1021_n N_A_1212_100#_c_1022_n
+ N_A_1212_100#_c_999_n N_A_1212_100#_c_1023_n N_A_1212_100#_c_1000_n
+ N_A_1212_100#_c_1001_n PM_SKY130_FD_SC_HVL__SDFRTP_1%A_1212_100#
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%A_1510_100# N_A_1510_100#_M1007_d
+ N_A_1510_100#_M1009_d N_A_1510_100#_M1010_g N_A_1510_100#_M1015_g
+ N_A_1510_100#_c_1246_n N_A_1510_100#_c_1267_n N_A_1510_100#_c_1247_n
+ N_A_1510_100#_c_1253_n N_A_1510_100#_c_1292_n N_A_1510_100#_c_1248_n
+ N_A_1510_100#_c_1274_n N_A_1510_100#_c_1255_n N_A_1510_100#_c_1256_n
+ PM_SKY130_FD_SC_HVL__SDFRTP_1%A_1510_100#
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%RESET_B N_RESET_B_M1019_g N_RESET_B_M1024_g
+ N_RESET_B_c_1352_n N_RESET_B_c_1353_n N_RESET_B_M1013_g N_RESET_B_c_1364_n
+ N_RESET_B_c_1356_n N_RESET_B_c_1357_n RESET_B N_RESET_B_c_1365_n
+ N_RESET_B_c_1366_n N_RESET_B_c_1367_n N_RESET_B_c_1368_n N_RESET_B_c_1369_n
+ N_RESET_B_c_1370_n N_RESET_B_c_1358_n N_RESET_B_c_1387_n N_RESET_B_c_1359_n
+ N_RESET_B_c_1375_n N_RESET_B_M1027_g N_RESET_B_M1025_g N_RESET_B_c_1457_n
+ N_RESET_B_M1006_g PM_SKY130_FD_SC_HVL__SDFRTP_1%RESET_B
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%A_1312_126# N_A_1312_126#_M1022_d
+ N_A_1312_126#_M1026_d N_A_1312_126#_M1027_d N_A_1312_126#_M1007_g
+ N_A_1312_126#_c_1562_n N_A_1312_126#_M1009_g N_A_1312_126#_c_1563_n
+ N_A_1312_126#_c_1589_n N_A_1312_126#_c_1569_n N_A_1312_126#_c_1570_n
+ N_A_1312_126#_c_1571_n N_A_1312_126#_c_1572_n N_A_1312_126#_c_1573_n
+ N_A_1312_126#_c_1564_n N_A_1312_126#_c_1574_n N_A_1312_126#_c_1575_n
+ N_A_1312_126#_c_1611_n PM_SKY130_FD_SC_HVL__SDFRTP_1%A_1312_126#
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%A_2616_417# N_A_2616_417#_M1031_d
+ N_A_2616_417#_M1006_d N_A_2616_417#_M1039_g N_A_2616_417#_c_1693_n
+ N_A_2616_417#_c_1694_n N_A_2616_417#_c_1695_n N_A_2616_417#_c_1751_p
+ N_A_2616_417#_c_1696_n N_A_2616_417#_c_1689_n N_A_2616_417#_c_1707_n
+ N_A_2616_417#_c_1708_n N_A_2616_417#_c_1698_n N_A_2616_417#_c_1690_n
+ N_A_2616_417#_M1021_g PM_SKY130_FD_SC_HVL__SDFRTP_1%A_2616_417#
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%A_2360_115# N_A_2360_115#_M1030_d
+ N_A_2360_115#_M1036_d N_A_2360_115#_M1031_g N_A_2360_115#_M1028_g
+ N_A_2360_115#_M1029_g N_A_2360_115#_M1005_g N_A_2360_115#_c_1783_n
+ N_A_2360_115#_c_1784_n N_A_2360_115#_c_1785_n N_A_2360_115#_c_1786_n
+ N_A_2360_115#_c_1795_n N_A_2360_115#_c_1796_n N_A_2360_115#_c_1797_n
+ N_A_2360_115#_c_1798_n N_A_2360_115#_c_1799_n N_A_2360_115#_c_1800_n
+ N_A_2360_115#_c_1801_n N_A_2360_115#_c_1802_n N_A_2360_115#_c_1805_n
+ N_A_2360_115#_c_1902_n N_A_2360_115#_c_1905_n N_A_2360_115#_c_1808_n
+ N_A_2360_115#_c_1787_n N_A_2360_115#_c_1788_n N_A_2360_115#_c_1789_n
+ PM_SKY130_FD_SC_HVL__SDFRTP_1%A_2360_115#
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%CLK N_CLK_c_1958_n N_CLK_M1033_g CLK
+ N_CLK_c_1960_n N_CLK_c_1964_n N_CLK_M1018_g PM_SKY130_FD_SC_HVL__SDFRTP_1%CLK
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%A_3417_443# N_A_3417_443#_M1005_s
+ N_A_3417_443#_M1029_s N_A_3417_443#_M1017_g N_A_3417_443#_M1034_g
+ N_A_3417_443#_c_1997_n N_A_3417_443#_c_1998_n N_A_3417_443#_c_1999_n
+ N_A_3417_443#_c_2000_n N_A_3417_443#_c_2005_n N_A_3417_443#_c_2012_n
+ N_A_3417_443#_c_2014_n PM_SKY130_FD_SC_HVL__SDFRTP_1%A_3417_443#
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%A_65_649# N_A_65_649#_M1016_d
+ N_A_65_649#_M1022_s N_A_65_649#_M1008_s N_A_65_649#_M1037_d
+ N_A_65_649#_M1026_s N_A_65_649#_c_2046_n N_A_65_649#_c_2055_n
+ N_A_65_649#_c_2047_n N_A_65_649#_c_2048_n N_A_65_649#_c_2058_n
+ N_A_65_649#_c_2091_n N_A_65_649#_c_2122_n N_A_65_649#_c_2049_n
+ N_A_65_649#_c_2127_n N_A_65_649#_c_2059_n N_A_65_649#_c_2062_n
+ N_A_65_649#_c_2065_n N_A_65_649#_c_2066_n N_A_65_649#_c_2067_n
+ N_A_65_649#_c_2099_n N_A_65_649#_c_2068_n N_A_65_649#_c_2071_n
+ N_A_65_649#_c_2050_n N_A_65_649#_c_2074_n N_A_65_649#_c_2075_n
+ N_A_65_649#_c_2076_n N_A_65_649#_c_2052_n N_A_65_649#_c_2053_n
+ PM_SKY130_FD_SC_HVL__SDFRTP_1%A_65_649#
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%VPWR N_VPWR_M1011_d N_VPWR_M1019_d
+ N_VPWR_M1015_d N_VPWR_M1020_d N_VPWR_M1039_d N_VPWR_M1028_d N_VPWR_M1029_d
+ VPWR N_VPWR_c_2199_n N_VPWR_c_2202_n N_VPWR_c_2205_n N_VPWR_c_2208_n
+ N_VPWR_c_2211_n N_VPWR_c_2214_n N_VPWR_c_2217_n N_VPWR_c_2220_n
+ PM_SKY130_FD_SC_HVL__SDFRTP_1%VPWR
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%Q N_Q_M1034_d N_Q_M1017_d Q Q Q Q Q Q Q
+ N_Q_c_2350_n PM_SKY130_FD_SC_HVL__SDFRTP_1%Q
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%noxref_23 N_noxref_23_M1002_s
+ N_noxref_23_M1004_d N_noxref_23_c_2364_n N_noxref_23_c_2365_n
+ N_noxref_23_c_2367_n N_noxref_23_c_2369_n
+ PM_SKY130_FD_SC_HVL__SDFRTP_1%noxref_23
x_PM_SKY130_FD_SC_HVL__SDFRTP_1%VGND N_VGND_M1024_d N_VGND_M1013_d
+ N_VGND_M1032_d N_VGND_M1021_d N_VGND_M1033_d N_VGND_M1005_d VGND
+ N_VGND_c_2396_n N_VGND_c_2398_n N_VGND_c_2400_n N_VGND_c_2402_n
+ N_VGND_c_2404_n N_VGND_c_2406_n N_VGND_c_2408_n
+ PM_SKY130_FD_SC_HVL__SDFRTP_1%VGND
cc_1 N_VNB_M1002_b N_A_116_451#_c_339_n 0.0492856f $X=-0.33 $Y=-0.265 $X2=2.71
+ $Y2=1.315
cc_2 N_VNB_M1002_b N_A_116_451#_M1038_g 0.0486686f $X=-0.33 $Y=-0.265 $X2=2.71
+ $Y2=0.84
cc_3 N_VNB_M1002_b N_A_116_451#_c_341_n 0.00490686f $X=-0.33 $Y=-0.265 $X2=1.73
+ $Y2=2.755
cc_4 N_VNB_M1002_b N_A_116_451#_c_342_n 0.00608073f $X=-0.33 $Y=-0.265 $X2=2.48
+ $Y2=1.18
cc_5 N_VNB_M1002_b N_A_116_451#_c_343_n 0.00137292f $X=-0.33 $Y=-0.265 $X2=1.815
+ $Y2=1.18
cc_6 N_VNB_M1002_b N_A_116_451#_c_344_n 0.0223935f $X=-0.33 $Y=-0.265 $X2=5.285
+ $Y2=1.26
cc_7 N_VNB_M1002_b N_A_116_451#_c_345_n 0.0171391f $X=-0.33 $Y=-0.265 $X2=5.37
+ $Y2=0.84
cc_8 N_VNB_c_8_p N_A_116_451#_c_345_n 5.64934e-19 $X=0.24 $Y=0 $X2=5.37 $Y2=0.84
cc_9 N_VNB_M1002_b N_SCD_c_500_n 0.0427537f $X=-0.33 $Y=-0.265 $X2=5.23 $Y2=0.63
cc_10 N_VNB_M1002_b N_SCD_c_501_n 0.0354654f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_11 N_VNB_M1002_b N_SCD_c_502_n 0.109193f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_12 N_VNB_M1002_b N_SCD_c_503_n 0.028355f $X=-0.33 $Y=-0.265 $X2=2.71
+ $Y2=1.315
cc_13 N_VNB_M1002_b N_SCD_c_504_n 0.0133586f $X=-0.33 $Y=-0.265 $X2=2.48
+ $Y2=1.18
cc_14 N_VNB_M1002_b N_SCE_M1016_g 0.0448137f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_15 N_VNB_M1002_b N_SCE_c_552_n 0.00256375f $X=-0.33 $Y=-0.265 $X2=0.895
+ $Y2=2.42
cc_16 N_VNB_M1002_b N_SCE_c_553_n 0.060573f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_17 N_VNB_M1002_b N_SCE_c_554_n 0.00619829f $X=-0.33 $Y=-0.265 $X2=2.56
+ $Y2=2.84
cc_18 N_VNB_M1002_b N_SCE_c_555_n 0.00249711f $X=-0.33 $Y=-0.265 $X2=2.645
+ $Y2=2.48
cc_19 N_VNB_M1002_b SCE 0.00617497f $X=-0.33 $Y=-0.265 $X2=2.645 $Y2=2.755
cc_20 N_VNB_M1002_b SCE 0.012354f $X=-0.33 $Y=-0.265 $X2=2.81 $Y2=1.26
cc_21 N_VNB_M1002_b N_SCE_M1012_g 0.101921f $X=-0.33 $Y=-0.265 $X2=5.41 $Y2=0.84
cc_22 N_VNB_M1002_b N_SCE_c_559_n 0.0208142f $X=-0.33 $Y=-0.265 $X2=2.645
+ $Y2=1.57
cc_23 N_VNB_M1002_b N_D_M1004_g 0.0995061f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_24 N_VNB_M1002_b N_A_1212_471#_c_737_n 0.0811343f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=3.115
cc_25 N_VNB_M1002_b N_A_1212_471#_c_738_n 0.00163893f $X=-0.33 $Y=-0.265
+ $X2=2.71 $Y2=0.84
cc_26 N_VNB_M1002_b N_A_1212_471#_c_739_n 0.064348f $X=-0.33 $Y=-0.265 $X2=0.895
+ $Y2=2.755
cc_27 N_VNB_c_8_p N_A_1212_471#_c_739_n 0.00402054f $X=0.24 $Y=0 $X2=0.895
+ $Y2=2.755
cc_28 N_VNB_M1002_b N_A_1212_471#_c_741_n 0.0126949f $X=-0.33 $Y=-0.265
+ $X2=0.895 $Y2=2.42
cc_29 N_VNB_c_8_p N_A_1212_471#_c_741_n 8.18031e-19 $X=0.24 $Y=0 $X2=0.895
+ $Y2=2.42
cc_30 N_VNB_M1002_b N_A_1212_471#_c_743_n 0.00164171f $X=-0.33 $Y=-0.265
+ $X2=1.645 $Y2=2.84
cc_31 N_VNB_M1002_b N_A_1212_471#_c_744_n 0.00125919f $X=-0.33 $Y=-0.265
+ $X2=1.73 $Y2=2.755
cc_32 N_VNB_M1002_b N_A_1212_471#_c_745_n 0.0206396f $X=-0.33 $Y=-0.265
+ $X2=3.385 $Y2=2.395
cc_33 N_VNB_M1002_b N_A_1212_471#_c_746_n 0.0105885f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_M1002_b N_A_1212_471#_M1001_g 0.0828107f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_35 N_VNB_M1002_b N_A_1212_100#_M1022_g 0.0960701f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=3.455
cc_36 N_VNB_M1002_b N_A_1212_100#_c_977_n 0.0464356f $X=-0.33 $Y=-0.265
+ $X2=0.895 $Y2=2.42
cc_37 N_VNB_M1002_b N_A_1212_100#_c_978_n 0.0700245f $X=-0.33 $Y=-0.265
+ $X2=1.645 $Y2=2.84
cc_38 N_VNB_M1002_b N_A_1212_100#_c_979_n 0.00388201f $X=-0.33 $Y=-0.265
+ $X2=2.645 $Y2=2.48
cc_39 N_VNB_M1002_b N_A_1212_100#_M1000_g 0.0487114f $X=-0.33 $Y=-0.265 $X2=2.73
+ $Y2=2.395
cc_40 N_VNB_M1002_b N_A_1212_100#_c_981_n 0.00538479f $X=-0.33 $Y=-0.265
+ $X2=5.32 $Y2=3.37
cc_41 N_VNB_M1002_b N_A_1212_100#_c_982_n 0.0207377f $X=-0.33 $Y=-0.265 $X2=5.32
+ $Y2=3.37
cc_42 N_VNB_M1002_b N_A_1212_100#_c_983_n 0.00211404f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_M1002_b N_A_1212_100#_c_984_n 0.139475f $X=-0.33 $Y=-0.265 $X2=2.645
+ $Y2=1.18
cc_44 N_VNB_c_8_p N_A_1212_100#_c_984_n 0.0056467f $X=0.24 $Y=0 $X2=2.645
+ $Y2=1.18
cc_45 N_VNB_M1002_b N_A_1212_100#_c_986_n 0.013657f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_c_8_p N_A_1212_100#_c_986_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_47 N_VNB_M1002_b N_A_1212_100#_c_988_n 0.00132454f $X=-0.33 $Y=-0.265
+ $X2=2.645 $Y2=1.26
cc_48 N_VNB_M1002_b N_A_1212_100#_c_989_n 0.00854752f $X=-0.33 $Y=-0.265
+ $X2=2.71 $Y2=1.57
cc_49 N_VNB_M1002_b N_A_1212_100#_c_990_n 0.01797f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_M1002_b N_A_1212_100#_c_991_n 0.00302887f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_51 N_VNB_M1002_b N_A_1212_100#_c_992_n 0.081145f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_52 N_VNB_c_8_p N_A_1212_100#_c_992_n 0.00387355f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_53 N_VNB_M1002_b N_A_1212_100#_c_994_n 0.00699849f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_54 N_VNB_c_8_p N_A_1212_100#_c_994_n 3.76524e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_55 N_VNB_M1002_b N_A_1212_100#_c_996_n 0.0073834f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_56 N_VNB_M1002_b N_A_1212_100#_c_997_n 0.019981f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_57 N_VNB_M1002_b N_A_1212_100#_c_998_n 0.00229636f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_58 N_VNB_M1002_b N_A_1212_100#_c_999_n 0.0032059f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_59 N_VNB_M1002_b N_A_1212_100#_c_1000_n 0.0933385f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_60 N_VNB_M1002_b N_A_1212_100#_c_1001_n 4.5649e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_61 N_VNB_M1002_b N_A_1510_100#_M1010_g 0.0826366f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=3.455
cc_62 N_VNB_M1002_b N_A_1510_100#_c_1246_n 0.0089999f $X=-0.33 $Y=-0.265
+ $X2=0.895 $Y2=2.42
cc_63 N_VNB_M1002_b N_A_1510_100#_c_1247_n 0.0036955f $X=-0.33 $Y=-0.265
+ $X2=2.48 $Y2=1.18
cc_64 N_VNB_M1002_b N_A_1510_100#_c_1248_n 0.0060064f $X=-0.33 $Y=-0.265
+ $X2=2.645 $Y2=2.755
cc_65 N_VNB_M1002_b N_RESET_B_M1024_g 0.0563847f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=3.455
cc_66 N_VNB_M1002_b N_RESET_B_c_1352_n 0.245068f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=3.455
cc_67 N_VNB_M1002_b N_RESET_B_c_1353_n 0.168061f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_68 N_VNB_c_8_p N_RESET_B_c_1353_n 0.0723707f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_69 N_VNB_M1002_b N_RESET_B_M1013_g 0.0432866f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_70 N_VNB_M1002_b N_RESET_B_c_1356_n 0.0263363f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_71 N_VNB_M1002_b N_RESET_B_c_1357_n 0.0576097f $X=-0.33 $Y=-0.265 $X2=1.73
+ $Y2=1.265
cc_72 N_VNB_M1002_b N_RESET_B_c_1358_n 0.0231236f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_73 N_VNB_M1002_b N_RESET_B_c_1359_n 0.0274543f $X=-0.33 $Y=-0.265 $X2=5.37
+ $Y2=0.84
cc_74 N_VNB_M1002_b N_RESET_B_M1025_g 0.0797996f $X=-0.33 $Y=-0.265 $X2=2.645
+ $Y2=1.57
cc_75 N_VNB_M1002_b N_A_1312_126#_M1007_g 0.0645191f $X=-0.33 $Y=-0.265 $X2=2.71
+ $Y2=0.84
cc_76 N_VNB_c_8_p N_A_1312_126#_M1007_g 4.06814e-19 $X=0.24 $Y=0 $X2=2.71
+ $Y2=0.84
cc_77 N_VNB_M1002_b N_A_1312_126#_c_1562_n 0.0157393f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_78 N_VNB_M1002_b N_A_1312_126#_c_1563_n 0.0102875f $X=-0.33 $Y=-0.265
+ $X2=0.895 $Y2=2.42
cc_79 N_VNB_M1002_b N_A_1312_126#_c_1564_n 0.00101051f $X=-0.33 $Y=-0.265
+ $X2=5.155 $Y2=2.79
cc_80 N_VNB_M1002_b N_A_2616_417#_c_1689_n 0.00371478f $X=-0.33 $Y=-0.265
+ $X2=2.56 $Y2=2.84
cc_81 N_VNB_M1002_b N_A_2616_417#_c_1690_n 0.0096685f $X=-0.33 $Y=-0.265
+ $X2=2.73 $Y2=2.395
cc_82 N_VNB_M1002_b N_A_2616_417#_M1021_g 0.0776962f $X=-0.33 $Y=-0.265
+ $X2=5.155 $Y2=2.79
cc_83 N_VNB_M1002_b N_A_2360_115#_M1031_g 0.0373896f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=3.455
cc_84 N_VNB_M1002_b N_A_2360_115#_M1005_g 0.0595559f $X=-0.33 $Y=-0.265 $X2=1.06
+ $Y2=2.84
cc_85 N_VNB_M1002_b N_A_2360_115#_c_1783_n 0.0630517f $X=-0.33 $Y=-0.265
+ $X2=1.73 $Y2=2.755
cc_86 N_VNB_M1002_b N_A_2360_115#_c_1784_n 0.0295498f $X=-0.33 $Y=-0.265
+ $X2=2.48 $Y2=1.18
cc_87 N_VNB_M1002_b N_A_2360_115#_c_1785_n 0.00252127f $X=-0.33 $Y=-0.265
+ $X2=1.815 $Y2=2.84
cc_88 N_VNB_M1002_b N_A_2360_115#_c_1786_n 0.00415983f $X=-0.33 $Y=-0.265
+ $X2=3.385 $Y2=2.395
cc_89 N_VNB_M1002_b N_A_2360_115#_c_1787_n 0.0251951f $X=-0.33 $Y=-0.265
+ $X2=2.645 $Y2=1.57
cc_90 N_VNB_M1002_b N_A_2360_115#_c_1788_n 0.00346004f $X=-0.33 $Y=-0.265
+ $X2=2.71 $Y2=1.57
cc_91 N_VNB_M1002_b N_A_2360_115#_c_1789_n 0.0426543f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_92 N_VNB_M1002_b N_CLK_c_1958_n 0.0911742f $X=-0.33 $Y=-0.265 $X2=5.23
+ $Y2=0.63
cc_93 N_VNB_c_8_p N_CLK_c_1958_n 9.82187e-19 $X=0.24 $Y=0 $X2=5.23 $Y2=0.63
cc_94 N_VNB_M1002_b N_CLK_c_1960_n 0.0616573f $X=-0.33 $Y=-0.265 $X2=2.71
+ $Y2=0.84
cc_95 N_VNB_M1002_b N_A_3417_443#_M1034_g 0.0479335f $X=-0.33 $Y=-0.265 $X2=2.71
+ $Y2=0.84
cc_96 N_VNB_c_8_p N_A_3417_443#_M1034_g 6.79573e-19 $X=0.24 $Y=0 $X2=2.71
+ $Y2=0.84
cc_97 N_VNB_M1002_b N_A_3417_443#_c_1997_n 0.00673533f $X=-0.33 $Y=-0.265
+ $X2=0.895 $Y2=2.755
cc_98 N_VNB_M1002_b N_A_3417_443#_c_1998_n 0.00185187f $X=-0.33 $Y=-0.265
+ $X2=1.645 $Y2=2.84
cc_99 N_VNB_M1002_b N_A_3417_443#_c_1999_n 0.0078064f $X=-0.33 $Y=-0.265
+ $X2=1.815 $Y2=1.18
cc_100 N_VNB_M1002_b N_A_3417_443#_c_2000_n 0.046267f $X=-0.33 $Y=-0.265
+ $X2=2.56 $Y2=2.84
cc_101 N_VNB_M1002_b N_A_65_649#_c_2046_n 0.00128013f $X=-0.33 $Y=-0.265
+ $X2=0.895 $Y2=2.42
cc_102 N_VNB_M1002_b N_A_65_649#_c_2047_n 0.0124353f $X=-0.33 $Y=-0.265 $X2=1.73
+ $Y2=1.265
cc_103 N_VNB_M1002_b N_A_65_649#_c_2048_n 0.00903544f $X=-0.33 $Y=-0.265
+ $X2=1.73 $Y2=2.755
cc_104 N_VNB_M1002_b N_A_65_649#_c_2049_n 0.00176659f $X=-0.33 $Y=-0.265
+ $X2=3.385 $Y2=2.395
cc_105 N_VNB_M1002_b N_A_65_649#_c_2050_n 0.012636f $X=-0.33 $Y=-0.265 $X2=1.73
+ $Y2=2.84
cc_106 N_VNB_c_8_p N_A_65_649#_c_2050_n 5.66018e-19 $X=0.24 $Y=0 $X2=1.73
+ $Y2=2.84
cc_107 N_VNB_M1002_b N_A_65_649#_c_2052_n 0.00269919f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_108 N_VNB_M1002_b N_A_65_649#_c_2053_n 0.0183163f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_109 N_VNB_M1002_b N_Q_c_2350_n 0.066486f $X=-0.33 $Y=-0.265 $X2=1.73
+ $Y2=1.265
cc_110 N_VNB_c_8_p N_Q_c_2350_n 5.76324e-19 $X=0.24 $Y=0 $X2=1.73 $Y2=1.265
cc_111 N_VNB_M1002_b N_noxref_23_c_2364_n 0.0183118f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=3.455
cc_112 N_VNB_M1002_b N_noxref_23_c_2365_n 0.244042f $X=-0.33 $Y=-0.265 $X2=2.71
+ $Y2=1.315
cc_113 N_VNB_c_8_p N_noxref_23_c_2365_n 0.0100829f $X=0.24 $Y=0 $X2=2.71
+ $Y2=1.315
cc_114 N_VNB_M1002_b N_noxref_23_c_2367_n 0.0269123f $X=-0.33 $Y=-0.265 $X2=2.71
+ $Y2=0.84
cc_115 N_VNB_c_8_p N_noxref_23_c_2367_n 0.00109438f $X=0.24 $Y=0 $X2=2.71
+ $Y2=0.84
cc_116 N_VNB_M1002_b N_noxref_23_c_2369_n 8.23828e-19 $X=-0.33 $Y=-0.265
+ $X2=0.895 $Y2=2.755
cc_117 N_VNB_M1002_b N_VGND_c_2396_n 0.0449686f $X=-0.33 $Y=-0.265 $X2=1.73
+ $Y2=1.265
cc_118 N_VNB_c_8_p N_VGND_c_2396_n 0.00324287f $X=0.24 $Y=0 $X2=1.73 $Y2=1.265
cc_119 N_VNB_M1002_b N_VGND_c_2398_n 0.0585438f $X=-0.33 $Y=-0.265 $X2=2.73
+ $Y2=2.395
cc_120 N_VNB_c_8_p N_VGND_c_2398_n 0.00362764f $X=0.24 $Y=0 $X2=2.73 $Y2=2.395
cc_121 N_VNB_M1002_b N_VGND_c_2400_n 0.0467653f $X=-0.33 $Y=-0.265 $X2=5.32
+ $Y2=3.37
cc_122 N_VNB_c_8_p N_VGND_c_2400_n 0.00166879f $X=0.24 $Y=0 $X2=5.32 $Y2=3.37
cc_123 N_VNB_M1002_b N_VGND_c_2402_n 0.0690249f $X=-0.33 $Y=-0.265 $X2=2.645
+ $Y2=1.26
cc_124 N_VNB_c_8_p N_VGND_c_2402_n 0.00269049f $X=0.24 $Y=0 $X2=2.645 $Y2=1.26
cc_125 N_VNB_M1002_b N_VGND_c_2404_n 0.0439913f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_126 N_VNB_c_8_p N_VGND_c_2404_n 0.00167079f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_127 N_VNB_M1002_b N_VGND_c_2406_n 0.058498f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_128 N_VNB_c_8_p N_VGND_c_2406_n 0.00257697f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_129 N_VNB_M1002_b N_VGND_c_2408_n 0.28668f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_130 N_VNB_c_8_p N_VGND_c_2408_n 2.0446f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_131 N_VPB_M1008_b N_A_116_451#_c_347_n 0.0950601f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=3.115
cc_132 N_VPB_M1008_b N_A_116_451#_M1008_g 0.0412306f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=3.455
cc_133 VPB N_A_116_451#_M1008_g 0.00274588f $X=0 $Y=3.955 $X2=0.86 $Y2=3.455
cc_134 N_VPB_c_134_p N_A_116_451#_M1008_g 0.0142077f $X=18.96 $Y=4.07 $X2=0.86
+ $Y2=3.455
cc_135 N_VPB_M1008_b N_A_116_451#_c_351_n 0.00335562f $X=-0.33 $Y=1.885
+ $X2=0.895 $Y2=2.42
cc_136 N_VPB_M1008_b N_A_116_451#_c_352_n 0.00789107f $X=-0.33 $Y=1.885
+ $X2=1.645 $Y2=2.84
cc_137 N_VPB_M1008_b N_A_116_451#_c_341_n 0.00189781f $X=-0.33 $Y=1.885 $X2=1.73
+ $Y2=2.755
cc_138 N_VPB_M1008_b N_A_116_451#_c_354_n 0.01149f $X=-0.33 $Y=1.885 $X2=2.56
+ $Y2=2.84
cc_139 N_VPB_M1008_b N_A_116_451#_c_355_n 0.00209982f $X=-0.33 $Y=1.885
+ $X2=2.645 $Y2=2.755
cc_140 N_VPB_M1008_b N_A_116_451#_c_356_n 0.00994816f $X=-0.33 $Y=1.885
+ $X2=3.385 $Y2=2.395
cc_141 N_VPB_M1008_b N_A_116_451#_c_357_n 0.00101481f $X=-0.33 $Y=1.885 $X2=2.73
+ $Y2=2.395
cc_142 N_VPB_M1008_b N_A_116_451#_c_358_n 0.00401429f $X=-0.33 $Y=1.885 $X2=3.47
+ $Y2=2.705
cc_143 N_VPB_M1008_b N_A_116_451#_c_359_n 0.0119787f $X=-0.33 $Y=1.885 $X2=5.155
+ $Y2=2.79
cc_144 N_VPB_M1008_b N_A_116_451#_c_360_n 0.00281857f $X=-0.33 $Y=1.885
+ $X2=3.555 $Y2=2.79
cc_145 N_VPB_M1008_b N_A_116_451#_c_361_n 0.00723684f $X=-0.33 $Y=1.885 $X2=5.32
+ $Y2=3.37
cc_146 N_VPB_M1008_b N_SCD_c_501_n 0.0856942f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_147 N_VPB_M1008_b N_SCD_M1011_g 0.0983667f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=3.455
cc_148 VPB N_SCD_M1011_g 0.00274588f $X=0 $Y=3.955 $X2=0.86 $Y2=3.455
cc_149 N_VPB_c_134_p N_SCD_M1011_g 0.0102234f $X=18.96 $Y=4.07 $X2=0.86
+ $Y2=3.455
cc_150 N_VPB_M1008_b N_SCE_c_560_n 0.0760267f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_151 N_VPB_M1008_b N_SCE_M1035_g 0.0739022f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=3.115
cc_152 VPB N_SCE_M1035_g 0.00274588f $X=0 $Y=3.955 $X2=0.86 $Y2=3.115
cc_153 N_VPB_c_134_p N_SCE_M1035_g 0.0111766f $X=18.96 $Y=4.07 $X2=0.86
+ $Y2=3.115
cc_154 N_VPB_M1008_b N_SCE_M1014_g 0.100959f $X=-0.33 $Y=1.885 $X2=2.71
+ $Y2=1.315
cc_155 VPB N_SCE_M1014_g 7.03951e-19 $X=0 $Y=3.955 $X2=2.71 $Y2=1.315
cc_156 N_VPB_c_134_p N_SCE_M1014_g 0.00595623f $X=18.96 $Y=4.07 $X2=2.71
+ $Y2=1.315
cc_157 N_VPB_M1008_b N_SCE_c_567_n 0.0560973f $X=-0.33 $Y=1.885 $X2=0.895
+ $Y2=2.755
cc_158 N_VPB_M1008_b N_SCE_c_568_n 0.00386088f $X=-0.33 $Y=1.885 $X2=1.73
+ $Y2=2.755
cc_159 N_VPB_M1008_b N_SCE_c_554_n 0.00770083f $X=-0.33 $Y=1.885 $X2=2.56
+ $Y2=2.84
cc_160 N_VPB_M1008_b N_SCE_c_555_n 8.79775e-19 $X=-0.33 $Y=1.885 $X2=2.645
+ $Y2=2.48
cc_161 N_VPB_M1008_b SCE 0.00155029f $X=-0.33 $Y=1.885 $X2=2.645 $Y2=2.755
cc_162 N_VPB_M1008_b SCE 0.0186374f $X=-0.33 $Y=1.885 $X2=2.81 $Y2=1.26
cc_163 N_VPB_M1008_b N_SCE_M1012_g 0.0168861f $X=-0.33 $Y=1.885 $X2=5.41
+ $Y2=0.84
cc_164 N_VPB_M1008_b N_D_c_681_n 0.0340729f $X=-0.33 $Y=1.885 $X2=5.23 $Y2=0.63
cc_165 N_VPB_M1008_b N_D_M1004_g 0.0334433f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_166 N_VPB_M1008_b N_D_c_683_n 0.110942f $X=-0.33 $Y=1.885 $X2=0.895 $Y2=2.755
cc_167 VPB N_D_c_683_n 0.00274588f $X=0 $Y=3.955 $X2=0.895 $Y2=2.755
cc_168 N_VPB_c_134_p N_D_c_683_n 0.00916369f $X=18.96 $Y=4.07 $X2=0.895
+ $Y2=2.755
cc_169 N_VPB_M1008_b N_A_1212_471#_c_737_n 0.0332704f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=3.115
cc_170 N_VPB_M1008_b N_A_1212_471#_c_738_n 0.00376437f $X=-0.33 $Y=1.885
+ $X2=2.71 $Y2=0.84
cc_171 N_VPB_M1008_b N_A_1212_471#_c_750_n 0.111421f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_172 VPB N_A_1212_471#_c_750_n 6.67351e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_173 N_VPB_c_134_p N_A_1212_471#_c_750_n 0.00545833f $X=18.96 $Y=4.07 $X2=0
+ $Y2=0
cc_174 N_VPB_M1008_b N_A_1212_471#_c_753_n 0.00472847f $X=-0.33 $Y=1.885
+ $X2=0.895 $Y2=2.42
cc_175 VPB N_A_1212_471#_c_753_n 0.00290046f $X=0 $Y=3.955 $X2=0.895 $Y2=2.42
cc_176 N_VPB_c_134_p N_A_1212_471#_c_753_n 0.0568137f $X=18.96 $Y=4.07 $X2=0.895
+ $Y2=2.42
cc_177 N_VPB_M1008_b N_A_1212_471#_c_756_n 7.83871e-19 $X=-0.33 $Y=1.885
+ $X2=0.895 $Y2=2.42
cc_178 VPB N_A_1212_471#_c_756_n 5.70856e-19 $X=0 $Y=3.955 $X2=0.895 $Y2=2.42
cc_179 N_VPB_c_134_p N_A_1212_471#_c_756_n 0.0114989f $X=18.96 $Y=4.07 $X2=0.895
+ $Y2=2.42
cc_180 N_VPB_M1008_b N_A_1212_471#_c_759_n 0.00488603f $X=-0.33 $Y=1.885
+ $X2=2.645 $Y2=2.48
cc_181 N_VPB_M1008_b N_A_1212_471#_c_760_n 0.0125808f $X=-0.33 $Y=1.885 $X2=3.47
+ $Y2=2.48
cc_182 VPB N_A_1212_471#_c_760_n 0.00363377f $X=0 $Y=3.955 $X2=3.47 $Y2=2.48
cc_183 N_VPB_c_134_p N_A_1212_471#_c_760_n 0.0715819f $X=18.96 $Y=4.07 $X2=3.47
+ $Y2=2.48
cc_184 N_VPB_M1008_b N_A_1212_471#_c_763_n 0.00125214f $X=-0.33 $Y=1.885
+ $X2=3.47 $Y2=2.705
cc_185 VPB N_A_1212_471#_c_763_n 5.70856e-19 $X=0 $Y=3.955 $X2=3.47 $Y2=2.705
cc_186 N_VPB_c_134_p N_A_1212_471#_c_763_n 0.0114989f $X=18.96 $Y=4.07 $X2=3.47
+ $Y2=2.705
cc_187 N_VPB_M1008_b N_A_1212_471#_c_766_n 0.00612843f $X=-0.33 $Y=1.885
+ $X2=5.32 $Y2=2.875
cc_188 N_VPB_M1008_b N_A_1212_471#_c_767_n 0.00464967f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_189 N_VPB_M1008_b N_A_1212_471#_c_768_n 0.00279041f $X=-0.33 $Y=1.885
+ $X2=1.73 $Y2=2.84
cc_190 N_VPB_M1008_b N_A_1212_471#_c_769_n 0.0109653f $X=-0.33 $Y=1.885
+ $X2=2.645 $Y2=1.57
cc_191 N_VPB_M1008_b N_A_1212_471#_c_770_n 0.0880589f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_192 N_VPB_M1008_b N_A_1212_471#_c_771_n 0.00167974f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_193 N_VPB_M1008_b N_A_1212_471#_c_772_n 0.00458706f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_194 N_VPB_M1008_b N_A_1212_100#_M1022_g 0.00623548f $X=-0.33 $Y=1.885
+ $X2=0.86 $Y2=3.455
cc_195 N_VPB_M1008_b N_A_1212_100#_c_1003_n 0.0198854f $X=-0.33 $Y=1.885
+ $X2=2.71 $Y2=1.315
cc_196 N_VPB_M1008_b N_A_1212_100#_c_1004_n 0.0211544f $X=-0.33 $Y=1.885
+ $X2=2.71 $Y2=0.84
cc_197 N_VPB_M1008_b N_A_1212_100#_c_1005_n 0.0689635f $X=-0.33 $Y=1.885
+ $X2=2.71 $Y2=0.84
cc_198 N_VPB_M1008_b N_A_1212_100#_M1003_g 0.0706805f $X=-0.33 $Y=1.885
+ $X2=0.895 $Y2=2.755
cc_199 VPB N_A_1212_100#_M1003_g 6.67351e-19 $X=0 $Y=3.955 $X2=0.895 $Y2=2.755
cc_200 N_VPB_c_134_p N_A_1212_100#_M1003_g 0.00545833f $X=18.96 $Y=4.07
+ $X2=0.895 $Y2=2.755
cc_201 N_VPB_M1008_b N_A_1212_100#_c_978_n 0.120389f $X=-0.33 $Y=1.885 $X2=1.645
+ $Y2=2.84
cc_202 N_VPB_M1008_b N_A_1212_100#_M1020_g 0.0419015f $X=-0.33 $Y=1.885 $X2=1.73
+ $Y2=1.265
cc_203 VPB N_A_1212_100#_M1020_g 7.76601e-19 $X=0 $Y=3.955 $X2=1.73 $Y2=1.265
cc_204 N_VPB_c_134_p N_A_1212_100#_M1020_g 0.00498289f $X=18.96 $Y=4.07 $X2=1.73
+ $Y2=1.265
cc_205 N_VPB_M1008_b N_A_1212_100#_c_1013_n 0.037113f $X=-0.33 $Y=1.885 $X2=2.48
+ $Y2=1.18
cc_206 VPB N_A_1212_100#_c_1013_n 0.00970178f $X=0 $Y=3.955 $X2=2.48 $Y2=1.18
cc_207 N_VPB_c_134_p N_A_1212_100#_c_1013_n 0.0196751f $X=18.96 $Y=4.07 $X2=2.48
+ $Y2=1.18
cc_208 N_VPB_M1008_b N_A_1212_100#_c_979_n 0.0755202f $X=-0.33 $Y=1.885
+ $X2=2.645 $Y2=2.48
cc_209 N_VPB_M1008_b N_A_1212_100#_c_981_n 0.00133253f $X=-0.33 $Y=1.885
+ $X2=5.32 $Y2=3.37
cc_210 N_VPB_M1008_b N_A_1212_100#_c_1018_n 0.0442962f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_211 VPB N_A_1212_100#_c_1018_n 5.2689e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_212 N_VPB_c_134_p N_A_1212_100#_c_1018_n 0.00566149f $X=18.96 $Y=4.07 $X2=0
+ $Y2=0
cc_213 N_VPB_M1008_b N_A_1212_100#_c_1021_n 0.0178718f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_214 N_VPB_M1008_b N_A_1212_100#_c_1022_n 0.00231118f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_215 N_VPB_M1008_b N_A_1212_100#_c_1023_n 0.00795184f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_216 N_VPB_M1008_b N_A_1510_100#_M1015_g 0.0829281f $X=-0.33 $Y=1.885 $X2=2.71
+ $Y2=0.84
cc_217 VPB N_A_1510_100#_M1015_g 0.00260111f $X=0 $Y=3.955 $X2=2.71 $Y2=0.84
cc_218 N_VPB_c_134_p N_A_1510_100#_M1015_g 0.00850026f $X=18.96 $Y=4.07 $X2=2.71
+ $Y2=0.84
cc_219 N_VPB_M1008_b N_A_1510_100#_c_1246_n 0.00923706f $X=-0.33 $Y=1.885
+ $X2=0.895 $Y2=2.42
cc_220 N_VPB_M1008_b N_A_1510_100#_c_1253_n 0.00242911f $X=-0.33 $Y=1.885
+ $X2=2.56 $Y2=2.84
cc_221 N_VPB_M1008_b N_A_1510_100#_c_1248_n 0.0660905f $X=-0.33 $Y=1.885
+ $X2=2.645 $Y2=2.755
cc_222 N_VPB_M1008_b N_A_1510_100#_c_1255_n 9.67407e-19 $X=-0.33 $Y=1.885
+ $X2=2.73 $Y2=2.395
cc_223 N_VPB_M1008_b N_A_1510_100#_c_1256_n 0.00219526f $X=-0.33 $Y=1.885
+ $X2=3.47 $Y2=2.705
cc_224 N_VPB_M1008_b N_RESET_B_M1019_g 0.0401447f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_225 VPB N_RESET_B_M1019_g 0.00274588f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_226 N_VPB_c_134_p N_RESET_B_M1019_g 0.0104883f $X=18.96 $Y=4.07 $X2=0 $Y2=0
cc_227 N_VPB_M1008_b N_RESET_B_c_1364_n 0.0869413f $X=-0.33 $Y=1.885 $X2=0.895
+ $Y2=2.42
cc_228 N_VPB_M1008_b N_RESET_B_c_1365_n 0.0296814f $X=-0.33 $Y=1.885 $X2=1.815
+ $Y2=1.18
cc_229 N_VPB_M1008_b N_RESET_B_c_1366_n 0.00274587f $X=-0.33 $Y=1.885 $X2=2.56
+ $Y2=2.84
cc_230 N_VPB_M1008_b N_RESET_B_c_1367_n 0.0401431f $X=-0.33 $Y=1.885 $X2=1.815
+ $Y2=2.84
cc_231 N_VPB_M1008_b N_RESET_B_c_1368_n 0.00125284f $X=-0.33 $Y=1.885 $X2=2.645
+ $Y2=2.48
cc_232 N_VPB_M1008_b N_RESET_B_c_1369_n 0.00903646f $X=-0.33 $Y=1.885 $X2=2.73
+ $Y2=2.395
cc_233 N_VPB_M1008_b N_RESET_B_c_1370_n 8.73552e-19 $X=-0.33 $Y=1.885 $X2=3.555
+ $Y2=2.79
cc_234 N_VPB_M1008_b N_RESET_B_c_1358_n 0.0548933f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_235 N_VPB_M1008_b N_RESET_B_c_1359_n 0.150766f $X=-0.33 $Y=1.885 $X2=5.37
+ $Y2=0.84
cc_236 VPB N_RESET_B_c_1359_n 6.67351e-19 $X=0 $Y=3.955 $X2=5.37 $Y2=0.84
cc_237 N_VPB_c_134_p N_RESET_B_c_1359_n 0.00545833f $X=18.96 $Y=4.07 $X2=5.37
+ $Y2=0.84
cc_238 N_VPB_M1008_b N_RESET_B_c_1375_n 0.00329874f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_239 N_VPB_M1008_b N_RESET_B_M1025_g 0.101381f $X=-0.33 $Y=1.885 $X2=2.645
+ $Y2=1.57
cc_240 N_VPB_M1008_b N_A_1312_126#_c_1562_n 0.114783f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_241 VPB N_A_1312_126#_c_1562_n 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_242 N_VPB_c_134_p N_A_1312_126#_c_1562_n 0.0163911f $X=18.96 $Y=4.07 $X2=0
+ $Y2=0
cc_243 N_VPB_M1008_b N_A_1312_126#_c_1563_n 0.00765988f $X=-0.33 $Y=1.885
+ $X2=0.895 $Y2=2.42
cc_244 N_VPB_M1008_b N_A_1312_126#_c_1569_n 0.01103f $X=-0.33 $Y=1.885 $X2=1.73
+ $Y2=2.755
cc_245 N_VPB_M1008_b N_A_1312_126#_c_1570_n 0.00639551f $X=-0.33 $Y=1.885
+ $X2=1.815 $Y2=2.84
cc_246 N_VPB_M1008_b N_A_1312_126#_c_1571_n 0.00678755f $X=-0.33 $Y=1.885
+ $X2=3.385 $Y2=2.395
cc_247 N_VPB_M1008_b N_A_1312_126#_c_1572_n 0.00496598f $X=-0.33 $Y=1.885
+ $X2=2.73 $Y2=2.395
cc_248 N_VPB_M1008_b N_A_1312_126#_c_1573_n 0.00273461f $X=-0.33 $Y=1.885
+ $X2=5.285 $Y2=1.26
cc_249 N_VPB_M1008_b N_A_1312_126#_c_1574_n 6.92236e-19 $X=-0.33 $Y=1.885
+ $X2=5.32 $Y2=2.875
cc_250 N_VPB_M1008_b N_A_1312_126#_c_1575_n 0.00399078f $X=-0.33 $Y=1.885
+ $X2=5.32 $Y2=3.37
cc_251 N_VPB_M1008_b N_A_2616_417#_M1039_g 0.0347213f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=3.455
cc_252 N_VPB_M1008_b N_A_2616_417#_c_1693_n 0.0577263f $X=-0.33 $Y=1.885
+ $X2=2.71 $Y2=0.84
cc_253 N_VPB_M1008_b N_A_2616_417#_c_1694_n 9.80592e-19 $X=-0.33 $Y=1.885
+ $X2=0.895 $Y2=2.42
cc_254 N_VPB_M1008_b N_A_2616_417#_c_1695_n 0.00332854f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_255 N_VPB_M1008_b N_A_2616_417#_c_1696_n 0.00210811f $X=-0.33 $Y=1.885
+ $X2=1.73 $Y2=2.755
cc_256 N_VPB_M1008_b N_A_2616_417#_c_1689_n 0.00758668f $X=-0.33 $Y=1.885
+ $X2=2.56 $Y2=2.84
cc_257 N_VPB_M1008_b N_A_2616_417#_c_1698_n 0.00250004f $X=-0.33 $Y=1.885
+ $X2=2.645 $Y2=2.755
cc_258 N_VPB_M1008_b N_A_2616_417#_M1021_g 0.0207891f $X=-0.33 $Y=1.885
+ $X2=5.155 $Y2=2.79
cc_259 N_VPB_M1008_b N_A_2360_115#_M1028_g 0.0690498f $X=-0.33 $Y=1.885 $X2=2.71
+ $Y2=0.84
cc_260 N_VPB_M1008_b N_A_2360_115#_M1029_g 0.0489072f $X=-0.33 $Y=1.885
+ $X2=0.895 $Y2=2.42
cc_261 N_VPB_M1008_b N_A_2360_115#_c_1783_n 0.0453416f $X=-0.33 $Y=1.885
+ $X2=1.73 $Y2=2.755
cc_262 N_VPB_M1008_b N_A_2360_115#_c_1784_n 0.0170569f $X=-0.33 $Y=1.885
+ $X2=2.48 $Y2=1.18
cc_263 N_VPB_M1008_b N_A_2360_115#_c_1786_n 5.4194e-19 $X=-0.33 $Y=1.885
+ $X2=3.385 $Y2=2.395
cc_264 N_VPB_M1008_b N_A_2360_115#_c_1795_n 0.00563403f $X=-0.33 $Y=1.885
+ $X2=2.81 $Y2=1.26
cc_265 N_VPB_M1008_b N_A_2360_115#_c_1796_n 0.0153015f $X=-0.33 $Y=1.885
+ $X2=3.47 $Y2=2.705
cc_266 N_VPB_M1008_b N_A_2360_115#_c_1797_n 0.00603245f $X=-0.33 $Y=1.885
+ $X2=5.155 $Y2=2.79
cc_267 N_VPB_M1008_b N_A_2360_115#_c_1798_n 0.00418149f $X=-0.33 $Y=1.885
+ $X2=5.32 $Y2=2.875
cc_268 N_VPB_M1008_b N_A_2360_115#_c_1799_n 0.00141351f $X=-0.33 $Y=1.885
+ $X2=5.32 $Y2=3.37
cc_269 N_VPB_M1008_b N_A_2360_115#_c_1800_n 7.61606e-19 $X=-0.33 $Y=1.885
+ $X2=5.32 $Y2=3.37
cc_270 N_VPB_M1008_b N_A_2360_115#_c_1801_n 0.00433192f $X=-0.33 $Y=1.885
+ $X2=5.41 $Y2=1.175
cc_271 N_VPB_M1008_b N_A_2360_115#_c_1802_n 0.0168129f $X=-0.33 $Y=1.885
+ $X2=5.41 $Y2=0.84
cc_272 VPB N_A_2360_115#_c_1802_n 0.00173699f $X=0 $Y=3.955 $X2=5.41 $Y2=0.84
cc_273 N_VPB_c_134_p N_A_2360_115#_c_1802_n 0.0184698f $X=18.96 $Y=4.07 $X2=5.41
+ $Y2=0.84
cc_274 N_VPB_M1008_b N_A_2360_115#_c_1805_n 0.00342771f $X=-0.33 $Y=1.885
+ $X2=5.37 $Y2=0.84
cc_275 VPB N_A_2360_115#_c_1805_n 3.7339e-19 $X=0 $Y=3.955 $X2=5.37 $Y2=0.84
cc_276 N_VPB_c_134_p N_A_2360_115#_c_1805_n 0.00409372f $X=18.96 $Y=4.07
+ $X2=5.37 $Y2=0.84
cc_277 N_VPB_M1008_b N_A_2360_115#_c_1808_n 0.00197943f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_278 N_VPB_M1008_b N_A_2360_115#_c_1789_n 0.0433562f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_279 N_VPB_M1008_b N_CLK_c_1960_n 0.110765f $X=-0.33 $Y=1.885 $X2=2.71
+ $Y2=0.84
cc_280 VPB N_CLK_c_1960_n 5.41292e-19 $X=0 $Y=3.955 $X2=2.71 $Y2=0.84
cc_281 N_VPB_c_134_p N_CLK_c_1960_n 0.00416385f $X=18.96 $Y=4.07 $X2=2.71
+ $Y2=0.84
cc_282 N_VPB_M1008_b N_CLK_c_1964_n 0.0122988f $X=-0.33 $Y=1.885 $X2=2.71
+ $Y2=0.84
cc_283 N_VPB_M1008_b N_A_3417_443#_M1017_g 0.042212f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=3.455
cc_284 VPB N_A_3417_443#_M1017_g 0.00970178f $X=0 $Y=3.955 $X2=0.86 $Y2=3.455
cc_285 N_VPB_c_134_p N_A_3417_443#_M1017_g 0.0152133f $X=18.96 $Y=4.07 $X2=0.86
+ $Y2=3.455
cc_286 N_VPB_M1008_b N_A_3417_443#_c_2000_n 0.0214997f $X=-0.33 $Y=1.885
+ $X2=2.56 $Y2=2.84
cc_287 N_VPB_M1008_b N_A_3417_443#_c_2005_n 0.0161907f $X=-0.33 $Y=1.885
+ $X2=2.645 $Y2=2.755
cc_288 N_VPB_M1008_b N_A_65_649#_c_2046_n 0.0643478f $X=-0.33 $Y=1.885 $X2=0.895
+ $Y2=2.42
cc_289 N_VPB_M1008_b N_A_65_649#_c_2055_n 0.011693f $X=-0.33 $Y=1.885 $X2=1.645
+ $Y2=2.84
cc_290 VPB N_A_65_649#_c_2055_n 9.76027e-19 $X=0 $Y=3.955 $X2=1.645 $Y2=2.84
cc_291 N_VPB_c_134_p N_A_65_649#_c_2055_n 0.0140766f $X=18.96 $Y=4.07 $X2=1.645
+ $Y2=2.84
cc_292 N_VPB_M1008_b N_A_65_649#_c_2058_n 0.00645809f $X=-0.33 $Y=1.885 $X2=2.48
+ $Y2=1.18
cc_293 N_VPB_M1008_b N_A_65_649#_c_2059_n 0.00188552f $X=-0.33 $Y=1.885 $X2=3.47
+ $Y2=2.48
cc_294 VPB N_A_65_649#_c_2059_n 0.00303599f $X=0 $Y=3.955 $X2=3.47 $Y2=2.48
cc_295 N_VPB_c_134_p N_A_65_649#_c_2059_n 0.0332751f $X=18.96 $Y=4.07 $X2=3.47
+ $Y2=2.48
cc_296 N_VPB_M1008_b N_A_65_649#_c_2062_n 5.72166e-19 $X=-0.33 $Y=1.885 $X2=3.47
+ $Y2=2.705
cc_297 VPB N_A_65_649#_c_2062_n 5.96002e-19 $X=0 $Y=3.955 $X2=3.47 $Y2=2.705
cc_298 N_VPB_c_134_p N_A_65_649#_c_2062_n 0.00708252f $X=18.96 $Y=4.07 $X2=3.47
+ $Y2=2.705
cc_299 N_VPB_M1008_b N_A_65_649#_c_2065_n 3.00334e-19 $X=-0.33 $Y=1.885 $X2=5.32
+ $Y2=3.37
cc_300 N_VPB_M1008_b N_A_65_649#_c_2066_n 0.00898534f $X=-0.33 $Y=1.885 $X2=5.32
+ $Y2=3.37
cc_301 N_VPB_M1008_b N_A_65_649#_c_2067_n 0.00292981f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_302 N_VPB_M1008_b N_A_65_649#_c_2068_n 0.0117287f $X=-0.33 $Y=1.885 $X2=5.37
+ $Y2=0.84
cc_303 VPB N_A_65_649#_c_2068_n 0.00346584f $X=0 $Y=3.955 $X2=5.37 $Y2=0.84
cc_304 N_VPB_c_134_p N_A_65_649#_c_2068_n 0.0681035f $X=18.96 $Y=4.07 $X2=5.37
+ $Y2=0.84
cc_305 N_VPB_M1008_b N_A_65_649#_c_2071_n 7.34254e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_306 VPB N_A_65_649#_c_2071_n 5.70856e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_307 N_VPB_c_134_p N_A_65_649#_c_2071_n 0.0114989f $X=18.96 $Y=4.07 $X2=0
+ $Y2=0
cc_308 N_VPB_M1008_b N_A_65_649#_c_2074_n 0.00494559f $X=-0.33 $Y=1.885
+ $X2=2.645 $Y2=1.26
cc_309 N_VPB_M1008_b N_A_65_649#_c_2075_n 0.00404383f $X=-0.33 $Y=1.885
+ $X2=2.645 $Y2=1.57
cc_310 N_VPB_M1008_b N_A_65_649#_c_2076_n 0.0116495f $X=-0.33 $Y=1.885 $X2=2.71
+ $Y2=1.57
cc_311 N_VPB_M1008_b N_A_65_649#_c_2053_n 0.0276245f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_312 N_VPB_M1008_b N_VPWR_c_2199_n 0.00157286f $X=-0.33 $Y=1.885 $X2=2.73
+ $Y2=2.395
cc_313 VPB N_VPWR_c_2199_n 0.00367725f $X=0 $Y=3.955 $X2=2.73 $Y2=2.395
cc_314 N_VPB_c_134_p N_VPWR_c_2199_n 0.0380315f $X=18.96 $Y=4.07 $X2=2.73
+ $Y2=2.395
cc_315 N_VPB_M1008_b N_VPWR_c_2202_n 0.00332161f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_316 VPB N_VPWR_c_2202_n 0.00312753f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_317 N_VPB_c_134_p N_VPWR_c_2202_n 0.0365091f $X=18.96 $Y=4.07 $X2=0 $Y2=0
cc_318 N_VPB_M1008_b N_VPWR_c_2205_n 0.00330298f $X=-0.33 $Y=1.885 $X2=2.645
+ $Y2=1.26
cc_319 VPB N_VPWR_c_2205_n 0.00348466f $X=0 $Y=3.955 $X2=2.645 $Y2=1.26
cc_320 N_VPB_c_134_p N_VPWR_c_2205_n 0.0386046f $X=18.96 $Y=4.07 $X2=2.645
+ $Y2=1.26
cc_321 N_VPB_M1008_b N_VPWR_c_2208_n 0.00411021f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_322 VPB N_VPWR_c_2208_n 0.00324688f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_323 N_VPB_c_134_p N_VPWR_c_2208_n 0.0442811f $X=18.96 $Y=4.07 $X2=0 $Y2=0
cc_324 N_VPB_M1008_b N_VPWR_c_2211_n 0.0290724f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_325 VPB N_VPWR_c_2211_n 0.0027231f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_326 N_VPB_c_134_p N_VPWR_c_2211_n 0.0404583f $X=18.96 $Y=4.07 $X2=0 $Y2=0
cc_327 N_VPB_M1008_b N_VPWR_c_2214_n 0.0245002f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_328 VPB N_VPWR_c_2214_n 0.00252021f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_329 N_VPB_c_134_p N_VPWR_c_2214_n 0.0384021f $X=18.96 $Y=4.07 $X2=0 $Y2=0
cc_330 N_VPB_M1008_b N_VPWR_c_2217_n 0.0301039f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_2217_n 0.00343155f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_332 N_VPB_c_134_p N_VPWR_c_2217_n 0.0465008f $X=18.96 $Y=4.07 $X2=0 $Y2=0
cc_333 N_VPB_M1008_b N_VPWR_c_2220_n 0.197405f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_334 VPB N_VPWR_c_2220_n 2.05015f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_335 N_VPB_c_134_p N_VPWR_c_2220_n 0.0962444f $X=18.96 $Y=4.07 $X2=0 $Y2=0
cc_336 N_VPB_M1008_b N_Q_c_2350_n 0.069368f $X=-0.33 $Y=1.885 $X2=1.73 $Y2=1.265
cc_337 VPB N_Q_c_2350_n 7.75439e-19 $X=0 $Y=3.955 $X2=1.73 $Y2=1.265
cc_338 N_VPB_c_134_p N_Q_c_2350_n 0.0133691f $X=18.96 $Y=4.07 $X2=1.73 $Y2=1.265
cc_339 N_A_116_451#_c_343_n N_SCD_c_500_n 0.00113903f $X=1.815 $Y=1.18 $X2=0
+ $Y2=0
cc_340 N_A_116_451#_c_347_n N_SCD_c_501_n 0.0181218f $X=0.86 $Y=3.115 $X2=-0.33
+ $Y2=-0.265
cc_341 N_A_116_451#_c_351_n N_SCD_c_501_n 0.00111141f $X=0.895 $Y=2.42 $X2=-0.33
+ $Y2=-0.265
cc_342 N_A_116_451#_c_352_n N_SCD_c_501_n 0.00171371f $X=1.645 $Y=2.84 $X2=-0.33
+ $Y2=-0.265
cc_343 N_A_116_451#_c_341_n N_SCD_c_501_n 0.0249802f $X=1.73 $Y=2.755 $X2=-0.33
+ $Y2=-0.265
cc_344 N_A_116_451#_c_347_n N_SCD_M1011_g 0.0956367f $X=0.86 $Y=3.115 $X2=0
+ $Y2=0
cc_345 N_A_116_451#_c_351_n N_SCD_M1011_g 0.00157268f $X=0.895 $Y=2.42 $X2=0
+ $Y2=0
cc_346 N_A_116_451#_c_352_n N_SCD_M1011_g 0.0255331f $X=1.645 $Y=2.84 $X2=0
+ $Y2=0
cc_347 N_A_116_451#_c_341_n N_SCD_M1011_g 0.0156407f $X=1.73 $Y=2.755 $X2=0
+ $Y2=0
cc_348 N_A_116_451#_c_354_n N_SCD_M1011_g 0.00217858f $X=2.56 $Y=2.84 $X2=0
+ $Y2=0
cc_349 N_A_116_451#_c_372_p N_SCD_M1011_g 0.00521703f $X=1.73 $Y=2.84 $X2=0
+ $Y2=0
cc_350 N_A_116_451#_c_347_n N_SCD_c_502_n 0.00412465f $X=0.86 $Y=3.115 $X2=0.24
+ $Y2=0
cc_351 N_A_116_451#_c_341_n N_SCD_c_503_n 0.00993f $X=1.73 $Y=2.755 $X2=0.24
+ $Y2=0
cc_352 N_A_116_451#_M1038_g N_SCE_M1016_g 0.0198169f $X=2.71 $Y=0.84 $X2=0 $Y2=0
cc_353 N_A_116_451#_c_341_n N_SCE_M1016_g 2.99507e-19 $X=1.73 $Y=2.755 $X2=0
+ $Y2=0
cc_354 N_A_116_451#_c_342_n N_SCE_M1016_g 0.0229683f $X=2.48 $Y=1.18 $X2=0 $Y2=0
cc_355 N_A_116_451#_c_343_n N_SCE_M1016_g 0.00455662f $X=1.815 $Y=1.18 $X2=0
+ $Y2=0
cc_356 N_A_116_451#_c_339_n N_SCE_c_560_n 0.00394785f $X=2.71 $Y=1.315 $X2=-0.33
+ $Y2=-0.265
cc_357 N_A_116_451#_c_341_n N_SCE_c_560_n 0.00143911f $X=1.73 $Y=2.755 $X2=-0.33
+ $Y2=-0.265
cc_358 N_A_116_451#_c_354_n N_SCE_c_560_n 0.0026244f $X=2.56 $Y=2.84 $X2=-0.33
+ $Y2=-0.265
cc_359 N_A_116_451#_c_355_n N_SCE_c_560_n 0.00749364f $X=2.645 $Y=2.755
+ $X2=-0.33 $Y2=-0.265
cc_360 N_A_116_451#_c_357_n N_SCE_c_560_n 0.00574754f $X=2.73 $Y=2.395 $X2=-0.33
+ $Y2=-0.265
cc_361 N_A_116_451#_c_341_n N_SCE_M1035_g 5.55637e-19 $X=1.73 $Y=2.755 $X2=0
+ $Y2=0
cc_362 N_A_116_451#_c_354_n N_SCE_M1035_g 0.029134f $X=2.56 $Y=2.84 $X2=0 $Y2=0
cc_363 N_A_116_451#_c_355_n N_SCE_M1035_g 0.00401359f $X=2.645 $Y=2.755 $X2=0
+ $Y2=0
cc_364 N_A_116_451#_c_359_n N_SCE_M1014_g 0.0294644f $X=5.155 $Y=2.79 $X2=0.24
+ $Y2=0
cc_365 N_A_116_451#_c_361_n N_SCE_M1014_g 0.0226209f $X=5.32 $Y=3.37 $X2=0.24
+ $Y2=0
cc_366 N_A_116_451#_c_359_n N_SCE_c_567_n 0.00138583f $X=5.155 $Y=2.79 $X2=0
+ $Y2=0
cc_367 N_A_116_451#_c_339_n N_SCE_c_552_n 0.00149363f $X=2.71 $Y=1.315 $X2=0
+ $Y2=0
cc_368 N_A_116_451#_c_341_n N_SCE_c_552_n 0.0264498f $X=1.73 $Y=2.755 $X2=0
+ $Y2=0
cc_369 N_A_116_451#_c_342_n N_SCE_c_552_n 0.0182807f $X=2.48 $Y=1.18 $X2=0 $Y2=0
cc_370 N_A_116_451#_c_393_p N_SCE_c_552_n 0.0119131f $X=2.645 $Y=1.18 $X2=0
+ $Y2=0
cc_371 N_A_116_451#_M1038_g N_SCE_c_553_n 0.0327726f $X=2.71 $Y=0.84 $X2=0 $Y2=0
cc_372 N_A_116_451#_c_341_n N_SCE_c_553_n 0.0171723f $X=1.73 $Y=2.755 $X2=0
+ $Y2=0
cc_373 N_A_116_451#_c_342_n N_SCE_c_553_n 0.00212313f $X=2.48 $Y=1.18 $X2=0
+ $Y2=0
cc_374 N_A_116_451#_c_393_p N_SCE_c_553_n 0.00158394f $X=2.645 $Y=1.18 $X2=0
+ $Y2=0
cc_375 N_A_116_451#_c_341_n N_SCE_c_568_n 0.0416999f $X=1.73 $Y=2.755 $X2=9.6
+ $Y2=0.057
cc_376 N_A_116_451#_c_354_n N_SCE_c_568_n 0.0284833f $X=2.56 $Y=2.84 $X2=9.6
+ $Y2=0.057
cc_377 N_A_116_451#_c_355_n N_SCE_c_568_n 0.00652916f $X=2.645 $Y=2.755 $X2=9.6
+ $Y2=0.057
cc_378 N_A_116_451#_c_357_n N_SCE_c_568_n 0.0131048f $X=2.73 $Y=2.395 $X2=9.6
+ $Y2=0.057
cc_379 N_A_116_451#_c_339_n N_SCE_c_554_n 0.0097199f $X=2.71 $Y=1.315 $X2=0
+ $Y2=0
cc_380 N_A_116_451#_c_342_n N_SCE_c_554_n 0.00315629f $X=2.48 $Y=1.18 $X2=0
+ $Y2=0
cc_381 N_A_116_451#_c_356_n N_SCE_c_554_n 0.0130981f $X=3.385 $Y=2.395 $X2=0
+ $Y2=0
cc_382 N_A_116_451#_c_357_n N_SCE_c_554_n 0.00919594f $X=2.73 $Y=2.395 $X2=0
+ $Y2=0
cc_383 N_A_116_451#_c_344_n N_SCE_c_554_n 0.00647822f $X=5.285 $Y=1.26 $X2=0
+ $Y2=0
cc_384 N_A_116_451#_c_393_p N_SCE_c_554_n 0.0247095f $X=2.645 $Y=1.18 $X2=0
+ $Y2=0
cc_385 N_A_116_451#_c_341_n N_SCE_c_555_n 0.0137116f $X=1.73 $Y=2.755 $X2=0
+ $Y2=0
cc_386 N_A_116_451#_c_342_n N_SCE_c_555_n 0.00490722f $X=2.48 $Y=1.18 $X2=0
+ $Y2=0
cc_387 N_A_116_451#_c_339_n SCE 0.00297688f $X=2.71 $Y=1.315 $X2=0 $Y2=0
cc_388 N_A_116_451#_c_356_n SCE 0.00846076f $X=3.385 $Y=2.395 $X2=0 $Y2=0
cc_389 N_A_116_451#_c_344_n SCE 0.0119984f $X=5.285 $Y=1.26 $X2=0 $Y2=0
cc_390 N_A_116_451#_c_393_p SCE 0.00711763f $X=2.645 $Y=1.18 $X2=0 $Y2=0
cc_391 N_A_116_451#_c_344_n SCE 0.0474159f $X=5.285 $Y=1.26 $X2=0 $Y2=0
cc_392 N_A_116_451#_c_359_n SCE 0.0448683f $X=5.155 $Y=2.79 $X2=0 $Y2=0
cc_393 N_A_116_451#_c_344_n N_SCE_M1012_g 0.0288863f $X=5.285 $Y=1.26 $X2=0
+ $Y2=0
cc_394 N_A_116_451#_c_345_n N_SCE_M1012_g 0.00907758f $X=5.37 $Y=0.84 $X2=0
+ $Y2=0
cc_395 N_A_116_451#_c_356_n N_SCE_c_559_n 0.0130674f $X=3.385 $Y=2.395 $X2=0
+ $Y2=0
cc_396 N_A_116_451#_c_344_n N_SCE_c_559_n 0.108059f $X=5.285 $Y=1.26 $X2=0 $Y2=0
cc_397 N_A_116_451#_c_339_n N_D_c_681_n 0.00184116f $X=2.71 $Y=1.315 $X2=0 $Y2=0
cc_398 N_A_116_451#_c_356_n N_D_c_681_n 0.00860421f $X=3.385 $Y=2.395 $X2=0
+ $Y2=0
cc_399 N_A_116_451#_c_359_n N_D_c_681_n 0.00210555f $X=5.155 $Y=2.79 $X2=0 $Y2=0
cc_400 N_A_116_451#_c_339_n N_D_M1004_g 0.00633826f $X=2.71 $Y=1.315 $X2=0 $Y2=0
cc_401 N_A_116_451#_M1038_g N_D_M1004_g 0.0777906f $X=2.71 $Y=0.84 $X2=0 $Y2=0
cc_402 N_A_116_451#_c_344_n N_D_M1004_g 0.0299403f $X=5.285 $Y=1.26 $X2=0 $Y2=0
cc_403 N_A_116_451#_c_393_p N_D_M1004_g 0.0016937f $X=2.645 $Y=1.18 $X2=0 $Y2=0
cc_404 N_A_116_451#_c_354_n D 0.0136267f $X=2.56 $Y=2.84 $X2=0.24 $Y2=0
cc_405 N_A_116_451#_c_355_n D 0.00674399f $X=2.645 $Y=2.755 $X2=0.24 $Y2=0
cc_406 N_A_116_451#_c_356_n D 0.0210912f $X=3.385 $Y=2.395 $X2=0.24 $Y2=0
cc_407 N_A_116_451#_c_358_n D 0.00317534f $X=3.47 $Y=2.705 $X2=0.24 $Y2=0
cc_408 N_A_116_451#_c_360_n D 0.013626f $X=3.555 $Y=2.79 $X2=0.24 $Y2=0
cc_409 N_A_116_451#_c_354_n N_D_c_683_n 0.00129355f $X=2.56 $Y=2.84 $X2=0 $Y2=0
cc_410 N_A_116_451#_c_355_n N_D_c_683_n 0.00274836f $X=2.645 $Y=2.755 $X2=0
+ $Y2=0
cc_411 N_A_116_451#_c_356_n N_D_c_683_n 0.0330757f $X=3.385 $Y=2.395 $X2=0 $Y2=0
cc_412 N_A_116_451#_c_358_n N_D_c_683_n 0.00326035f $X=3.47 $Y=2.705 $X2=0 $Y2=0
cc_413 N_A_116_451#_c_360_n N_D_c_683_n 0.00163512f $X=3.555 $Y=2.79 $X2=0 $Y2=0
cc_414 N_A_116_451#_c_344_n N_RESET_B_M1024_g 0.0184198f $X=5.285 $Y=1.26 $X2=0
+ $Y2=0
cc_415 N_A_116_451#_c_345_n N_RESET_B_c_1352_n 0.00404708f $X=5.37 $Y=0.84 $X2=0
+ $Y2=0
cc_416 N_A_116_451#_c_358_n N_RESET_B_c_1364_n 0.00408543f $X=3.47 $Y=2.705
+ $X2=18.96 $Y2=0
cc_417 N_A_116_451#_c_359_n N_RESET_B_c_1364_n 0.0425349f $X=5.155 $Y=2.79
+ $X2=18.96 $Y2=0
cc_418 N_A_116_451#_c_344_n N_RESET_B_c_1356_n 0.00960336f $X=5.285 $Y=1.26
+ $X2=0 $Y2=0
cc_419 N_A_116_451#_c_359_n N_RESET_B_c_1365_n 0.0104418f $X=5.155 $Y=2.79 $X2=0
+ $Y2=0
cc_420 N_A_116_451#_c_359_n N_RESET_B_c_1366_n 0.00316724f $X=5.155 $Y=2.79
+ $X2=0 $Y2=0
cc_421 N_A_116_451#_c_359_n N_RESET_B_c_1369_n 0.0257566f $X=5.155 $Y=2.79 $X2=0
+ $Y2=0
cc_422 N_A_116_451#_c_356_n N_RESET_B_c_1358_n 0.00167275f $X=3.385 $Y=2.395
+ $X2=0 $Y2=0
cc_423 N_A_116_451#_c_358_n N_RESET_B_c_1358_n 7.58469e-19 $X=3.47 $Y=2.705
+ $X2=0 $Y2=0
cc_424 N_A_116_451#_c_356_n N_RESET_B_c_1387_n 0.00745183f $X=3.385 $Y=2.395
+ $X2=0 $Y2=0
cc_425 N_A_116_451#_c_358_n N_RESET_B_c_1387_n 0.0017329f $X=3.47 $Y=2.705 $X2=0
+ $Y2=0
cc_426 N_A_116_451#_c_359_n N_RESET_B_c_1387_n 0.0236495f $X=5.155 $Y=2.79 $X2=0
+ $Y2=0
cc_427 N_A_116_451#_c_347_n N_A_65_649#_c_2046_n 0.0261109f $X=0.86 $Y=3.115
+ $X2=18.96 $Y2=0
cc_428 N_A_116_451#_c_351_n N_A_65_649#_c_2046_n 0.0277155f $X=0.895 $Y=2.42
+ $X2=18.96 $Y2=0
cc_429 N_A_116_451#_c_452_p N_A_65_649#_c_2046_n 0.0100032f $X=1.06 $Y=2.84
+ $X2=18.96 $Y2=0
cc_430 N_A_116_451#_M1008_g N_A_65_649#_c_2055_n 0.0118374f $X=0.86 $Y=3.455
+ $X2=0 $Y2=0
cc_431 N_A_116_451#_c_347_n N_A_65_649#_c_2047_n 0.0041515f $X=0.86 $Y=3.115
+ $X2=0 $Y2=0
cc_432 N_A_116_451#_c_351_n N_A_65_649#_c_2047_n 0.0135354f $X=0.895 $Y=2.42
+ $X2=0 $Y2=0
cc_433 N_A_116_451#_c_341_n N_A_65_649#_c_2047_n 0.0130075f $X=1.73 $Y=2.755
+ $X2=0 $Y2=0
cc_434 N_A_116_451#_c_347_n N_A_65_649#_c_2058_n 0.00998495f $X=0.86 $Y=3.115
+ $X2=0 $Y2=0
cc_435 N_A_116_451#_M1008_g N_A_65_649#_c_2058_n 0.0155095f $X=0.86 $Y=3.455
+ $X2=0 $Y2=0
cc_436 N_A_116_451#_c_352_n N_A_65_649#_c_2058_n 0.0378998f $X=1.645 $Y=2.84
+ $X2=0 $Y2=0
cc_437 N_A_116_451#_c_452_p N_A_65_649#_c_2058_n 0.0229739f $X=1.06 $Y=2.84
+ $X2=0 $Y2=0
cc_438 N_A_116_451#_c_354_n N_A_65_649#_c_2058_n 0.0623673f $X=2.56 $Y=2.84
+ $X2=0 $Y2=0
cc_439 N_A_116_451#_c_372_p N_A_65_649#_c_2058_n 0.0117748f $X=1.73 $Y=2.84
+ $X2=0 $Y2=0
cc_440 N_A_116_451#_c_341_n N_A_65_649#_c_2091_n 0.0290194f $X=1.73 $Y=2.755
+ $X2=0 $Y2=0
cc_441 N_A_116_451#_c_343_n N_A_65_649#_c_2091_n 0.0131076f $X=1.815 $Y=1.18
+ $X2=0 $Y2=0
cc_442 N_A_116_451#_M1038_g N_A_65_649#_c_2049_n 0.00857942f $X=2.71 $Y=0.84
+ $X2=0 $Y2=0
cc_443 N_A_116_451#_c_342_n N_A_65_649#_c_2049_n 0.0403313f $X=2.48 $Y=1.18
+ $X2=0 $Y2=0
cc_444 N_A_116_451#_c_343_n N_A_65_649#_c_2049_n 0.0111603f $X=1.815 $Y=1.18
+ $X2=0 $Y2=0
cc_445 N_A_116_451#_c_359_n N_A_65_649#_c_2066_n 0.0919255f $X=5.155 $Y=2.79
+ $X2=0 $Y2=0
cc_446 N_A_116_451#_c_361_n N_A_65_649#_c_2066_n 0.0129587f $X=5.32 $Y=3.37
+ $X2=0 $Y2=0
cc_447 N_A_116_451#_c_360_n N_A_65_649#_c_2067_n 0.0145715f $X=3.555 $Y=2.79
+ $X2=0 $Y2=0
cc_448 N_A_116_451#_c_361_n N_A_65_649#_c_2099_n 0.0155852f $X=5.32 $Y=3.37
+ $X2=0 $Y2=0
cc_449 N_A_116_451#_M1014_d N_A_65_649#_c_2068_n 0.00130674f $X=5.18 $Y=3.245
+ $X2=0 $Y2=0
cc_450 N_A_116_451#_c_361_n N_A_65_649#_c_2068_n 0.019827f $X=5.32 $Y=3.37 $X2=0
+ $Y2=0
cc_451 N_A_116_451#_c_345_n N_A_65_649#_c_2050_n 0.0313963f $X=5.37 $Y=0.84
+ $X2=0 $Y2=0
cc_452 N_A_116_451#_c_361_n N_A_65_649#_c_2074_n 0.0169823f $X=5.32 $Y=3.37
+ $X2=0 $Y2=0
cc_453 N_A_116_451#_c_347_n N_A_65_649#_c_2076_n 0.00370874f $X=0.86 $Y=3.115
+ $X2=0 $Y2=0
cc_454 N_A_116_451#_M1008_g N_A_65_649#_c_2076_n 0.00328219f $X=0.86 $Y=3.455
+ $X2=0 $Y2=0
cc_455 N_A_116_451#_c_344_n N_A_65_649#_c_2053_n 0.00966566f $X=5.285 $Y=1.26
+ $X2=0 $Y2=0
cc_456 N_A_116_451#_c_359_n N_A_65_649#_c_2053_n 0.00869453f $X=5.155 $Y=2.79
+ $X2=0 $Y2=0
cc_457 N_A_116_451#_c_361_n N_A_65_649#_c_2053_n 0.0139058f $X=5.32 $Y=3.37
+ $X2=0 $Y2=0
cc_458 N_A_116_451#_c_345_n N_A_65_649#_c_2053_n 0.00877683f $X=5.37 $Y=0.84
+ $X2=0 $Y2=0
cc_459 N_A_116_451#_M1008_g N_VPWR_c_2199_n 0.00239781f $X=0.86 $Y=3.455 $X2=0
+ $Y2=0
cc_460 N_A_116_451#_M1008_g N_VPWR_c_2220_n 0.017656f $X=0.86 $Y=3.455 $X2=0
+ $Y2=0
cc_461 N_A_116_451#_c_354_n N_VPWR_c_2220_n 6.81464e-19 $X=2.56 $Y=2.84 $X2=0
+ $Y2=0
cc_462 N_A_116_451#_c_359_n N_VPWR_c_2220_n 0.00567298f $X=5.155 $Y=2.79 $X2=0
+ $Y2=0
cc_463 N_A_116_451#_c_360_n N_VPWR_c_2220_n 6.46954e-19 $X=3.555 $Y=2.79 $X2=0
+ $Y2=0
cc_464 N_A_116_451#_c_361_n N_VPWR_c_2220_n 0.0228159f $X=5.32 $Y=3.37 $X2=0
+ $Y2=0
cc_465 N_A_116_451#_M1038_g N_noxref_23_c_2365_n 0.0146952f $X=2.71 $Y=0.84
+ $X2=0.24 $Y2=0
cc_466 N_A_116_451#_c_393_p N_noxref_23_c_2365_n 0.00450421f $X=2.645 $Y=1.18
+ $X2=0.24 $Y2=0
cc_467 N_A_116_451#_M1038_g N_noxref_23_c_2369_n 0.00169006f $X=2.71 $Y=0.84
+ $X2=0 $Y2=0
cc_468 N_A_116_451#_c_344_n N_noxref_23_c_2369_n 0.0199202f $X=5.285 $Y=1.26
+ $X2=0 $Y2=0
cc_469 N_A_116_451#_c_344_n N_VGND_c_2396_n 0.0632635f $X=5.285 $Y=1.26 $X2=0
+ $Y2=0
cc_470 N_A_116_451#_c_345_n N_VGND_c_2396_n 0.0220683f $X=5.37 $Y=0.84 $X2=0
+ $Y2=0
cc_471 N_A_116_451#_M1038_g N_VGND_c_2408_n 0.015669f $X=2.71 $Y=0.84 $X2=0
+ $Y2=0
cc_472 N_A_116_451#_c_342_n N_VGND_c_2408_n 0.00254638f $X=2.48 $Y=1.18 $X2=0
+ $Y2=0
cc_473 N_A_116_451#_c_343_n N_VGND_c_2408_n 7.26677e-19 $X=1.815 $Y=1.18 $X2=0
+ $Y2=0
cc_474 N_A_116_451#_c_344_n N_VGND_c_2408_n 0.0394516f $X=5.285 $Y=1.26 $X2=0
+ $Y2=0
cc_475 N_A_116_451#_c_345_n N_VGND_c_2408_n 0.0238816f $X=5.37 $Y=0.84 $X2=0
+ $Y2=0
cc_476 N_A_116_451#_c_393_p N_VGND_c_2408_n 0.00725212f $X=2.645 $Y=1.18 $X2=0
+ $Y2=0
cc_477 N_SCD_c_500_n N_SCE_M1016_g 0.0427115f $X=1.22 $Y=1.16 $X2=0 $Y2=0
cc_478 N_SCD_c_501_n N_SCE_c_560_n 0.04568f $X=1.22 $Y=1.985 $X2=-0.33
+ $Y2=-0.265
cc_479 N_SCD_M1011_g N_SCE_M1035_g 0.0385464f $X=1.57 $Y=3.455 $X2=0 $Y2=0
cc_480 N_SCD_c_501_n N_SCE_c_553_n 0.00926648f $X=1.22 $Y=1.985 $X2=0 $Y2=0
cc_481 N_SCD_c_503_n N_SCE_c_553_n 0.0427115f $X=1.22 $Y=1.362 $X2=0 $Y2=0
cc_482 N_SCD_c_501_n N_SCE_c_568_n 0.00351783f $X=1.22 $Y=1.985 $X2=9.6
+ $Y2=0.057
cc_483 N_SCD_c_501_n N_A_65_649#_c_2046_n 0.00526067f $X=1.22 $Y=1.985 $X2=18.96
+ $Y2=0
cc_484 N_SCD_M1011_g N_A_65_649#_c_2055_n 0.00168413f $X=1.57 $Y=3.455 $X2=0
+ $Y2=0
cc_485 N_SCD_c_501_n N_A_65_649#_c_2047_n 0.0417103f $X=1.22 $Y=1.985 $X2=0
+ $Y2=0
cc_486 N_SCD_c_502_n N_A_65_649#_c_2047_n 0.00733691f $X=0.97 $Y=1.362 $X2=0
+ $Y2=0
cc_487 N_SCD_c_504_n N_A_65_649#_c_2047_n 0.0454503f $X=0.95 $Y=1.345 $X2=0
+ $Y2=0
cc_488 N_SCD_c_502_n N_A_65_649#_c_2048_n 0.00438532f $X=0.97 $Y=1.362 $X2=9.6
+ $Y2=0.057
cc_489 N_SCD_c_504_n N_A_65_649#_c_2048_n 0.0137314f $X=0.95 $Y=1.345 $X2=9.6
+ $Y2=0.057
cc_490 N_SCD_M1011_g N_A_65_649#_c_2058_n 0.025466f $X=1.57 $Y=3.455 $X2=0 $Y2=0
cc_491 N_SCD_c_500_n N_A_65_649#_c_2091_n 0.0143872f $X=1.22 $Y=1.16 $X2=0 $Y2=0
cc_492 N_SCD_c_501_n N_A_65_649#_c_2091_n 0.00747058f $X=1.22 $Y=1.985 $X2=0
+ $Y2=0
cc_493 N_SCD_c_503_n N_A_65_649#_c_2091_n 0.016295f $X=1.22 $Y=1.362 $X2=0 $Y2=0
cc_494 N_SCD_c_504_n N_A_65_649#_c_2091_n 0.0238596f $X=0.95 $Y=1.345 $X2=0
+ $Y2=0
cc_495 N_SCD_c_500_n N_A_65_649#_c_2122_n 0.0114237f $X=1.22 $Y=1.16 $X2=0 $Y2=0
cc_496 N_SCD_c_500_n N_A_65_649#_c_2049_n 0.00283201f $X=1.22 $Y=1.16 $X2=0
+ $Y2=0
cc_497 N_SCD_M1011_g N_VPWR_c_2199_n 0.0198048f $X=1.57 $Y=3.455 $X2=0 $Y2=0
cc_498 N_SCD_M1011_g N_VPWR_c_2220_n 0.011273f $X=1.57 $Y=3.455 $X2=0 $Y2=0
cc_499 N_SCD_c_500_n N_noxref_23_c_2364_n 0.0143864f $X=1.22 $Y=1.16 $X2=0 $Y2=0
cc_500 N_SCD_c_502_n N_noxref_23_c_2364_n 0.00728568f $X=0.97 $Y=1.362 $X2=0
+ $Y2=0
cc_501 N_SCD_c_504_n N_noxref_23_c_2364_n 0.0220358f $X=0.95 $Y=1.345 $X2=0
+ $Y2=0
cc_502 N_SCD_c_500_n N_noxref_23_c_2365_n 0.0146562f $X=1.22 $Y=1.16 $X2=0.24
+ $Y2=0
cc_503 N_SCD_c_500_n N_VGND_c_2408_n 0.0165804f $X=1.22 $Y=1.16 $X2=0 $Y2=0
cc_504 N_SCD_c_502_n N_VGND_c_2408_n 0.0129994f $X=0.97 $Y=1.362 $X2=0 $Y2=0
cc_505 N_SCD_c_504_n N_VGND_c_2408_n 0.0233861f $X=0.95 $Y=1.345 $X2=0 $Y2=0
cc_506 N_SCE_c_560_n N_D_c_681_n 0.0543283f $X=2.37 $Y=2.675 $X2=0 $Y2=0
cc_507 N_SCE_c_568_n N_D_c_681_n 6.30109e-19 $X=2.215 $Y=2.15 $X2=0 $Y2=0
cc_508 N_SCE_c_554_n N_D_c_681_n 0.00293558f $X=3.005 $Y=1.92 $X2=0 $Y2=0
cc_509 SCE N_D_c_681_n 0.00473256f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_510 N_SCE_c_554_n N_D_M1004_g 8.29566e-19 $X=3.005 $Y=1.92 $X2=0 $Y2=0
cc_511 SCE N_D_M1004_g 0.0144117f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_512 N_SCE_c_559_n N_D_M1004_g 0.038843f $X=4.88 $Y=1.692 $X2=0 $Y2=0
cc_513 N_SCE_c_560_n D 2.37558e-19 $X=2.37 $Y=2.675 $X2=0.24 $Y2=0
cc_514 N_SCE_M1035_g D 0.00124877f $X=2.37 $Y=3.455 $X2=0.24 $Y2=0
cc_515 N_SCE_M1035_g N_D_c_683_n 0.0543283f $X=2.37 $Y=3.455 $X2=0 $Y2=0
cc_516 N_SCE_M1014_g N_RESET_B_M1019_g 0.0108857f $X=4.93 $Y=3.455 $X2=0 $Y2=0
cc_517 N_SCE_M1012_g N_RESET_B_M1024_g 0.0360909f $X=4.98 $Y=0.84 $X2=0 $Y2=0
cc_518 N_SCE_M1012_g N_RESET_B_c_1352_n 0.034112f $X=4.98 $Y=0.84 $X2=0 $Y2=0
cc_519 N_SCE_M1014_g N_RESET_B_c_1364_n 0.021247f $X=4.93 $Y=3.455 $X2=18.96
+ $Y2=0
cc_520 N_SCE_c_559_n N_RESET_B_c_1356_n 0.0112649f $X=4.88 $Y=1.692 $X2=0 $Y2=0
cc_521 N_SCE_c_567_n N_RESET_B_c_1365_n 0.0039871f $X=4.955 $Y=2.545 $X2=0 $Y2=0
cc_522 SCE N_RESET_B_c_1365_n 0.0686615f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_523 N_SCE_c_559_n N_RESET_B_c_1365_n 0.00495303f $X=4.88 $Y=1.692 $X2=0 $Y2=0
cc_524 N_SCE_c_567_n N_RESET_B_c_1366_n 0.0022337f $X=4.955 $Y=2.545 $X2=0 $Y2=0
cc_525 SCE N_RESET_B_c_1366_n 0.00230712f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_526 N_SCE_c_559_n N_RESET_B_c_1366_n 0.00714324f $X=4.88 $Y=1.692 $X2=0 $Y2=0
cc_527 N_SCE_c_567_n N_RESET_B_c_1369_n 0.00225016f $X=4.955 $Y=2.545 $X2=0
+ $Y2=0
cc_528 SCE N_RESET_B_c_1369_n 0.0133949f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_529 N_SCE_c_559_n N_RESET_B_c_1369_n 0.011092f $X=4.88 $Y=1.692 $X2=0 $Y2=0
cc_530 N_SCE_c_567_n N_RESET_B_c_1358_n 0.021247f $X=4.955 $Y=2.545 $X2=0 $Y2=0
cc_531 SCE N_RESET_B_c_1358_n 0.00206317f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_532 N_SCE_M1012_g N_RESET_B_c_1358_n 0.0147161f $X=4.98 $Y=0.84 $X2=0 $Y2=0
cc_533 N_SCE_c_559_n N_RESET_B_c_1358_n 0.0227586f $X=4.88 $Y=1.692 $X2=0 $Y2=0
cc_534 N_SCE_c_567_n N_RESET_B_c_1387_n 0.00116218f $X=4.955 $Y=2.545 $X2=0
+ $Y2=0
cc_535 SCE N_RESET_B_c_1387_n 0.00797999f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_536 N_SCE_c_559_n N_RESET_B_c_1387_n 0.0245438f $X=4.88 $Y=1.692 $X2=0 $Y2=0
cc_537 N_SCE_M1035_g N_A_65_649#_c_2058_n 0.0240499f $X=2.37 $Y=3.455 $X2=0
+ $Y2=0
cc_538 N_SCE_M1016_g N_A_65_649#_c_2091_n 0.00201788f $X=1.93 $Y=0.84 $X2=0
+ $Y2=0
cc_539 N_SCE_M1016_g N_A_65_649#_c_2049_n 0.0263564f $X=1.93 $Y=0.84 $X2=0 $Y2=0
cc_540 N_SCE_M1035_g N_A_65_649#_c_2127_n 0.0105058f $X=2.37 $Y=3.455 $X2=0
+ $Y2=0
cc_541 N_SCE_M1035_g N_A_65_649#_c_2062_n 0.00424052f $X=2.37 $Y=3.455 $X2=0
+ $Y2=0
cc_542 N_SCE_M1014_g N_A_65_649#_c_2066_n 0.0163883f $X=4.93 $Y=3.455 $X2=0
+ $Y2=0
cc_543 N_SCE_M1014_g N_A_65_649#_c_2099_n 0.017945f $X=4.93 $Y=3.455 $X2=0 $Y2=0
cc_544 N_SCE_M1014_g N_A_65_649#_c_2068_n 0.0143804f $X=4.93 $Y=3.455 $X2=0
+ $Y2=0
cc_545 N_SCE_M1014_g N_A_65_649#_c_2071_n 0.00702623f $X=4.93 $Y=3.455 $X2=0
+ $Y2=0
cc_546 N_SCE_M1014_g N_A_65_649#_c_2074_n 6.61814e-19 $X=4.93 $Y=3.455 $X2=0
+ $Y2=0
cc_547 N_SCE_M1014_g N_A_65_649#_c_2075_n 0.00179017f $X=4.93 $Y=3.455 $X2=0
+ $Y2=0
cc_548 N_SCE_M1014_g N_A_65_649#_c_2053_n 0.00546712f $X=4.93 $Y=3.455 $X2=0
+ $Y2=0
cc_549 N_SCE_c_567_n N_A_65_649#_c_2053_n 5.10276e-19 $X=4.955 $Y=2.545 $X2=0
+ $Y2=0
cc_550 SCE N_A_65_649#_c_2053_n 0.0712561f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_551 N_SCE_M1012_g N_A_65_649#_c_2053_n 0.00899417f $X=4.98 $Y=0.84 $X2=0
+ $Y2=0
cc_552 N_SCE_M1035_g N_VPWR_c_2199_n 0.011721f $X=2.37 $Y=3.455 $X2=0 $Y2=0
cc_553 N_SCE_M1014_g N_VPWR_c_2202_n 0.00279807f $X=4.93 $Y=3.455 $X2=0 $Y2=0
cc_554 N_SCE_M1035_g N_VPWR_c_2220_n 0.00942952f $X=2.37 $Y=3.455 $X2=0 $Y2=0
cc_555 N_SCE_M1014_g N_VPWR_c_2220_n 0.0100282f $X=4.93 $Y=3.455 $X2=0 $Y2=0
cc_556 N_SCE_M1016_g N_noxref_23_c_2364_n 6.66769e-19 $X=1.93 $Y=0.84 $X2=0
+ $Y2=0
cc_557 N_SCE_M1016_g N_noxref_23_c_2365_n 0.0110269f $X=1.93 $Y=0.84 $X2=0.24
+ $Y2=0
cc_558 N_SCE_M1012_g N_VGND_c_2396_n 0.0306975f $X=4.98 $Y=0.84 $X2=0 $Y2=0
cc_559 N_SCE_M1016_g N_VGND_c_2408_n 0.00724706f $X=1.93 $Y=0.84 $X2=0 $Y2=0
cc_560 N_SCE_M1012_g N_VGND_c_2408_n 0.00463336f $X=4.98 $Y=0.84 $X2=0 $Y2=0
cc_561 N_D_M1004_g N_RESET_B_M1024_g 0.0371745f $X=3.42 $Y=0.84 $X2=0 $Y2=0
cc_562 N_D_c_681_n N_RESET_B_c_1364_n 0.00409093f $X=3.42 $Y=2.175 $X2=18.96
+ $Y2=0
cc_563 D N_RESET_B_c_1364_n 0.00131501f $X=3.035 $Y=2.69 $X2=18.96 $Y2=0
cc_564 N_D_c_683_n N_RESET_B_c_1364_n 0.040721f $X=3.06 $Y=2.825 $X2=18.96 $Y2=0
cc_565 N_D_c_681_n N_RESET_B_c_1356_n 0.0371745f $X=3.42 $Y=2.175 $X2=0 $Y2=0
cc_566 N_D_c_683_n N_RESET_B_c_1358_n 0.00325217f $X=3.06 $Y=2.825 $X2=0 $Y2=0
cc_567 N_D_M1004_g N_RESET_B_c_1387_n 0.00203633f $X=3.42 $Y=0.84 $X2=0 $Y2=0
cc_568 D N_A_65_649#_c_2058_n 0.0123978f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_569 N_D_c_683_n N_A_65_649#_c_2058_n 0.00140466f $X=3.06 $Y=2.825 $X2=0 $Y2=0
cc_570 N_D_M1004_g N_A_65_649#_c_2049_n 9.1669e-19 $X=3.42 $Y=0.84 $X2=0 $Y2=0
cc_571 N_D_c_683_n N_A_65_649#_c_2127_n 0.00285181f $X=3.06 $Y=2.825 $X2=0 $Y2=0
cc_572 D N_A_65_649#_c_2059_n 0.0108958f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_573 N_D_c_683_n N_A_65_649#_c_2059_n 0.0210703f $X=3.06 $Y=2.825 $X2=0 $Y2=0
cc_574 D N_A_65_649#_c_2065_n 0.00188352f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_575 N_D_c_683_n N_A_65_649#_c_2065_n 5.74689e-19 $X=3.06 $Y=2.825 $X2=0 $Y2=0
cc_576 D N_A_65_649#_c_2067_n 0.013626f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_577 N_D_c_683_n N_A_65_649#_c_2067_n 0.00163512f $X=3.06 $Y=2.825 $X2=0 $Y2=0
cc_578 N_D_c_683_n N_VPWR_c_2199_n 2.17204e-19 $X=3.06 $Y=2.825 $X2=0 $Y2=0
cc_579 D N_VPWR_c_2220_n 0.00804915f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_580 N_D_c_683_n N_VPWR_c_2220_n 0.0177209f $X=3.06 $Y=2.825 $X2=0 $Y2=0
cc_581 N_D_M1004_g N_noxref_23_c_2365_n 0.0171077f $X=3.42 $Y=0.84 $X2=0.24
+ $Y2=0
cc_582 N_D_M1004_g N_noxref_23_c_2369_n 0.0146315f $X=3.42 $Y=0.84 $X2=0 $Y2=0
cc_583 N_D_M1004_g N_VGND_c_2396_n 2.15619e-19 $X=3.42 $Y=0.84 $X2=0 $Y2=0
cc_584 N_D_M1004_g N_VGND_c_2408_n 0.0150913f $X=3.42 $Y=0.84 $X2=0 $Y2=0
cc_585 N_A_1212_471#_c_738_n N_A_1212_100#_M1022_g 0.0569691f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_586 N_A_1212_471#_c_739_n N_A_1212_100#_M1022_g 0.00367584f $X=7.045 $Y=0.35
+ $X2=0 $Y2=0
cc_587 N_A_1212_471#_c_743_n N_A_1212_100#_M1022_g 0.00100082f $X=7.15 $Y=1.175
+ $X2=0 $Y2=0
cc_588 N_A_1212_471#_c_744_n N_A_1212_100#_M1022_g 3.11135e-19 $X=7.15 $Y=1.57
+ $X2=0 $Y2=0
cc_589 N_A_1212_471#_M1001_g N_A_1212_100#_M1022_g 0.0385598f $X=7.09 $Y=0.84
+ $X2=0 $Y2=0
cc_590 N_A_1212_471#_c_738_n N_A_1212_100#_c_1004_n 0.00831103f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_591 N_A_1212_471#_c_750_n N_A_1212_100#_c_1004_n 0.031f $X=6.27 $Y=2.54 $X2=0
+ $Y2=0
cc_592 N_A_1212_471#_c_750_n N_A_1212_100#_c_1005_n 0.0157004f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_593 N_A_1212_471#_c_744_n N_A_1212_100#_c_1005_n 2.41421e-19 $X=7.15 $Y=1.57
+ $X2=0 $Y2=0
cc_594 N_A_1212_471#_M1001_g N_A_1212_100#_c_1005_n 0.0332258f $X=7.09 $Y=0.84
+ $X2=0 $Y2=0
cc_595 N_A_1212_471#_c_738_n N_A_1212_100#_M1003_g 0.0014021f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_596 N_A_1212_471#_c_750_n N_A_1212_100#_M1003_g 0.0360406f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_597 N_A_1212_471#_c_753_n N_A_1212_100#_M1003_g 0.0170833f $X=7.045 $Y=3.72
+ $X2=0 $Y2=0
cc_598 N_A_1212_471#_c_786_p N_A_1212_100#_M1003_g 0.0165468f $X=7.13 $Y=3.635
+ $X2=0 $Y2=0
cc_599 N_A_1212_471#_c_759_n N_A_1212_100#_M1003_g 0.00714723f $X=8.535 $Y=3.15
+ $X2=0 $Y2=0
cc_600 N_A_1212_471#_c_788_p N_A_1212_100#_M1003_g 0.00766182f $X=7.215 $Y=3.15
+ $X2=0 $Y2=0
cc_601 N_A_1212_471#_c_746_n N_A_1212_100#_c_977_n 0.0101838f $X=9.47 $Y=1.115
+ $X2=18.96 $Y2=0
cc_602 N_A_1212_471#_c_745_n N_A_1212_100#_c_978_n 0.00218131f $X=9.305 $Y=1.26
+ $X2=0 $Y2=0
cc_603 N_A_1212_471#_c_766_n N_A_1212_100#_c_978_n 0.00959677f $X=9.62 $Y=2.86
+ $X2=0 $Y2=0
cc_604 N_A_1212_471#_c_746_n N_A_1212_100#_c_978_n 0.00906084f $X=9.47 $Y=1.115
+ $X2=0 $Y2=0
cc_605 N_A_1212_471#_c_766_n N_A_1212_100#_M1020_g 0.0228703f $X=9.62 $Y=2.86
+ $X2=0 $Y2=0
cc_606 N_A_1212_471#_c_767_n N_A_1212_100#_M1020_g 0.0117163f $X=9.62 $Y=3.635
+ $X2=0 $Y2=0
cc_607 N_A_1212_471#_c_795_p N_A_1212_100#_M1020_g 0.0374019f $X=11.62 $Y=3.22
+ $X2=0 $Y2=0
cc_608 N_A_1212_471#_c_771_n N_A_1212_100#_M1020_g 3.84191e-19 $X=9.62 $Y=3.22
+ $X2=0 $Y2=0
cc_609 N_A_1212_471#_c_795_p N_A_1212_100#_c_1013_n 0.0164437f $X=11.62 $Y=3.22
+ $X2=0 $Y2=0
cc_610 N_A_1212_471#_c_798_p N_A_1212_100#_c_1013_n 0.0222007f $X=11.705
+ $Y=3.135 $X2=0 $Y2=0
cc_611 N_A_1212_471#_c_769_n N_A_1212_100#_c_1013_n 0.0123959f $X=12.48 $Y=3.22
+ $X2=0 $Y2=0
cc_612 N_A_1212_471#_c_800_p N_A_1212_100#_c_1013_n 0.00103903f $X=12.645
+ $Y=2.39 $X2=0 $Y2=0
cc_613 N_A_1212_471#_c_770_n N_A_1212_100#_c_1013_n 0.0149132f $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_614 N_A_1212_471#_c_802_p N_A_1212_100#_c_1013_n 0.00555541f $X=11.705
+ $Y=3.22 $X2=0 $Y2=0
cc_615 N_A_1212_471#_c_737_n N_A_1212_100#_c_979_n 0.0215974f $X=11.55 $Y=1.445
+ $X2=0 $Y2=0
cc_616 N_A_1212_471#_c_768_n N_A_1212_100#_c_979_n 0.00273438f $X=11.395 $Y=1.63
+ $X2=0 $Y2=0
cc_617 N_A_1212_471#_c_798_p N_A_1212_100#_c_979_n 0.00669732f $X=11.705
+ $Y=3.135 $X2=0 $Y2=0
cc_618 N_A_1212_471#_c_769_n N_A_1212_100#_c_979_n 6.25698e-19 $X=12.48 $Y=3.22
+ $X2=0 $Y2=0
cc_619 N_A_1212_471#_c_800_p N_A_1212_100#_c_979_n 3.25741e-19 $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_620 N_A_1212_471#_c_770_n N_A_1212_100#_c_979_n 0.0325075f $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_621 N_A_1212_471#_c_772_n N_A_1212_100#_c_979_n 0.013315f $X=11.705 $Y=2.37
+ $X2=0 $Y2=0
cc_622 N_A_1212_471#_c_737_n N_A_1212_100#_M1000_g 0.0121851f $X=11.55 $Y=1.445
+ $X2=0 $Y2=0
cc_623 N_A_1212_471#_c_750_n N_A_1212_100#_c_1062_n 2.1042e-19 $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_624 N_A_1212_471#_c_744_n N_A_1212_100#_c_981_n 0.00274704f $X=7.15 $Y=1.57
+ $X2=0 $Y2=0
cc_625 N_A_1212_471#_M1001_g N_A_1212_100#_c_981_n 2.62551e-19 $X=7.09 $Y=0.84
+ $X2=0 $Y2=0
cc_626 N_A_1212_471#_c_745_n N_A_1212_100#_c_982_n 0.114334f $X=9.305 $Y=1.26
+ $X2=0 $Y2=0
cc_627 N_A_1212_471#_c_746_n N_A_1212_100#_c_982_n 0.0244077f $X=9.47 $Y=1.115
+ $X2=0 $Y2=0
cc_628 N_A_1212_471#_c_744_n N_A_1212_100#_c_983_n 0.013321f $X=7.15 $Y=1.57
+ $X2=0 $Y2=0
cc_629 N_A_1212_471#_c_745_n N_A_1212_100#_c_983_n 0.0127422f $X=9.305 $Y=1.26
+ $X2=0 $Y2=0
cc_630 N_A_1212_471#_M1001_g N_A_1212_100#_c_983_n 0.00130695f $X=7.09 $Y=0.84
+ $X2=0 $Y2=0
cc_631 N_A_1212_471#_c_737_n N_A_1212_100#_c_1070_n 0.00117255f $X=11.55
+ $Y=1.445 $X2=0 $Y2=0
cc_632 N_A_1212_471#_c_737_n N_A_1212_100#_c_984_n 0.0173691f $X=11.55 $Y=1.445
+ $X2=0 $Y2=0
cc_633 N_A_1212_471#_c_737_n N_A_1212_100#_c_988_n 2.42178e-19 $X=11.55 $Y=1.445
+ $X2=0 $Y2=0
cc_634 N_A_1212_471#_c_737_n N_A_1212_100#_c_989_n 0.0028884f $X=11.55 $Y=1.445
+ $X2=0 $Y2=0
cc_635 N_A_1212_471#_c_744_n N_A_1212_100#_c_1023_n 0.015439f $X=7.15 $Y=1.57
+ $X2=0 $Y2=0
cc_636 N_A_1212_471#_c_745_n N_A_1212_100#_c_1023_n 0.00552447f $X=9.305 $Y=1.26
+ $X2=0 $Y2=0
cc_637 N_A_1212_471#_M1001_g N_A_1212_100#_c_1023_n 0.00357027f $X=7.09 $Y=0.84
+ $X2=0 $Y2=0
cc_638 N_A_1212_471#_c_737_n N_A_1212_100#_c_1000_n 0.0316057f $X=11.55 $Y=1.445
+ $X2=0 $Y2=0
cc_639 N_A_1212_471#_c_770_n N_A_1212_100#_c_1000_n 0.0230135f $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_640 N_A_1212_471#_c_795_p N_A_1510_100#_M1009_d 0.00390627f $X=11.62 $Y=3.22
+ $X2=0 $Y2=0
cc_641 N_A_1212_471#_c_743_n N_A_1510_100#_M1010_g 0.00450474f $X=7.15 $Y=1.175
+ $X2=0 $Y2=0
cc_642 N_A_1212_471#_c_744_n N_A_1510_100#_M1010_g 0.00128775f $X=7.15 $Y=1.57
+ $X2=0 $Y2=0
cc_643 N_A_1212_471#_c_745_n N_A_1510_100#_M1010_g 0.0292526f $X=9.305 $Y=1.26
+ $X2=0 $Y2=0
cc_644 N_A_1212_471#_M1001_g N_A_1510_100#_M1010_g 0.0868283f $X=7.09 $Y=0.84
+ $X2=0 $Y2=0
cc_645 N_A_1212_471#_c_753_n N_A_1510_100#_M1015_g 5.61619e-19 $X=7.045 $Y=3.72
+ $X2=0 $Y2=0
cc_646 N_A_1212_471#_c_786_p N_A_1510_100#_M1015_g 0.00127662f $X=7.13 $Y=3.635
+ $X2=0 $Y2=0
cc_647 N_A_1212_471#_c_759_n N_A_1510_100#_M1015_g 0.0257143f $X=8.535 $Y=3.15
+ $X2=0 $Y2=0
cc_648 N_A_1212_471#_c_836_p N_A_1510_100#_M1015_g 7.57207e-19 $X=8.62 $Y=3.635
+ $X2=0 $Y2=0
cc_649 N_A_1212_471#_c_763_n N_A_1510_100#_M1015_g 4.59593e-19 $X=8.705 $Y=3.72
+ $X2=0 $Y2=0
cc_650 N_A_1212_471#_c_737_n N_A_1510_100#_c_1267_n 0.0124309f $X=11.55 $Y=1.445
+ $X2=9.6 $Y2=0
cc_651 N_A_1212_471#_c_737_n N_A_1510_100#_c_1247_n 0.00441813f $X=11.55
+ $Y=1.445 $X2=0 $Y2=0
cc_652 N_A_1212_471#_c_768_n N_A_1510_100#_c_1247_n 0.0280532f $X=11.395 $Y=1.63
+ $X2=0 $Y2=0
cc_653 N_A_1212_471#_c_737_n N_A_1510_100#_c_1253_n 6.64643e-19 $X=11.55
+ $Y=1.445 $X2=0 $Y2=0
cc_654 N_A_1212_471#_c_768_n N_A_1510_100#_c_1253_n 0.0169593f $X=11.395 $Y=1.63
+ $X2=0 $Y2=0
cc_655 N_A_1212_471#_c_798_p N_A_1510_100#_c_1253_n 0.00601479f $X=11.705
+ $Y=3.135 $X2=0 $Y2=0
cc_656 N_A_1212_471#_c_772_n N_A_1510_100#_c_1253_n 0.0116702f $X=11.705 $Y=2.37
+ $X2=0 $Y2=0
cc_657 N_A_1212_471#_c_737_n N_A_1510_100#_c_1274_n 0.00684719f $X=11.55
+ $Y=1.445 $X2=0 $Y2=0
cc_658 N_A_1212_471#_c_768_n N_A_1510_100#_c_1274_n 0.0010494f $X=11.395 $Y=1.63
+ $X2=0 $Y2=0
cc_659 N_A_1212_471#_c_737_n N_A_1510_100#_c_1255_n 0.00134037f $X=11.55
+ $Y=1.445 $X2=0 $Y2=0
cc_660 N_A_1212_471#_c_768_n N_A_1510_100#_c_1255_n 0.0131385f $X=11.395 $Y=1.63
+ $X2=0 $Y2=0
cc_661 N_A_1212_471#_c_737_n N_A_1510_100#_c_1256_n 0.00239177f $X=11.55
+ $Y=1.445 $X2=0 $Y2=0
cc_662 N_A_1212_471#_c_795_p N_A_1510_100#_c_1256_n 0.0242527f $X=11.62 $Y=3.22
+ $X2=0 $Y2=0
cc_663 N_A_1212_471#_c_798_p N_A_1510_100#_c_1256_n 0.0196451f $X=11.705
+ $Y=3.135 $X2=0 $Y2=0
cc_664 N_A_1212_471#_c_772_n N_A_1510_100#_c_1256_n 0.00665983f $X=11.705
+ $Y=2.37 $X2=0 $Y2=0
cc_665 N_A_1212_471#_c_739_n N_RESET_B_c_1352_n 0.0159638f $X=7.045 $Y=0.35
+ $X2=0 $Y2=0
cc_666 N_A_1212_471#_c_741_n N_RESET_B_c_1352_n 0.00333865f $X=6.355 $Y=0.35
+ $X2=0 $Y2=0
cc_667 N_A_1212_471#_M1001_g N_RESET_B_c_1352_n 0.0337051f $X=7.09 $Y=0.84 $X2=0
+ $Y2=0
cc_668 N_A_1212_471#_c_746_n N_RESET_B_M1013_g 0.00288781f $X=9.47 $Y=1.115
+ $X2=0 $Y2=0
cc_669 N_A_1212_471#_c_745_n N_RESET_B_c_1357_n 0.0320286f $X=9.305 $Y=1.26
+ $X2=0 $Y2=0
cc_670 N_A_1212_471#_c_746_n N_RESET_B_c_1357_n 0.00132414f $X=9.47 $Y=1.115
+ $X2=0 $Y2=0
cc_671 N_A_1212_471#_c_738_n N_RESET_B_c_1365_n 0.0188f $X=6.27 $Y=2.54 $X2=0
+ $Y2=0
cc_672 N_A_1212_471#_c_750_n N_RESET_B_c_1365_n 0.0146417f $X=6.27 $Y=2.54 $X2=0
+ $Y2=0
cc_673 N_A_1212_471#_M1001_g N_RESET_B_c_1365_n 4.28754e-19 $X=7.09 $Y=0.84
+ $X2=0 $Y2=0
cc_674 N_A_1212_471#_c_737_n N_RESET_B_c_1367_n 0.00220001f $X=11.55 $Y=1.445
+ $X2=0 $Y2=0
cc_675 N_A_1212_471#_c_766_n N_RESET_B_c_1367_n 0.00766432f $X=9.62 $Y=2.86
+ $X2=0 $Y2=0
cc_676 N_A_1212_471#_c_768_n N_RESET_B_c_1367_n 0.00178896f $X=11.395 $Y=1.63
+ $X2=0 $Y2=0
cc_677 N_A_1212_471#_c_798_p N_RESET_B_c_1367_n 0.0099513f $X=11.705 $Y=3.135
+ $X2=0 $Y2=0
cc_678 N_A_1212_471#_c_800_p N_RESET_B_c_1367_n 0.0294764f $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_679 N_A_1212_471#_c_770_n N_RESET_B_c_1367_n 0.00990881f $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_680 N_A_1212_471#_c_772_n N_RESET_B_c_1367_n 0.0188276f $X=11.705 $Y=2.37
+ $X2=0 $Y2=0
cc_681 N_A_1212_471#_c_759_n N_RESET_B_c_1359_n 0.0158362f $X=8.535 $Y=3.15
+ $X2=0 $Y2=0
cc_682 N_A_1212_471#_c_836_p N_RESET_B_c_1359_n 0.0170271f $X=8.62 $Y=3.635
+ $X2=0 $Y2=0
cc_683 N_A_1212_471#_c_760_n N_RESET_B_c_1359_n 0.0128285f $X=9.455 $Y=3.72
+ $X2=0 $Y2=0
cc_684 N_A_1212_471#_c_763_n N_RESET_B_c_1359_n 0.00579092f $X=8.705 $Y=3.72
+ $X2=0 $Y2=0
cc_685 N_A_1212_471#_c_766_n N_RESET_B_c_1359_n 0.00163271f $X=9.62 $Y=2.86
+ $X2=0 $Y2=0
cc_686 N_A_1212_471#_c_767_n N_RESET_B_c_1359_n 0.00209476f $X=9.62 $Y=3.635
+ $X2=0 $Y2=0
cc_687 N_A_1212_471#_c_771_n N_RESET_B_c_1359_n 5.06755e-19 $X=9.62 $Y=3.22
+ $X2=0 $Y2=0
cc_688 N_A_1212_471#_c_737_n N_A_1312_126#_M1007_g 0.0500283f $X=11.55 $Y=1.445
+ $X2=0 $Y2=0
cc_689 N_A_1212_471#_c_768_n N_A_1312_126#_M1007_g 4.41214e-19 $X=11.395 $Y=1.63
+ $X2=0 $Y2=0
cc_690 N_A_1212_471#_c_737_n N_A_1312_126#_c_1562_n 0.00874305f $X=11.55
+ $Y=1.445 $X2=0 $Y2=0
cc_691 N_A_1212_471#_c_795_p N_A_1312_126#_c_1562_n 0.0369003f $X=11.62 $Y=3.22
+ $X2=0 $Y2=0
cc_692 N_A_1212_471#_c_768_n N_A_1312_126#_c_1562_n 8.48736e-19 $X=11.395
+ $Y=1.63 $X2=0 $Y2=0
cc_693 N_A_1212_471#_c_798_p N_A_1312_126#_c_1562_n 0.00141636f $X=11.705
+ $Y=3.135 $X2=0 $Y2=0
cc_694 N_A_1212_471#_c_772_n N_A_1312_126#_c_1562_n 8.61122e-19 $X=11.705
+ $Y=2.37 $X2=0 $Y2=0
cc_695 N_A_1212_471#_c_738_n N_A_1312_126#_c_1563_n 0.112506f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_696 N_A_1212_471#_c_750_n N_A_1312_126#_c_1563_n 0.00773145f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_697 N_A_1212_471#_c_743_n N_A_1312_126#_c_1563_n 0.00769944f $X=7.15 $Y=1.175
+ $X2=0 $Y2=0
cc_698 N_A_1212_471#_c_744_n N_A_1312_126#_c_1563_n 0.0168768f $X=7.15 $Y=1.57
+ $X2=0 $Y2=0
cc_699 N_A_1212_471#_c_887_p N_A_1312_126#_c_1563_n 0.00805772f $X=7.15 $Y=1.26
+ $X2=0 $Y2=0
cc_700 N_A_1212_471#_M1001_g N_A_1312_126#_c_1563_n 0.00646356f $X=7.09 $Y=0.84
+ $X2=0 $Y2=0
cc_701 N_A_1212_471#_c_738_n N_A_1312_126#_c_1589_n 0.0387742f $X=6.27 $Y=2.54
+ $X2=9.6 $Y2=0
cc_702 N_A_1212_471#_c_750_n N_A_1312_126#_c_1589_n 0.0134172f $X=6.27 $Y=2.54
+ $X2=9.6 $Y2=0
cc_703 N_A_1212_471#_c_753_n N_A_1312_126#_c_1589_n 0.0199321f $X=7.045 $Y=3.72
+ $X2=9.6 $Y2=0
cc_704 N_A_1212_471#_c_786_p N_A_1312_126#_c_1589_n 0.014903f $X=7.13 $Y=3.635
+ $X2=9.6 $Y2=0
cc_705 N_A_1212_471#_c_788_p N_A_1312_126#_c_1589_n 0.0129587f $X=7.215 $Y=3.15
+ $X2=9.6 $Y2=0
cc_706 N_A_1212_471#_c_759_n N_A_1312_126#_c_1569_n 0.0955579f $X=8.535 $Y=3.15
+ $X2=9.6 $Y2=0.057
cc_707 N_A_1212_471#_c_788_p N_A_1312_126#_c_1569_n 0.011601f $X=7.215 $Y=3.15
+ $X2=9.6 $Y2=0.057
cc_708 N_A_1212_471#_c_759_n N_A_1312_126#_c_1570_n 0.0129587f $X=8.535 $Y=3.15
+ $X2=0 $Y2=0
cc_709 N_A_1212_471#_c_836_p N_A_1312_126#_c_1570_n 0.014903f $X=8.62 $Y=3.635
+ $X2=0 $Y2=0
cc_710 N_A_1212_471#_c_760_n N_A_1312_126#_c_1570_n 0.0209781f $X=9.455 $Y=3.72
+ $X2=0 $Y2=0
cc_711 N_A_1212_471#_c_766_n N_A_1312_126#_c_1570_n 0.0163009f $X=9.62 $Y=2.86
+ $X2=0 $Y2=0
cc_712 N_A_1212_471#_c_767_n N_A_1312_126#_c_1570_n 0.00964628f $X=9.62 $Y=3.635
+ $X2=0 $Y2=0
cc_713 N_A_1212_471#_c_771_n N_A_1312_126#_c_1570_n 0.0118078f $X=9.62 $Y=3.22
+ $X2=0 $Y2=0
cc_714 N_A_1212_471#_c_766_n N_A_1312_126#_c_1571_n 0.00121706f $X=9.62 $Y=2.86
+ $X2=0 $Y2=0
cc_715 N_A_1212_471#_c_766_n N_A_1312_126#_c_1572_n 0.0120276f $X=9.62 $Y=2.86
+ $X2=0 $Y2=0
cc_716 N_A_1212_471#_c_738_n N_A_1312_126#_c_1564_n 0.0258485f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_717 N_A_1212_471#_c_739_n N_A_1312_126#_c_1564_n 0.0220953f $X=7.045 $Y=0.35
+ $X2=0 $Y2=0
cc_718 N_A_1212_471#_c_743_n N_A_1312_126#_c_1564_n 0.0262454f $X=7.15 $Y=1.175
+ $X2=0 $Y2=0
cc_719 N_A_1212_471#_M1001_g N_A_1312_126#_c_1564_n 0.00800283f $X=7.09 $Y=0.84
+ $X2=0 $Y2=0
cc_720 N_A_1212_471#_c_738_n N_A_1312_126#_c_1574_n 0.0123662f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_721 N_A_1212_471#_c_750_n N_A_1312_126#_c_1574_n 0.00495995f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_722 N_A_1212_471#_c_766_n N_A_1312_126#_c_1575_n 0.0118078f $X=9.62 $Y=2.86
+ $X2=0 $Y2=0
cc_723 N_A_1212_471#_c_795_p N_A_1312_126#_c_1611_n 0.00698065f $X=11.62 $Y=3.22
+ $X2=0 $Y2=0
cc_724 N_A_1212_471#_c_769_n N_A_2616_417#_M1039_g 5.35189e-19 $X=12.48 $Y=3.22
+ $X2=0 $Y2=0
cc_725 N_A_1212_471#_c_800_p N_A_2616_417#_c_1693_n 9.74726e-19 $X=12.645
+ $Y=2.39 $X2=0 $Y2=0
cc_726 N_A_1212_471#_c_770_n N_A_2616_417#_c_1693_n 0.076016f $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_727 N_A_1212_471#_c_769_n N_A_2360_115#_M1036_d 0.00743978f $X=12.48 $Y=3.22
+ $X2=0 $Y2=0
cc_728 N_A_1212_471#_c_737_n N_A_2360_115#_c_1785_n 0.0195159f $X=11.55 $Y=1.445
+ $X2=0 $Y2=0
cc_729 N_A_1212_471#_c_737_n N_A_2360_115#_c_1786_n 0.0178577f $X=11.55 $Y=1.445
+ $X2=0 $Y2=0
cc_730 N_A_1212_471#_c_768_n N_A_2360_115#_c_1786_n 0.0304295f $X=11.395 $Y=1.63
+ $X2=0 $Y2=0
cc_731 N_A_1212_471#_c_737_n N_A_2360_115#_c_1795_n 2.90797e-19 $X=11.55
+ $Y=1.445 $X2=0 $Y2=0
cc_732 N_A_1212_471#_c_768_n N_A_2360_115#_c_1795_n 0.00618173f $X=11.395
+ $Y=1.63 $X2=0 $Y2=0
cc_733 N_A_1212_471#_c_798_p N_A_2360_115#_c_1795_n 0.0257423f $X=11.705
+ $Y=3.135 $X2=0 $Y2=0
cc_734 N_A_1212_471#_c_769_n N_A_2360_115#_c_1795_n 0.0243646f $X=12.48 $Y=3.22
+ $X2=0 $Y2=0
cc_735 N_A_1212_471#_c_800_p N_A_2360_115#_c_1795_n 0.0488574f $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_736 N_A_1212_471#_c_770_n N_A_2360_115#_c_1795_n 0.0109388f $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_737 N_A_1212_471#_c_772_n N_A_2360_115#_c_1795_n 0.0112449f $X=11.705 $Y=2.37
+ $X2=0 $Y2=0
cc_738 N_A_1212_471#_c_800_p N_A_2360_115#_c_1796_n 0.0229371f $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_739 N_A_1212_471#_c_770_n N_A_2360_115#_c_1796_n 0.00794057f $X=12.645
+ $Y=2.39 $X2=0 $Y2=0
cc_740 N_A_1212_471#_c_737_n N_A_2360_115#_c_1797_n 0.00391904f $X=11.55
+ $Y=1.445 $X2=0 $Y2=0
cc_741 N_A_1212_471#_c_768_n N_A_2360_115#_c_1797_n 0.0129427f $X=11.395 $Y=1.63
+ $X2=0 $Y2=0
cc_742 N_A_1212_471#_c_772_n N_A_2360_115#_c_1797_n 0.00854125f $X=11.705
+ $Y=2.37 $X2=0 $Y2=0
cc_743 N_A_1212_471#_c_800_p N_A_2360_115#_c_1798_n 0.0345071f $X=12.645 $Y=2.39
+ $X2=0 $Y2=0
cc_744 N_A_1212_471#_c_770_n N_A_2360_115#_c_1798_n 0.00728856f $X=12.645
+ $Y=2.39 $X2=0 $Y2=0
cc_745 N_A_1212_471#_c_769_n N_A_2360_115#_c_1800_n 0.00399632f $X=12.48 $Y=3.22
+ $X2=0 $Y2=0
cc_746 N_A_1212_471#_c_770_n N_A_2360_115#_c_1800_n 8.00152e-19 $X=12.645
+ $Y=2.39 $X2=0 $Y2=0
cc_747 N_A_1212_471#_c_737_n N_A_2360_115#_c_1788_n 0.00783081f $X=11.55
+ $Y=1.445 $X2=0 $Y2=0
cc_748 N_A_1212_471#_c_750_n N_A_65_649#_c_2068_n 0.0026513f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_749 N_A_1212_471#_c_756_n N_A_65_649#_c_2068_n 0.0114843f $X=6.355 $Y=3.72
+ $X2=0 $Y2=0
cc_750 N_A_1212_471#_c_738_n N_A_65_649#_c_2050_n 0.185627f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_751 N_A_1212_471#_c_750_n N_A_65_649#_c_2053_n 0.024249f $X=6.27 $Y=2.54
+ $X2=0 $Y2=0
cc_752 N_A_1212_471#_c_759_n N_VPWR_M1015_d 0.00246135f $X=8.535 $Y=3.15 $X2=0
+ $Y2=0
cc_753 N_A_1212_471#_c_795_p N_VPWR_M1020_d 0.0103009f $X=11.62 $Y=3.22 $X2=0
+ $Y2=0
cc_754 N_A_1212_471#_c_753_n N_VPWR_c_2205_n 0.00432577f $X=7.045 $Y=3.72 $X2=0
+ $Y2=0
cc_755 N_A_1212_471#_c_786_p N_VPWR_c_2205_n 0.0135786f $X=7.13 $Y=3.635 $X2=0
+ $Y2=0
cc_756 N_A_1212_471#_c_759_n N_VPWR_c_2205_n 0.0526181f $X=8.535 $Y=3.15 $X2=0
+ $Y2=0
cc_757 N_A_1212_471#_c_836_p N_VPWR_c_2205_n 0.0102154f $X=8.62 $Y=3.635 $X2=0
+ $Y2=0
cc_758 N_A_1212_471#_c_763_n N_VPWR_c_2205_n 0.00457995f $X=8.705 $Y=3.72 $X2=0
+ $Y2=0
cc_759 N_A_1212_471#_c_760_n N_VPWR_c_2208_n 0.00696789f $X=9.455 $Y=3.72 $X2=0
+ $Y2=0
cc_760 N_A_1212_471#_c_767_n N_VPWR_c_2208_n 0.00946989f $X=9.62 $Y=3.635 $X2=0
+ $Y2=0
cc_761 N_A_1212_471#_c_795_p N_VPWR_c_2208_n 0.0507008f $X=11.62 $Y=3.22 $X2=0
+ $Y2=0
cc_762 N_A_1212_471#_c_738_n N_VPWR_c_2220_n 0.0199629f $X=6.27 $Y=2.54 $X2=0
+ $Y2=0
cc_763 N_A_1212_471#_c_750_n N_VPWR_c_2220_n 0.0179039f $X=6.27 $Y=2.54 $X2=0
+ $Y2=0
cc_764 N_A_1212_471#_c_753_n N_VPWR_c_2220_n 0.0312412f $X=7.045 $Y=3.72 $X2=0
+ $Y2=0
cc_765 N_A_1212_471#_c_756_n N_VPWR_c_2220_n 0.00522478f $X=6.355 $Y=3.72 $X2=0
+ $Y2=0
cc_766 N_A_1212_471#_c_786_p N_VPWR_c_2220_n 0.0137523f $X=7.13 $Y=3.635 $X2=0
+ $Y2=0
cc_767 N_A_1212_471#_c_759_n N_VPWR_c_2220_n 0.0220875f $X=8.535 $Y=3.15 $X2=0
+ $Y2=0
cc_768 N_A_1212_471#_c_836_p N_VPWR_c_2220_n 0.013657f $X=8.62 $Y=3.635 $X2=0
+ $Y2=0
cc_769 N_A_1212_471#_c_760_n N_VPWR_c_2220_n 0.0390924f $X=9.455 $Y=3.72 $X2=0
+ $Y2=0
cc_770 N_A_1212_471#_c_763_n N_VPWR_c_2220_n 0.00732918f $X=8.705 $Y=3.72 $X2=0
+ $Y2=0
cc_771 N_A_1212_471#_c_767_n N_VPWR_c_2220_n 0.0348182f $X=9.62 $Y=3.635 $X2=0
+ $Y2=0
cc_772 N_A_1212_471#_c_795_p N_VPWR_c_2220_n 0.0678272f $X=11.62 $Y=3.22 $X2=0
+ $Y2=0
cc_773 N_A_1212_471#_c_769_n N_VPWR_c_2220_n 0.0540969f $X=12.48 $Y=3.22 $X2=0
+ $Y2=0
cc_774 N_A_1212_471#_c_770_n N_VPWR_c_2220_n 0.00189764f $X=12.645 $Y=2.39 $X2=0
+ $Y2=0
cc_775 N_A_1212_471#_c_802_p N_VPWR_c_2220_n 0.00862856f $X=11.705 $Y=3.22 $X2=0
+ $Y2=0
cc_776 N_A_1212_471#_c_759_n A_1468_641# 9.88449e-19 $X=8.535 $Y=3.15 $X2=0
+ $Y2=0
cc_777 N_A_1212_471#_c_745_n N_VGND_c_2398_n 0.0638635f $X=9.305 $Y=1.26 $X2=0
+ $Y2=0
cc_778 N_A_1212_471#_c_746_n N_VGND_c_2398_n 0.00761835f $X=9.47 $Y=1.115 $X2=0
+ $Y2=0
cc_779 N_A_1212_471#_c_746_n N_VGND_c_2400_n 0.0310984f $X=9.47 $Y=1.115 $X2=0
+ $Y2=0
cc_780 N_A_1212_471#_c_737_n N_VGND_c_2408_n 0.024275f $X=11.55 $Y=1.445 $X2=0
+ $Y2=0
cc_781 N_A_1212_471#_c_738_n N_VGND_c_2408_n 0.0222636f $X=6.27 $Y=2.54 $X2=0
+ $Y2=0
cc_782 N_A_1212_471#_c_739_n N_VGND_c_2408_n 0.037633f $X=7.045 $Y=0.35 $X2=0
+ $Y2=0
cc_783 N_A_1212_471#_c_741_n N_VGND_c_2408_n 0.00925191f $X=6.355 $Y=0.35 $X2=0
+ $Y2=0
cc_784 N_A_1212_471#_c_743_n N_VGND_c_2408_n 0.027332f $X=7.15 $Y=1.175 $X2=0
+ $Y2=0
cc_785 N_A_1212_471#_c_745_n N_VGND_c_2408_n 0.0374186f $X=9.305 $Y=1.26 $X2=0
+ $Y2=0
cc_786 N_A_1212_471#_c_746_n N_VGND_c_2408_n 0.0164336f $X=9.47 $Y=1.115 $X2=0
+ $Y2=0
cc_787 N_A_1212_471#_M1001_g N_VGND_c_2408_n 0.0122633f $X=7.09 $Y=0.84 $X2=0
+ $Y2=0
cc_788 N_A_1212_100#_c_981_n N_A_1510_100#_M1010_g 0.00917694f $X=7.52 $Y=1.915
+ $X2=0 $Y2=0
cc_789 N_A_1212_100#_c_982_n N_A_1510_100#_M1010_g 0.0270427f $X=10.61 $Y=1.61
+ $X2=0 $Y2=0
cc_790 N_A_1212_100#_c_983_n N_A_1510_100#_M1010_g 0.00247675f $X=7.605 $Y=1.61
+ $X2=0 $Y2=0
cc_791 N_A_1212_100#_M1003_g N_A_1510_100#_M1015_g 0.0575237f $X=7.09 $Y=3.415
+ $X2=0 $Y2=0
cc_792 N_A_1212_100#_c_978_n N_A_1510_100#_c_1246_n 0.0479886f $X=10.01 $Y=2.585
+ $X2=18.96 $Y2=0
cc_793 N_A_1212_100#_c_982_n N_A_1510_100#_c_1246_n 0.180867f $X=10.61 $Y=1.61
+ $X2=18.96 $Y2=0
cc_794 N_A_1212_100#_c_1070_n N_A_1510_100#_c_1267_n 0.0614367f $X=10.695
+ $Y=1.525 $X2=9.6 $Y2=0
cc_795 N_A_1212_100#_c_984_n N_A_1510_100#_c_1267_n 0.0223253f $X=12.285 $Y=0.35
+ $X2=9.6 $Y2=0
cc_796 N_A_1212_100#_c_982_n N_A_1510_100#_c_1247_n 0.0123662f $X=10.61 $Y=1.61
+ $X2=0 $Y2=0
cc_797 N_A_1212_100#_c_979_n N_A_1510_100#_c_1253_n 0.00120882f $X=12.085
+ $Y=2.155 $X2=0 $Y2=0
cc_798 N_A_1212_100#_c_1005_n N_A_1510_100#_c_1292_n 0.00127398f $X=7.09
+ $Y=2.635 $X2=0 $Y2=0
cc_799 N_A_1212_100#_c_1062_n N_A_1510_100#_c_1292_n 0.0117f $X=7.115 $Y=2.11
+ $X2=0 $Y2=0
cc_800 N_A_1212_100#_c_981_n N_A_1510_100#_c_1292_n 0.0029097f $X=7.52 $Y=1.915
+ $X2=0 $Y2=0
cc_801 N_A_1212_100#_c_982_n N_A_1510_100#_c_1292_n 0.0241903f $X=10.61 $Y=1.61
+ $X2=0 $Y2=0
cc_802 N_A_1212_100#_c_1023_n N_A_1510_100#_c_1292_n 0.0133233f $X=7.52 $Y=2
+ $X2=0 $Y2=0
cc_803 N_A_1212_100#_c_1005_n N_A_1510_100#_c_1248_n 0.0677606f $X=7.09 $Y=2.635
+ $X2=0 $Y2=0
cc_804 N_A_1212_100#_c_1062_n N_A_1510_100#_c_1248_n 0.00186963f $X=7.115
+ $Y=2.11 $X2=0 $Y2=0
cc_805 N_A_1212_100#_c_981_n N_A_1510_100#_c_1248_n 0.00317498f $X=7.52 $Y=1.915
+ $X2=0 $Y2=0
cc_806 N_A_1212_100#_c_982_n N_A_1510_100#_c_1248_n 0.00228287f $X=10.61 $Y=1.61
+ $X2=0 $Y2=0
cc_807 N_A_1212_100#_c_1023_n N_A_1510_100#_c_1248_n 0.00707302f $X=7.52 $Y=2
+ $X2=0 $Y2=0
cc_808 N_A_1212_100#_M1020_g N_A_1510_100#_c_1256_n 0.00108976f $X=10.01 $Y=3.09
+ $X2=0 $Y2=0
cc_809 N_A_1212_100#_c_1013_n N_A_1510_100#_c_1256_n 0.00588296f $X=11.665
+ $Y=2.605 $X2=0 $Y2=0
cc_810 N_A_1212_100#_M1022_g N_RESET_B_c_1352_n 0.0339467f $X=6.31 $Y=0.84 $X2=0
+ $Y2=0
cc_811 N_A_1212_100#_c_977_n N_RESET_B_c_1357_n 0.00370456f $X=9.86 $Y=1.435
+ $X2=0 $Y2=0
cc_812 N_A_1212_100#_c_978_n N_RESET_B_c_1357_n 0.0523495f $X=10.01 $Y=2.585
+ $X2=0 $Y2=0
cc_813 N_A_1212_100#_c_982_n N_RESET_B_c_1357_n 0.0165681f $X=10.61 $Y=1.61
+ $X2=0 $Y2=0
cc_814 N_A_1212_100#_c_1004_n N_RESET_B_c_1365_n 0.00599363f $X=6.56 $Y=2.03
+ $X2=0 $Y2=0
cc_815 N_A_1212_100#_c_1005_n N_RESET_B_c_1365_n 0.00803019f $X=7.09 $Y=2.635
+ $X2=0 $Y2=0
cc_816 N_A_1212_100#_c_1062_n N_RESET_B_c_1365_n 0.0178259f $X=7.115 $Y=2.11
+ $X2=0 $Y2=0
cc_817 N_A_1212_100#_c_1023_n N_RESET_B_c_1365_n 0.0100035f $X=7.52 $Y=2 $X2=0
+ $Y2=0
cc_818 N_A_1212_100#_c_978_n N_RESET_B_c_1367_n 0.0313364f $X=10.01 $Y=2.585
+ $X2=0 $Y2=0
cc_819 N_A_1212_100#_c_979_n N_RESET_B_c_1367_n 0.0166454f $X=12.085 $Y=2.155
+ $X2=0 $Y2=0
cc_820 N_A_1212_100#_c_990_n N_RESET_B_c_1370_n 0.00156416f $X=14.225 $Y=1.63
+ $X2=0 $Y2=0
cc_821 N_A_1212_100#_c_982_n N_RESET_B_c_1359_n 0.0151242f $X=10.61 $Y=1.61
+ $X2=0 $Y2=0
cc_822 N_A_1212_100#_c_978_n N_RESET_B_c_1375_n 2.64494e-19 $X=10.01 $Y=2.585
+ $X2=0 $Y2=0
cc_823 N_A_1212_100#_c_990_n N_RESET_B_M1025_g 0.0244469f $X=14.225 $Y=1.63
+ $X2=0 $Y2=0
cc_824 N_A_1212_100#_c_991_n N_RESET_B_M1025_g 0.0350248f $X=14.31 $Y=1.545
+ $X2=0 $Y2=0
cc_825 N_A_1212_100#_c_992_n N_RESET_B_M1025_g 0.00576606f $X=15.755 $Y=0.62
+ $X2=0 $Y2=0
cc_826 N_A_1212_100#_c_990_n N_RESET_B_c_1457_n 0.0241181f $X=14.225 $Y=1.63
+ $X2=0 $Y2=0
cc_827 N_A_1212_100#_c_977_n N_A_1312_126#_M1007_g 0.0172069f $X=9.86 $Y=1.435
+ $X2=0 $Y2=0
cc_828 N_A_1212_100#_c_982_n N_A_1312_126#_M1007_g 0.0168869f $X=10.61 $Y=1.61
+ $X2=0 $Y2=0
cc_829 N_A_1212_100#_c_1070_n N_A_1312_126#_M1007_g 0.0447675f $X=10.695
+ $Y=1.525 $X2=0 $Y2=0
cc_830 N_A_1212_100#_c_984_n N_A_1312_126#_M1007_g 0.00861305f $X=12.285 $Y=0.35
+ $X2=0 $Y2=0
cc_831 N_A_1212_100#_c_978_n N_A_1312_126#_c_1562_n 0.0553689f $X=10.01 $Y=2.585
+ $X2=0 $Y2=0
cc_832 N_A_1212_100#_M1020_g N_A_1312_126#_c_1562_n 0.0361537f $X=10.01 $Y=3.09
+ $X2=0 $Y2=0
cc_833 N_A_1212_100#_c_979_n N_A_1312_126#_c_1562_n 0.0601121f $X=12.085
+ $Y=2.155 $X2=0 $Y2=0
cc_834 N_A_1212_100#_M1022_g N_A_1312_126#_c_1563_n 0.0242357f $X=6.31 $Y=0.84
+ $X2=0 $Y2=0
cc_835 N_A_1212_100#_c_1003_n N_A_1312_126#_c_1563_n 0.0120078f $X=6.8 $Y=2.03
+ $X2=0 $Y2=0
cc_836 N_A_1212_100#_c_1004_n N_A_1312_126#_c_1563_n 0.00303105f $X=6.56 $Y=2.03
+ $X2=0 $Y2=0
cc_837 N_A_1212_100#_c_1005_n N_A_1312_126#_c_1563_n 0.0101641f $X=7.09 $Y=2.635
+ $X2=0 $Y2=0
cc_838 N_A_1212_100#_M1003_g N_A_1312_126#_c_1563_n 0.00179481f $X=7.09 $Y=3.415
+ $X2=0 $Y2=0
cc_839 N_A_1212_100#_c_1062_n N_A_1312_126#_c_1563_n 0.0240909f $X=7.115 $Y=2.11
+ $X2=0 $Y2=0
cc_840 N_A_1212_100#_c_1023_n N_A_1312_126#_c_1563_n 0.0097606f $X=7.52 $Y=2
+ $X2=0 $Y2=0
cc_841 N_A_1212_100#_M1003_g N_A_1312_126#_c_1589_n 0.0146041f $X=7.09 $Y=3.415
+ $X2=9.6 $Y2=0
cc_842 N_A_1212_100#_M1003_g N_A_1312_126#_c_1569_n 0.0246725f $X=7.09 $Y=3.415
+ $X2=9.6 $Y2=0.057
cc_843 N_A_1212_100#_c_1062_n N_A_1312_126#_c_1569_n 0.0211693f $X=7.115 $Y=2.11
+ $X2=9.6 $Y2=0.057
cc_844 N_A_1212_100#_c_1023_n N_A_1312_126#_c_1569_n 0.00360334f $X=7.52 $Y=2
+ $X2=9.6 $Y2=0.057
cc_845 N_A_1212_100#_M1020_g N_A_1312_126#_c_1570_n 0.00114747f $X=10.01 $Y=3.09
+ $X2=0 $Y2=0
cc_846 N_A_1212_100#_c_978_n N_A_1312_126#_c_1571_n 0.0049249f $X=10.01 $Y=2.585
+ $X2=0 $Y2=0
cc_847 N_A_1212_100#_M1020_g N_A_1312_126#_c_1571_n 0.00299899f $X=10.01 $Y=3.09
+ $X2=0 $Y2=0
cc_848 N_A_1212_100#_c_978_n N_A_1312_126#_c_1572_n 0.0521579f $X=10.01 $Y=2.585
+ $X2=0 $Y2=0
cc_849 N_A_1212_100#_M1022_g N_A_1312_126#_c_1564_n 0.00703965f $X=6.31 $Y=0.84
+ $X2=0 $Y2=0
cc_850 N_A_1212_100#_c_1003_n N_A_1312_126#_c_1574_n 0.00251763f $X=6.8 $Y=2.03
+ $X2=0 $Y2=0
cc_851 N_A_1212_100#_c_1005_n N_A_1312_126#_c_1574_n 0.00212434f $X=7.09
+ $Y=2.635 $X2=0 $Y2=0
cc_852 N_A_1212_100#_M1003_g N_A_1312_126#_c_1574_n 0.00291322f $X=7.09 $Y=3.415
+ $X2=0 $Y2=0
cc_853 N_A_1212_100#_c_978_n N_A_1312_126#_c_1611_n 0.00155157f $X=10.01
+ $Y=2.585 $X2=0 $Y2=0
cc_854 N_A_1212_100#_c_990_n N_A_2616_417#_c_1693_n 0.00157741f $X=14.225
+ $Y=1.63 $X2=0 $Y2=0
cc_855 N_A_1212_100#_c_990_n N_A_2616_417#_c_1694_n 0.0238596f $X=14.225 $Y=1.63
+ $X2=18.96 $Y2=0
cc_856 N_A_1212_100#_c_990_n N_A_2616_417#_c_1689_n 0.0130055f $X=14.225 $Y=1.63
+ $X2=0 $Y2=0
cc_857 N_A_1212_100#_c_991_n N_A_2616_417#_c_1689_n 0.0136329f $X=14.31 $Y=1.545
+ $X2=0 $Y2=0
cc_858 N_A_1212_100#_c_992_n N_A_2616_417#_c_1707_n 0.0128852f $X=15.755 $Y=0.62
+ $X2=0 $Y2=0
cc_859 N_A_1212_100#_c_991_n N_A_2616_417#_c_1708_n 0.00636915f $X=14.31
+ $Y=1.545 $X2=0 $Y2=0
cc_860 N_A_1212_100#_c_992_n N_A_2616_417#_c_1708_n 0.0046542f $X=15.755 $Y=0.62
+ $X2=0 $Y2=0
cc_861 N_A_1212_100#_c_992_n N_A_2616_417#_c_1690_n 0.0233376f $X=15.755 $Y=0.62
+ $X2=0 $Y2=0
cc_862 N_A_1212_100#_c_996_n N_A_2616_417#_c_1690_n 0.0256874f $X=15.92 $Y=0.765
+ $X2=0 $Y2=0
cc_863 N_A_1212_100#_c_998_n N_A_2616_417#_c_1690_n 0.00663941f $X=16.085
+ $Y=1.34 $X2=0 $Y2=0
cc_864 N_A_1212_100#_M1000_g N_A_2616_417#_M1021_g 0.0136465f $X=12.445 $Y=1.115
+ $X2=0 $Y2=0
cc_865 N_A_1212_100#_c_990_n N_A_2616_417#_M1021_g 0.0307464f $X=14.225 $Y=1.63
+ $X2=0 $Y2=0
cc_866 N_A_1212_100#_c_991_n N_A_2616_417#_M1021_g 0.00109266f $X=14.31 $Y=1.545
+ $X2=0 $Y2=0
cc_867 N_A_1212_100#_c_1000_n N_A_2616_417#_M1021_g 0.027576f $X=12.855 $Y=1.65
+ $X2=0 $Y2=0
cc_868 N_A_1212_100#_c_1001_n N_A_2616_417#_M1021_g 2.86787e-19 $X=13.02 $Y=1.65
+ $X2=0 $Y2=0
cc_869 N_A_1212_100#_c_991_n N_A_2360_115#_M1031_g 0.00255495f $X=14.31 $Y=1.545
+ $X2=0 $Y2=0
cc_870 N_A_1212_100#_c_992_n N_A_2360_115#_M1031_g 0.0166587f $X=15.755 $Y=0.62
+ $X2=0 $Y2=0
cc_871 N_A_1212_100#_c_996_n N_A_2360_115#_M1031_g 0.0039208f $X=15.92 $Y=0.765
+ $X2=0 $Y2=0
cc_872 N_A_1212_100#_c_998_n N_A_2360_115#_M1031_g 0.00188093f $X=16.085 $Y=1.34
+ $X2=0 $Y2=0
cc_873 N_A_1212_100#_c_1021_n N_A_2360_115#_M1029_g 9.96725e-19 $X=17.03 $Y=2.04
+ $X2=18.96 $Y2=0
cc_874 N_A_1212_100#_c_997_n N_A_2360_115#_M1005_g 0.00122828f $X=17.03 $Y=1.34
+ $X2=9.6 $Y2=0
cc_875 N_A_1212_100#_c_999_n N_A_2360_115#_M1005_g 5.20907e-19 $X=17.115
+ $Y=1.955 $X2=9.6 $Y2=0
cc_876 N_A_1212_100#_c_997_n N_A_2360_115#_c_1783_n 0.0144407f $X=17.03 $Y=1.34
+ $X2=9.6 $Y2=0.057
cc_877 N_A_1212_100#_c_1021_n N_A_2360_115#_c_1783_n 0.0258322f $X=17.03 $Y=2.04
+ $X2=9.6 $Y2=0.057
cc_878 N_A_1212_100#_c_1022_n N_A_2360_115#_c_1783_n 0.00567965f $X=16.595
+ $Y=2.04 $X2=9.6 $Y2=0.057
cc_879 N_A_1212_100#_c_999_n N_A_2360_115#_c_1783_n 0.0308239f $X=17.115
+ $Y=1.955 $X2=9.6 $Y2=0.057
cc_880 N_A_1212_100#_M1000_g N_A_2360_115#_c_1785_n 0.00609395f $X=12.445
+ $Y=1.115 $X2=0 $Y2=0
cc_881 N_A_1212_100#_c_984_n N_A_2360_115#_c_1785_n 0.0284636f $X=12.285 $Y=0.35
+ $X2=0 $Y2=0
cc_882 N_A_1212_100#_c_989_n N_A_2360_115#_c_1785_n 0.0554217f $X=12.37 $Y=1.545
+ $X2=0 $Y2=0
cc_883 N_A_1212_100#_M1000_g N_A_2360_115#_c_1786_n 6.96423e-19 $X=12.445
+ $Y=1.115 $X2=0 $Y2=0
cc_884 N_A_1212_100#_c_988_n N_A_2360_115#_c_1786_n 0.0159151f $X=12.285 $Y=1.65
+ $X2=0 $Y2=0
cc_885 N_A_1212_100#_c_989_n N_A_2360_115#_c_1786_n 0.00613112f $X=12.37
+ $Y=1.545 $X2=0 $Y2=0
cc_886 N_A_1212_100#_c_1000_n N_A_2360_115#_c_1786_n 0.00506841f $X=12.855
+ $Y=1.65 $X2=0 $Y2=0
cc_887 N_A_1212_100#_c_1013_n N_A_2360_115#_c_1795_n 0.00329083f $X=11.665
+ $Y=2.605 $X2=0 $Y2=0
cc_888 N_A_1212_100#_c_979_n N_A_2360_115#_c_1795_n 0.0225238f $X=12.085
+ $Y=2.155 $X2=0 $Y2=0
cc_889 N_A_1212_100#_c_990_n N_A_2360_115#_c_1796_n 0.0125419f $X=14.225 $Y=1.63
+ $X2=0 $Y2=0
cc_890 N_A_1212_100#_c_1001_n N_A_2360_115#_c_1796_n 0.0337608f $X=13.02 $Y=1.65
+ $X2=0 $Y2=0
cc_891 N_A_1212_100#_c_979_n N_A_2360_115#_c_1797_n 0.0185069f $X=12.085
+ $Y=2.155 $X2=0 $Y2=0
cc_892 N_A_1212_100#_c_988_n N_A_2360_115#_c_1797_n 0.0337608f $X=12.285 $Y=1.65
+ $X2=0 $Y2=0
cc_893 N_A_1212_100#_c_1000_n N_A_2360_115#_c_1797_n 0.0135537f $X=12.855
+ $Y=1.65 $X2=0 $Y2=0
cc_894 N_A_1212_100#_c_997_n N_A_2360_115#_c_1787_n 0.0524061f $X=17.03 $Y=1.34
+ $X2=0 $Y2=0
cc_895 N_A_1212_100#_c_998_n N_A_2360_115#_c_1787_n 0.0242977f $X=16.085 $Y=1.34
+ $X2=0 $Y2=0
cc_896 N_A_1212_100#_c_1021_n N_A_2360_115#_c_1787_n 0.0164773f $X=17.03 $Y=2.04
+ $X2=0 $Y2=0
cc_897 N_A_1212_100#_c_1022_n N_A_2360_115#_c_1787_n 0.0194818f $X=16.595
+ $Y=2.04 $X2=0 $Y2=0
cc_898 N_A_1212_100#_c_999_n N_A_2360_115#_c_1787_n 0.0122207f $X=17.115
+ $Y=1.955 $X2=0 $Y2=0
cc_899 N_A_1212_100#_c_988_n N_A_2360_115#_c_1788_n 0.00736567f $X=12.285
+ $Y=1.65 $X2=0 $Y2=0
cc_900 N_A_1212_100#_c_1000_n N_A_2360_115#_c_1788_n 0.00283623f $X=12.855
+ $Y=1.65 $X2=0 $Y2=0
cc_901 N_A_1212_100#_c_992_n N_CLK_c_1958_n 0.00346924f $X=15.755 $Y=0.62 $X2=0
+ $Y2=0
cc_902 N_A_1212_100#_c_996_n N_CLK_c_1958_n 0.0314829f $X=15.92 $Y=0.765 $X2=0
+ $Y2=0
cc_903 N_A_1212_100#_c_997_n N_CLK_c_1958_n 0.0179735f $X=17.03 $Y=1.34 $X2=0
+ $Y2=0
cc_904 N_A_1212_100#_c_998_n N_CLK_c_1958_n 3.68883e-19 $X=16.085 $Y=1.34 $X2=0
+ $Y2=0
cc_905 N_A_1212_100#_c_997_n N_CLK_c_1960_n 0.00984354f $X=17.03 $Y=1.34 $X2=0
+ $Y2=0
cc_906 N_A_1212_100#_c_998_n N_CLK_c_1960_n 0.0102612f $X=16.085 $Y=1.34 $X2=0
+ $Y2=0
cc_907 N_A_1212_100#_c_1018_n N_CLK_c_1960_n 0.0238722f $X=16.43 $Y=2.84 $X2=0
+ $Y2=0
cc_908 N_A_1212_100#_c_1022_n N_CLK_c_1960_n 0.00236515f $X=16.595 $Y=2.04 $X2=0
+ $Y2=0
cc_909 N_A_1212_100#_c_1018_n N_CLK_c_1964_n 0.0262078f $X=16.43 $Y=2.84 $X2=0
+ $Y2=0
cc_910 N_A_1212_100#_c_1022_n N_CLK_c_1964_n 0.013038f $X=16.595 $Y=2.04 $X2=0
+ $Y2=0
cc_911 N_A_1212_100#_c_997_n N_A_3417_443#_M1005_s 0.00124783f $X=17.03 $Y=1.34
+ $X2=0 $Y2=0
cc_912 N_A_1212_100#_c_997_n N_A_3417_443#_c_1997_n 0.00766824f $X=17.03 $Y=1.34
+ $X2=0 $Y2=0
cc_913 N_A_1212_100#_c_997_n N_A_3417_443#_c_1998_n 0.0126061f $X=17.03 $Y=1.34
+ $X2=0 $Y2=0
cc_914 N_A_1212_100#_c_999_n N_A_3417_443#_c_1998_n 0.00426653f $X=17.115
+ $Y=1.955 $X2=0 $Y2=0
cc_915 N_A_1212_100#_c_1018_n N_A_3417_443#_c_2005_n 0.0291309f $X=16.43 $Y=2.84
+ $X2=0 $Y2=0
cc_916 N_A_1212_100#_c_1021_n N_A_3417_443#_c_2005_n 0.0118721f $X=17.03 $Y=2.04
+ $X2=0 $Y2=0
cc_917 N_A_1212_100#_c_1021_n N_A_3417_443#_c_2012_n 0.0125158f $X=17.03 $Y=2.04
+ $X2=0 $Y2=0
cc_918 N_A_1212_100#_c_999_n N_A_3417_443#_c_2012_n 0.00899938f $X=17.115
+ $Y=1.955 $X2=0 $Y2=0
cc_919 N_A_1212_100#_c_999_n N_A_3417_443#_c_2014_n 0.024172f $X=17.115 $Y=1.955
+ $X2=0 $Y2=0
cc_920 N_A_1212_100#_M1022_g N_A_65_649#_c_2050_n 0.0167967f $X=6.31 $Y=0.84
+ $X2=0 $Y2=0
cc_921 N_A_1212_100#_c_1004_n N_A_65_649#_c_2053_n 0.0167967f $X=6.56 $Y=2.03
+ $X2=0 $Y2=0
cc_922 N_A_1212_100#_M1003_g N_VPWR_c_2205_n 0.0018477f $X=7.09 $Y=3.415 $X2=0
+ $Y2=0
cc_923 N_A_1212_100#_M1020_g N_VPWR_c_2208_n 0.0129328f $X=10.01 $Y=3.09 $X2=0
+ $Y2=0
cc_924 N_A_1212_100#_c_1013_n N_VPWR_c_2208_n 0.00174346f $X=11.665 $Y=2.605
+ $X2=0 $Y2=0
cc_925 N_A_1212_100#_c_1018_n N_VPWR_c_2214_n 0.0358477f $X=16.43 $Y=2.84 $X2=0
+ $Y2=0
cc_926 N_A_1212_100#_M1018_d N_VPWR_c_2220_n 0.00221032f $X=16.29 $Y=2.715 $X2=0
+ $Y2=0
cc_927 N_A_1212_100#_M1003_g N_VPWR_c_2220_n 0.00732976f $X=7.09 $Y=3.415 $X2=0
+ $Y2=0
cc_928 N_A_1212_100#_M1020_g N_VPWR_c_2220_n 0.00693371f $X=10.01 $Y=3.09 $X2=0
+ $Y2=0
cc_929 N_A_1212_100#_c_1013_n N_VPWR_c_2220_n 0.0227189f $X=11.665 $Y=2.605
+ $X2=0 $Y2=0
cc_930 N_A_1212_100#_c_1018_n N_VPWR_c_2220_n 0.023158f $X=16.43 $Y=2.84 $X2=0
+ $Y2=0
cc_931 N_A_1212_100#_c_977_n N_VGND_c_2398_n 0.00375778f $X=9.86 $Y=1.435 $X2=0
+ $Y2=0
cc_932 N_A_1212_100#_c_977_n N_VGND_c_2400_n 0.0442036f $X=9.86 $Y=1.435 $X2=0
+ $Y2=0
cc_933 N_A_1212_100#_c_982_n N_VGND_c_2400_n 0.0454403f $X=10.61 $Y=1.61 $X2=0
+ $Y2=0
cc_934 N_A_1212_100#_c_1070_n N_VGND_c_2400_n 0.0658068f $X=10.695 $Y=1.525
+ $X2=0 $Y2=0
cc_935 N_A_1212_100#_c_986_n N_VGND_c_2400_n 0.00488837f $X=10.78 $Y=0.35 $X2=0
+ $Y2=0
cc_936 N_A_1212_100#_M1000_g N_VGND_c_2402_n 0.00683356f $X=12.445 $Y=1.115
+ $X2=0 $Y2=0
cc_937 N_A_1212_100#_c_984_n N_VGND_c_2402_n 0.00116639f $X=12.285 $Y=0.35 $X2=0
+ $Y2=0
cc_938 N_A_1212_100#_c_989_n N_VGND_c_2402_n 0.0250512f $X=12.37 $Y=1.545 $X2=0
+ $Y2=0
cc_939 N_A_1212_100#_c_990_n N_VGND_c_2402_n 0.0725893f $X=14.225 $Y=1.63 $X2=0
+ $Y2=0
cc_940 N_A_1212_100#_c_991_n N_VGND_c_2402_n 0.0463275f $X=14.31 $Y=1.545 $X2=0
+ $Y2=0
cc_941 N_A_1212_100#_c_994_n N_VGND_c_2402_n 0.0128696f $X=14.395 $Y=0.62 $X2=0
+ $Y2=0
cc_942 N_A_1212_100#_c_992_n N_VGND_c_2404_n 0.0113439f $X=15.755 $Y=0.62 $X2=0
+ $Y2=0
cc_943 N_A_1212_100#_c_996_n N_VGND_c_2404_n 0.020798f $X=15.92 $Y=0.765 $X2=0
+ $Y2=0
cc_944 N_A_1212_100#_c_997_n N_VGND_c_2404_n 0.0342373f $X=17.03 $Y=1.34 $X2=0
+ $Y2=0
cc_945 N_A_1212_100#_M1022_g N_VGND_c_2408_n 0.0182708f $X=6.31 $Y=0.84 $X2=0
+ $Y2=0
cc_946 N_A_1212_100#_c_977_n N_VGND_c_2408_n 0.00736889f $X=9.86 $Y=1.435 $X2=0
+ $Y2=0
cc_947 N_A_1212_100#_M1000_g N_VGND_c_2408_n 0.0105908f $X=12.445 $Y=1.115 $X2=0
+ $Y2=0
cc_948 N_A_1212_100#_c_1070_n N_VGND_c_2408_n 0.0200372f $X=10.695 $Y=1.525
+ $X2=0 $Y2=0
cc_949 N_A_1212_100#_c_984_n N_VGND_c_2408_n 0.0676967f $X=12.285 $Y=0.35 $X2=0
+ $Y2=0
cc_950 N_A_1212_100#_c_986_n N_VGND_c_2408_n 0.00777234f $X=10.78 $Y=0.35 $X2=0
+ $Y2=0
cc_951 N_A_1212_100#_c_989_n N_VGND_c_2408_n 0.0192112f $X=12.37 $Y=1.545 $X2=0
+ $Y2=0
cc_952 N_A_1212_100#_c_992_n N_VGND_c_2408_n 0.0895572f $X=15.755 $Y=0.62 $X2=0
+ $Y2=0
cc_953 N_A_1212_100#_c_994_n N_VGND_c_2408_n 0.0103782f $X=14.395 $Y=0.62 $X2=0
+ $Y2=0
cc_954 N_A_1510_100#_M1010_g N_RESET_B_c_1352_n 0.0354633f $X=7.8 $Y=0.84 $X2=0
+ $Y2=0
cc_955 N_A_1510_100#_M1010_g N_RESET_B_M1013_g 0.0760414f $X=7.8 $Y=0.84 $X2=0
+ $Y2=0
cc_956 N_A_1510_100#_c_1246_n N_RESET_B_c_1357_n 7.86069e-19 $X=10.96 $Y=1.96
+ $X2=0 $Y2=0
cc_957 N_A_1510_100#_c_1246_n N_RESET_B_c_1365_n 0.0037303f $X=10.96 $Y=1.96
+ $X2=0 $Y2=0
cc_958 N_A_1510_100#_c_1292_n N_RESET_B_c_1365_n 0.02923f $X=7.95 $Y=2.035 $X2=0
+ $Y2=0
cc_959 N_A_1510_100#_c_1248_n N_RESET_B_c_1365_n 0.0130501f $X=7.95 $Y=2.035
+ $X2=0 $Y2=0
cc_960 N_A_1510_100#_c_1246_n N_RESET_B_c_1367_n 0.0239427f $X=10.96 $Y=1.96
+ $X2=0 $Y2=0
cc_961 N_A_1510_100#_c_1253_n N_RESET_B_c_1367_n 0.0152129f $X=11.045 $Y=2.675
+ $X2=0 $Y2=0
cc_962 N_A_1510_100#_c_1256_n N_RESET_B_c_1367_n 0.0123023f $X=11.275 $Y=2.855
+ $X2=0 $Y2=0
cc_963 N_A_1510_100#_c_1246_n N_RESET_B_c_1368_n 0.00278225f $X=10.96 $Y=1.96
+ $X2=0 $Y2=0
cc_964 N_A_1510_100#_c_1292_n N_RESET_B_c_1368_n 0.00266896f $X=7.95 $Y=2.035
+ $X2=0 $Y2=0
cc_965 N_A_1510_100#_c_1248_n N_RESET_B_c_1368_n 0.00152404f $X=7.95 $Y=2.035
+ $X2=0 $Y2=0
cc_966 N_A_1510_100#_M1010_g N_RESET_B_c_1359_n 0.0110927f $X=7.8 $Y=0.84 $X2=0
+ $Y2=0
cc_967 N_A_1510_100#_M1015_g N_RESET_B_c_1359_n 0.0418765f $X=7.8 $Y=3.415 $X2=0
+ $Y2=0
cc_968 N_A_1510_100#_c_1246_n N_RESET_B_c_1359_n 0.0279257f $X=10.96 $Y=1.96
+ $X2=0 $Y2=0
cc_969 N_A_1510_100#_c_1292_n N_RESET_B_c_1359_n 0.00161527f $X=7.95 $Y=2.035
+ $X2=0 $Y2=0
cc_970 N_A_1510_100#_c_1248_n N_RESET_B_c_1359_n 0.0359015f $X=7.95 $Y=2.035
+ $X2=0 $Y2=0
cc_971 N_A_1510_100#_c_1246_n N_RESET_B_c_1375_n 0.0298699f $X=10.96 $Y=1.96
+ $X2=0 $Y2=0
cc_972 N_A_1510_100#_c_1292_n N_RESET_B_c_1375_n 0.0209121f $X=7.95 $Y=2.035
+ $X2=0 $Y2=0
cc_973 N_A_1510_100#_c_1248_n N_RESET_B_c_1375_n 0.00193279f $X=7.95 $Y=2.035
+ $X2=0 $Y2=0
cc_974 N_A_1510_100#_c_1267_n N_A_1312_126#_M1007_g 0.0113724f $X=11.16 $Y=0.7
+ $X2=0 $Y2=0
cc_975 N_A_1510_100#_c_1247_n N_A_1312_126#_M1007_g 0.0103674f $X=11.045
+ $Y=1.875 $X2=0 $Y2=0
cc_976 N_A_1510_100#_c_1274_n N_A_1312_126#_M1007_g 0.00364657f $X=11.142
+ $Y=1.285 $X2=0 $Y2=0
cc_977 N_A_1510_100#_c_1246_n N_A_1312_126#_c_1562_n 0.029346f $X=10.96 $Y=1.96
+ $X2=0 $Y2=0
cc_978 N_A_1510_100#_c_1247_n N_A_1312_126#_c_1562_n 0.00869612f $X=11.045
+ $Y=1.875 $X2=0 $Y2=0
cc_979 N_A_1510_100#_c_1253_n N_A_1312_126#_c_1562_n 0.0322884f $X=11.045
+ $Y=2.675 $X2=0 $Y2=0
cc_980 N_A_1510_100#_c_1255_n N_A_1312_126#_c_1562_n 0.00232734f $X=11.045
+ $Y=1.96 $X2=0 $Y2=0
cc_981 N_A_1510_100#_c_1256_n N_A_1312_126#_c_1562_n 0.0143833f $X=11.275
+ $Y=2.855 $X2=0 $Y2=0
cc_982 N_A_1510_100#_M1015_g N_A_1312_126#_c_1589_n 6.33174e-19 $X=7.8 $Y=3.415
+ $X2=9.6 $Y2=0
cc_983 N_A_1510_100#_M1015_g N_A_1312_126#_c_1569_n 0.0269315f $X=7.8 $Y=3.415
+ $X2=9.6 $Y2=0.057
cc_984 N_A_1510_100#_c_1246_n N_A_1312_126#_c_1569_n 0.00296611f $X=10.96
+ $Y=1.96 $X2=9.6 $Y2=0.057
cc_985 N_A_1510_100#_c_1292_n N_A_1312_126#_c_1569_n 0.0221115f $X=7.95 $Y=2.035
+ $X2=9.6 $Y2=0.057
cc_986 N_A_1510_100#_c_1248_n N_A_1312_126#_c_1569_n 0.00239678f $X=7.95
+ $Y=2.035 $X2=9.6 $Y2=0.057
cc_987 N_A_1510_100#_c_1246_n N_A_1312_126#_c_1572_n 0.0781323f $X=10.96 $Y=1.96
+ $X2=0 $Y2=0
cc_988 N_A_1510_100#_c_1246_n N_A_1312_126#_c_1573_n 0.0128271f $X=10.96 $Y=1.96
+ $X2=0 $Y2=0
cc_989 N_A_1510_100#_c_1246_n N_A_1312_126#_c_1575_n 0.00189909f $X=10.96
+ $Y=1.96 $X2=0 $Y2=0
cc_990 N_A_1510_100#_c_1246_n N_A_1312_126#_c_1611_n 0.0183772f $X=10.96 $Y=1.96
+ $X2=0 $Y2=0
cc_991 N_A_1510_100#_c_1253_n N_A_1312_126#_c_1611_n 0.0213714f $X=11.045
+ $Y=2.675 $X2=0 $Y2=0
cc_992 N_A_1510_100#_c_1267_n N_A_2360_115#_c_1785_n 0.014954f $X=11.16 $Y=0.7
+ $X2=0 $Y2=0
cc_993 N_A_1510_100#_c_1247_n N_A_2360_115#_c_1788_n 0.00552992f $X=11.045
+ $Y=1.875 $X2=0 $Y2=0
cc_994 N_A_1510_100#_c_1274_n N_A_2360_115#_c_1788_n 0.014954f $X=11.142
+ $Y=1.285 $X2=0 $Y2=0
cc_995 N_A_1510_100#_M1015_g N_VPWR_c_2205_n 0.0253653f $X=7.8 $Y=3.415 $X2=0
+ $Y2=0
cc_996 N_A_1510_100#_M1009_d N_VPWR_c_2220_n 0.00235311f $X=11.135 $Y=2.715
+ $X2=0 $Y2=0
cc_997 N_A_1510_100#_M1015_g N_VPWR_c_2220_n 0.00514822f $X=7.8 $Y=3.415 $X2=0
+ $Y2=0
cc_998 N_A_1510_100#_M1010_g N_VGND_c_2398_n 0.0144251f $X=7.8 $Y=0.84 $X2=0
+ $Y2=0
cc_999 N_A_1510_100#_M1010_g N_VGND_c_2408_n 0.0140299f $X=7.8 $Y=0.84 $X2=0
+ $Y2=0
cc_1000 N_A_1510_100#_c_1267_n N_VGND_c_2408_n 0.0252188f $X=11.16 $Y=0.7 $X2=0
+ $Y2=0
cc_1001 N_RESET_B_c_1367_n N_A_1312_126#_c_1562_n 0.0113988f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1002 N_RESET_B_c_1365_n N_A_1312_126#_c_1563_n 0.0193149f $X=8.255 $Y=2.405
+ $X2=0 $Y2=0
cc_1003 N_RESET_B_c_1365_n N_A_1312_126#_c_1569_n 0.0262255f $X=8.255 $Y=2.405
+ $X2=9.6 $Y2=0.057
cc_1004 N_RESET_B_c_1367_n N_A_1312_126#_c_1569_n 0.00432755f $X=14.015 $Y=2.405
+ $X2=9.6 $Y2=0.057
cc_1005 N_RESET_B_c_1368_n N_A_1312_126#_c_1569_n 0.00307561f $X=8.545 $Y=2.405
+ $X2=9.6 $Y2=0.057
cc_1006 N_RESET_B_c_1359_n N_A_1312_126#_c_1569_n 0.026216f $X=8.595 $Y=2.38
+ $X2=9.6 $Y2=0.057
cc_1007 N_RESET_B_c_1375_n N_A_1312_126#_c_1569_n 0.0295423f $X=8.595 $Y=2.38
+ $X2=9.6 $Y2=0.057
cc_1008 N_RESET_B_c_1359_n N_A_1312_126#_c_1570_n 0.02144f $X=8.595 $Y=2.38
+ $X2=0 $Y2=0
cc_1009 N_RESET_B_c_1367_n N_A_1312_126#_c_1571_n 0.0143502f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1010 N_RESET_B_c_1368_n N_A_1312_126#_c_1571_n 2.15736e-19 $X=8.545 $Y=2.405
+ $X2=0 $Y2=0
cc_1011 N_RESET_B_c_1359_n N_A_1312_126#_c_1571_n 0.00759078f $X=8.595 $Y=2.38
+ $X2=0 $Y2=0
cc_1012 N_RESET_B_c_1375_n N_A_1312_126#_c_1571_n 0.00600223f $X=8.595 $Y=2.38
+ $X2=0 $Y2=0
cc_1013 N_RESET_B_c_1367_n N_A_1312_126#_c_1572_n 0.0426866f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1014 N_RESET_B_c_1367_n N_A_1312_126#_c_1573_n 0.00421488f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1015 N_RESET_B_c_1368_n N_A_1312_126#_c_1573_n 2.52703e-19 $X=8.545 $Y=2.405
+ $X2=0 $Y2=0
cc_1016 N_RESET_B_c_1359_n N_A_1312_126#_c_1573_n 0.00162219f $X=8.595 $Y=2.38
+ $X2=0 $Y2=0
cc_1017 N_RESET_B_c_1375_n N_A_1312_126#_c_1573_n 0.00855983f $X=8.595 $Y=2.38
+ $X2=0 $Y2=0
cc_1018 N_RESET_B_c_1352_n N_A_1312_126#_c_1564_n 0.00135567f $X=8.26 $Y=0.215
+ $X2=0 $Y2=0
cc_1019 N_RESET_B_c_1365_n N_A_1312_126#_c_1574_n 0.00752338f $X=8.255 $Y=2.405
+ $X2=0 $Y2=0
cc_1020 N_RESET_B_c_1367_n N_A_1312_126#_c_1575_n 0.00496778f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1021 N_RESET_B_c_1359_n N_A_1312_126#_c_1575_n 0.00452678f $X=8.595 $Y=2.38
+ $X2=0 $Y2=0
cc_1022 N_RESET_B_c_1367_n N_A_1312_126#_c_1611_n 0.0241999f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1023 N_RESET_B_M1025_g N_A_2616_417#_M1039_g 0.0201678f $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1024 N_RESET_B_c_1367_n N_A_2616_417#_c_1693_n 0.0118025f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1025 N_RESET_B_c_1370_n N_A_2616_417#_c_1693_n 0.00136636f $X=14.16 $Y=2.405
+ $X2=0 $Y2=0
cc_1026 N_RESET_B_c_1367_n N_A_2616_417#_c_1694_n 0.0307358f $X=14.015 $Y=2.405
+ $X2=18.96 $Y2=0
cc_1027 N_RESET_B_c_1370_n N_A_2616_417#_c_1694_n 0.00283687f $X=14.16 $Y=2.405
+ $X2=18.96 $Y2=0
cc_1028 N_RESET_B_M1025_g N_A_2616_417#_c_1694_n 0.00483742f $X=14.27 $Y=1.115
+ $X2=18.96 $Y2=0
cc_1029 N_RESET_B_c_1457_n N_A_2616_417#_c_1694_n 0.0233474f $X=14.205 $Y=2.025
+ $X2=18.96 $Y2=0
cc_1030 N_RESET_B_c_1367_n N_A_2616_417#_c_1695_n 0.01339f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1031 N_RESET_B_c_1370_n N_A_2616_417#_c_1695_n 0.00741821f $X=14.16 $Y=2.405
+ $X2=0 $Y2=0
cc_1032 N_RESET_B_M1025_g N_A_2616_417#_c_1695_n 0.0286158f $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1033 N_RESET_B_c_1457_n N_A_2616_417#_c_1695_n 0.0195319f $X=14.205 $Y=2.025
+ $X2=0 $Y2=0
cc_1034 N_RESET_B_M1025_g N_A_2616_417#_c_1696_n 0.0113809f $X=14.27 $Y=1.115
+ $X2=9.6 $Y2=0.057
cc_1035 N_RESET_B_c_1370_n N_A_2616_417#_c_1689_n 0.00244354f $X=14.16 $Y=2.405
+ $X2=0 $Y2=0
cc_1036 N_RESET_B_M1025_g N_A_2616_417#_c_1689_n 0.0162376f $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1037 N_RESET_B_c_1457_n N_A_2616_417#_c_1689_n 0.0374859f $X=14.205 $Y=2.025
+ $X2=0 $Y2=0
cc_1038 N_RESET_B_M1025_g N_A_2616_417#_c_1708_n 8.04259e-19 $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1039 N_RESET_B_M1025_g N_A_2616_417#_c_1698_n 0.00213848f $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1040 N_RESET_B_M1025_g N_A_2616_417#_c_1690_n 8.88372e-19 $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1041 N_RESET_B_M1025_g N_A_2616_417#_M1021_g 0.0690079f $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1042 N_RESET_B_c_1457_n N_A_2616_417#_M1021_g 0.00253227f $X=14.205 $Y=2.025
+ $X2=0 $Y2=0
cc_1043 N_RESET_B_M1025_g N_A_2360_115#_M1031_g 0.100208f $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1044 N_RESET_B_M1025_g N_A_2360_115#_M1028_g 0.0251803f $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1045 N_RESET_B_c_1367_n N_A_2360_115#_c_1795_n 0.0281036f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1046 N_RESET_B_c_1367_n N_A_2360_115#_c_1796_n 0.011426f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1047 N_RESET_B_c_1367_n N_A_2360_115#_c_1797_n 0.0170464f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1048 N_RESET_B_c_1367_n N_A_2360_115#_c_1798_n 0.0227883f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1049 N_RESET_B_c_1367_n N_A_2360_115#_c_1799_n 0.00616205f $X=14.015 $Y=2.405
+ $X2=0 $Y2=0
cc_1050 N_RESET_B_M1025_g N_A_2360_115#_c_1799_n 0.0159669f $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1051 N_RESET_B_M1025_g N_A_2360_115#_c_1801_n 0.00707973f $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1052 N_RESET_B_M1025_g N_A_2360_115#_c_1802_n 0.00669605f $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1053 N_RESET_B_M1025_g N_A_2360_115#_c_1808_n 5.40048e-19 $X=14.27 $Y=1.115
+ $X2=0 $Y2=0
cc_1054 N_RESET_B_c_1457_n N_A_2360_115#_c_1789_n 3.05158e-19 $X=14.205 $Y=2.025
+ $X2=0 $Y2=0
cc_1055 N_RESET_B_M1019_g N_A_65_649#_c_2059_n 5.57277e-19 $X=3.86 $Y=3.455
+ $X2=0 $Y2=0
cc_1056 N_RESET_B_M1019_g N_A_65_649#_c_2065_n 6.5786e-19 $X=3.86 $Y=3.455 $X2=0
+ $Y2=0
cc_1057 N_RESET_B_M1019_g N_A_65_649#_c_2066_n 0.0152175f $X=3.86 $Y=3.455 $X2=0
+ $Y2=0
cc_1058 N_RESET_B_c_1364_n N_A_65_649#_c_2066_n 0.0187892f $X=3.965 $Y=3.115
+ $X2=0 $Y2=0
cc_1059 N_RESET_B_M1019_g N_A_65_649#_c_2099_n 6.20364e-19 $X=3.86 $Y=3.455
+ $X2=0 $Y2=0
cc_1060 N_RESET_B_M1019_g N_A_65_649#_c_2071_n 5.55461e-19 $X=3.86 $Y=3.455
+ $X2=0 $Y2=0
cc_1061 N_RESET_B_c_1352_n N_A_65_649#_c_2050_n 0.00403218f $X=8.26 $Y=0.215
+ $X2=0 $Y2=0
cc_1062 N_RESET_B_c_1365_n N_A_65_649#_c_2053_n 0.0236862f $X=8.255 $Y=2.405
+ $X2=0 $Y2=0
cc_1063 N_RESET_B_M1019_g N_VPWR_c_2202_n 0.020198f $X=3.86 $Y=3.455 $X2=0 $Y2=0
cc_1064 N_RESET_B_c_1364_n N_VPWR_c_2202_n 0.00103515f $X=3.965 $Y=3.115 $X2=0
+ $Y2=0
cc_1065 N_RESET_B_c_1359_n N_VPWR_c_2205_n 0.00205448f $X=8.595 $Y=2.38 $X2=0
+ $Y2=0
cc_1066 N_RESET_B_M1019_g N_VPWR_c_2220_n 0.0072521f $X=3.86 $Y=3.455 $X2=0
+ $Y2=0
cc_1067 N_RESET_B_c_1359_n N_VPWR_c_2220_n 0.00912067f $X=8.595 $Y=2.38 $X2=0
+ $Y2=0
cc_1068 N_RESET_B_M1025_g N_VPWR_c_2220_n 0.00395199f $X=14.27 $Y=1.115 $X2=0
+ $Y2=0
cc_1069 N_RESET_B_M1024_g N_noxref_23_c_2365_n 0.00616693f $X=4.2 $Y=0.84
+ $X2=0.24 $Y2=0
cc_1070 N_RESET_B_c_1353_n N_noxref_23_c_2365_n 0.00140362f $X=4.45 $Y=0.215
+ $X2=0.24 $Y2=0
cc_1071 N_RESET_B_M1024_g N_noxref_23_c_2369_n 0.0114708f $X=4.2 $Y=0.84 $X2=0
+ $Y2=0
cc_1072 N_RESET_B_M1024_g N_VGND_c_2396_n 0.0367801f $X=4.2 $Y=0.84 $X2=0 $Y2=0
cc_1073 N_RESET_B_c_1352_n N_VGND_c_2396_n 0.00634114f $X=8.26 $Y=0.215 $X2=0
+ $Y2=0
cc_1074 N_RESET_B_c_1352_n N_VGND_c_2398_n 0.00108269f $X=8.26 $Y=0.215 $X2=0
+ $Y2=0
cc_1075 N_RESET_B_M1013_g N_VGND_c_2398_n 0.0528841f $X=8.51 $Y=0.84 $X2=0 $Y2=0
cc_1076 N_RESET_B_c_1357_n N_VGND_c_2398_n 0.00410388f $X=8.585 $Y=1.585 $X2=0
+ $Y2=0
cc_1077 N_RESET_B_M1025_g N_VGND_c_2402_n 0.0125737f $X=14.27 $Y=1.115 $X2=0
+ $Y2=0
cc_1078 N_RESET_B_M1024_g N_VGND_c_2408_n 0.00401816f $X=4.2 $Y=0.84 $X2=0 $Y2=0
cc_1079 N_RESET_B_c_1352_n N_VGND_c_2408_n 0.0392709f $X=8.26 $Y=0.215 $X2=0
+ $Y2=0
cc_1080 N_RESET_B_c_1353_n N_VGND_c_2408_n 0.00177478f $X=4.45 $Y=0.215 $X2=0
+ $Y2=0
cc_1081 N_RESET_B_M1013_g N_VGND_c_2408_n 0.00245024f $X=8.51 $Y=0.84 $X2=0
+ $Y2=0
cc_1082 N_RESET_B_M1025_g N_VGND_c_2408_n 0.00612806f $X=14.27 $Y=1.115 $X2=0
+ $Y2=0
cc_1083 N_A_1312_126#_M1007_g N_A_2360_115#_c_1785_n 4.26829e-19 $X=10.77
+ $Y=0.95 $X2=0 $Y2=0
cc_1084 N_A_1312_126#_c_1562_n N_VPWR_c_2208_n 0.0158699f $X=10.885 $Y=2.605
+ $X2=0 $Y2=0
cc_1085 N_A_1312_126#_c_1562_n N_VPWR_c_2220_n 0.0116266f $X=10.885 $Y=2.605
+ $X2=0 $Y2=0
cc_1086 N_A_1312_126#_c_1589_n N_VPWR_c_2220_n 0.0227597f $X=6.7 $Y=3.35 $X2=0
+ $Y2=0
cc_1087 N_A_1312_126#_c_1569_n N_VPWR_c_2220_n 0.0114897f $X=8.885 $Y=2.8 $X2=0
+ $Y2=0
cc_1088 N_A_1312_126#_c_1570_n N_VPWR_c_2220_n 0.0228033f $X=9.05 $Y=3.35 $X2=0
+ $Y2=0
cc_1089 N_A_1312_126#_M1007_g N_VGND_c_2400_n 0.00606092f $X=10.77 $Y=0.95 $X2=0
+ $Y2=0
cc_1090 N_A_1312_126#_M1007_g N_VGND_c_2408_n 0.0189078f $X=10.77 $Y=0.95 $X2=0
+ $Y2=0
cc_1091 N_A_1312_126#_c_1563_n N_VGND_c_2408_n 4.53408e-19 $X=6.62 $Y=2.715
+ $X2=0 $Y2=0
cc_1092 N_A_1312_126#_c_1564_n N_VGND_c_2408_n 0.0149545f $X=6.7 $Y=0.86 $X2=0
+ $Y2=0
cc_1093 N_A_2616_417#_c_1689_n N_A_2360_115#_M1031_g 0.00526294f $X=14.66
+ $Y=2.67 $X2=0 $Y2=0
cc_1094 N_A_2616_417#_c_1707_n N_A_2360_115#_M1031_g 0.0299464f $X=15.205
+ $Y=1.26 $X2=0 $Y2=0
cc_1095 N_A_2616_417#_c_1708_n N_A_2360_115#_M1031_g 0.00153054f $X=14.745
+ $Y=1.26 $X2=0 $Y2=0
cc_1096 N_A_2616_417#_c_1690_n N_A_2360_115#_M1031_g 0.00979817f $X=15.37
+ $Y=1.115 $X2=0 $Y2=0
cc_1097 N_A_2616_417#_c_1696_n N_A_2360_115#_M1028_g 4.29417e-19 $X=14.66
+ $Y=2.925 $X2=0 $Y2=0
cc_1098 N_A_2616_417#_c_1689_n N_A_2360_115#_M1028_g 0.00316641f $X=14.66
+ $Y=2.67 $X2=0 $Y2=0
cc_1099 N_A_2616_417#_c_1698_n N_A_2360_115#_M1028_g 5.12014e-19 $X=14.62
+ $Y=2.755 $X2=0 $Y2=0
cc_1100 N_A_2616_417#_c_1693_n N_A_2360_115#_c_1796_n 0.00310954f $X=13.405
+ $Y=2.585 $X2=0 $Y2=0
cc_1101 N_A_2616_417#_c_1694_n N_A_2360_115#_c_1796_n 0.0136032f $X=13.545
+ $Y=2.05 $X2=0 $Y2=0
cc_1102 N_A_2616_417#_M1021_g N_A_2360_115#_c_1796_n 0.00450905f $X=13.48
+ $Y=1.115 $X2=0 $Y2=0
cc_1103 N_A_2616_417#_M1039_g N_A_2360_115#_c_1798_n 0.0169362f $X=13.33
+ $Y=2.925 $X2=0 $Y2=0
cc_1104 N_A_2616_417#_c_1693_n N_A_2360_115#_c_1798_n 0.0126059f $X=13.405
+ $Y=2.585 $X2=0 $Y2=0
cc_1105 N_A_2616_417#_c_1694_n N_A_2360_115#_c_1798_n 0.0374031f $X=13.545
+ $Y=2.05 $X2=0 $Y2=0
cc_1106 N_A_2616_417#_c_1751_p N_A_2360_115#_c_1798_n 0.0123662f $X=13.71
+ $Y=2.755 $X2=0 $Y2=0
cc_1107 N_A_2616_417#_M1039_g N_A_2360_115#_c_1799_n 0.018418f $X=13.33 $Y=2.925
+ $X2=0 $Y2=0
cc_1108 N_A_2616_417#_c_1693_n N_A_2360_115#_c_1799_n 4.73083e-19 $X=13.405
+ $Y=2.585 $X2=0 $Y2=0
cc_1109 N_A_2616_417#_c_1695_n N_A_2360_115#_c_1799_n 0.0352242f $X=14.495
+ $Y=2.755 $X2=0 $Y2=0
cc_1110 N_A_2616_417#_c_1751_p N_A_2360_115#_c_1799_n 0.0189511f $X=13.71
+ $Y=2.755 $X2=0 $Y2=0
cc_1111 N_A_2616_417#_c_1696_n N_A_2360_115#_c_1799_n 0.0115828f $X=14.66
+ $Y=2.925 $X2=0 $Y2=0
cc_1112 N_A_2616_417#_M1039_g N_A_2360_115#_c_1800_n 0.00324687f $X=13.33
+ $Y=2.925 $X2=0 $Y2=0
cc_1113 N_A_2616_417#_M1039_g N_A_2360_115#_c_1801_n 3.97786e-19 $X=13.33
+ $Y=2.925 $X2=0 $Y2=0
cc_1114 N_A_2616_417#_c_1695_n N_A_2360_115#_c_1802_n 0.00465659f $X=14.495
+ $Y=2.755 $X2=0 $Y2=0
cc_1115 N_A_2616_417#_c_1696_n N_A_2360_115#_c_1802_n 0.0180677f $X=14.66
+ $Y=2.925 $X2=0 $Y2=0
cc_1116 N_A_2616_417#_c_1689_n N_A_2360_115#_c_1902_n 0.0123662f $X=14.66
+ $Y=2.67 $X2=0 $Y2=0
cc_1117 N_A_2616_417#_c_1707_n N_A_2360_115#_c_1902_n 0.0151573f $X=15.205
+ $Y=1.26 $X2=0 $Y2=0
cc_1118 N_A_2616_417#_c_1690_n N_A_2360_115#_c_1902_n 0.00296609f $X=15.37
+ $Y=1.115 $X2=0 $Y2=0
cc_1119 N_A_2616_417#_c_1689_n N_A_2360_115#_c_1905_n 0.060919f $X=14.66 $Y=2.67
+ $X2=0 $Y2=0
cc_1120 N_A_2616_417#_c_1696_n N_A_2360_115#_c_1808_n 0.0123388f $X=14.66
+ $Y=2.925 $X2=0 $Y2=0
cc_1121 N_A_2616_417#_c_1698_n N_A_2360_115#_c_1808_n 0.00749745f $X=14.62
+ $Y=2.755 $X2=0 $Y2=0
cc_1122 N_A_2616_417#_c_1690_n N_A_2360_115#_c_1787_n 0.0167535f $X=15.37
+ $Y=1.115 $X2=0 $Y2=0
cc_1123 N_A_2616_417#_c_1689_n N_A_2360_115#_c_1789_n 0.0223091f $X=14.66
+ $Y=2.67 $X2=0 $Y2=0
cc_1124 N_A_2616_417#_c_1690_n N_A_2360_115#_c_1789_n 0.00212715f $X=15.37
+ $Y=1.115 $X2=0 $Y2=0
cc_1125 N_A_2616_417#_c_1690_n N_CLK_c_1958_n 0.00164654f $X=15.37 $Y=1.115
+ $X2=0 $Y2=0
cc_1126 N_A_2616_417#_c_1695_n N_VPWR_M1039_d 0.00304131f $X=14.495 $Y=2.755
+ $X2=-0.33 $Y2=-0.265
cc_1127 N_A_2616_417#_c_1751_p N_VPWR_M1039_d 8.18519e-19 $X=13.71 $Y=2.755
+ $X2=-0.33 $Y2=-0.265
cc_1128 N_A_2616_417#_M1039_g N_VPWR_c_2211_n 0.014507f $X=13.33 $Y=2.925 $X2=0
+ $Y2=0
cc_1129 N_A_2616_417#_c_1695_n N_VPWR_c_2220_n 0.00135862f $X=14.495 $Y=2.755
+ $X2=0 $Y2=0
cc_1130 N_A_2616_417#_c_1696_n N_VPWR_c_2220_n 0.00163907f $X=14.66 $Y=2.925
+ $X2=0 $Y2=0
cc_1131 N_A_2616_417#_M1021_g N_VGND_c_2402_n 0.0554918f $X=13.48 $Y=1.115 $X2=0
+ $Y2=0
cc_1132 N_A_2616_417#_c_1707_n N_VGND_c_2408_n 0.00228453f $X=15.205 $Y=1.26
+ $X2=0 $Y2=0
cc_1133 N_A_2616_417#_c_1708_n N_VGND_c_2408_n 0.00116248f $X=14.745 $Y=1.26
+ $X2=0 $Y2=0
cc_1134 N_A_2616_417#_c_1690_n N_VGND_c_2408_n 0.00215908f $X=15.37 $Y=1.115
+ $X2=0 $Y2=0
cc_1135 N_A_2616_417#_c_1708_n A_2904_181# 0.00168885f $X=14.745 $Y=1.26 $X2=0
+ $Y2=0
cc_1136 N_A_2360_115#_M1031_g N_CLK_c_1958_n 0.00459954f $X=14.98 $Y=1.115 $X2=0
+ $Y2=0
cc_1137 N_A_2360_115#_c_1783_n N_CLK_c_1958_n 0.00326769f $X=17.37 $Y=1.795
+ $X2=0 $Y2=0
cc_1138 N_A_2360_115#_c_1787_n N_CLK_c_1958_n 0.001039f $X=16.685 $Y=1.69 $X2=0
+ $Y2=0
cc_1139 N_A_2360_115#_c_1783_n N_CLK_c_1960_n 0.0422196f $X=17.37 $Y=1.795 $X2=0
+ $Y2=0
cc_1140 N_A_2360_115#_c_1802_n N_CLK_c_1960_n 2.59558e-19 $X=14.925 $Y=3.44
+ $X2=0 $Y2=0
cc_1141 N_A_2360_115#_c_1905_n N_CLK_c_1960_n 0.00131902f $X=15.09 $Y=2.11 $X2=0
+ $Y2=0
cc_1142 N_A_2360_115#_c_1808_n N_CLK_c_1960_n 0.00112809f $X=15.01 $Y=3.355
+ $X2=0 $Y2=0
cc_1143 N_A_2360_115#_c_1787_n N_CLK_c_1960_n 0.0310234f $X=16.685 $Y=1.69 $X2=0
+ $Y2=0
cc_1144 N_A_2360_115#_c_1789_n N_CLK_c_1960_n 0.0382182f $X=15.09 $Y=1.77 $X2=0
+ $Y2=0
cc_1145 N_A_2360_115#_c_1905_n N_CLK_c_1964_n 0.021362f $X=15.09 $Y=2.11 $X2=0
+ $Y2=0
cc_1146 N_A_2360_115#_c_1808_n N_CLK_c_1964_n 0.00946801f $X=15.01 $Y=3.355
+ $X2=0 $Y2=0
cc_1147 N_A_2360_115#_c_1787_n N_CLK_c_1964_n 0.0490251f $X=16.685 $Y=1.69 $X2=0
+ $Y2=0
cc_1148 N_A_2360_115#_c_1789_n N_CLK_c_1964_n 0.00634559f $X=15.09 $Y=1.77 $X2=0
+ $Y2=0
cc_1149 N_A_2360_115#_M1029_g N_A_3417_443#_M1017_g 0.0184541f $X=17.62 $Y=2.59
+ $X2=0 $Y2=0
cc_1150 N_A_2360_115#_M1005_g N_A_3417_443#_M1034_g 0.0152868f $X=17.66 $Y=1.075
+ $X2=0 $Y2=0
cc_1151 N_A_2360_115#_M1005_g N_A_3417_443#_c_1997_n 0.00993368f $X=17.66
+ $Y=1.075 $X2=0 $Y2=0
cc_1152 N_A_2360_115#_c_1783_n N_A_3417_443#_c_1997_n 0.00574576f $X=17.37
+ $Y=1.795 $X2=0 $Y2=0
cc_1153 N_A_2360_115#_M1005_g N_A_3417_443#_c_1998_n 0.0201607f $X=17.66
+ $Y=1.075 $X2=0 $Y2=0
cc_1154 N_A_2360_115#_M1005_g N_A_3417_443#_c_1999_n 0.0120523f $X=17.66
+ $Y=1.075 $X2=0 $Y2=0
cc_1155 N_A_2360_115#_c_1784_n N_A_3417_443#_c_1999_n 0.027105f $X=17.64
+ $Y=1.795 $X2=0 $Y2=0
cc_1156 N_A_2360_115#_M1005_g N_A_3417_443#_c_2000_n 0.028171f $X=17.66 $Y=1.075
+ $X2=0 $Y2=0
cc_1157 N_A_2360_115#_M1029_g N_A_3417_443#_c_2005_n 0.0282534f $X=17.62 $Y=2.59
+ $X2=0 $Y2=0
cc_1158 N_A_2360_115#_c_1783_n N_A_3417_443#_c_2005_n 0.00719951f $X=17.37
+ $Y=1.795 $X2=0 $Y2=0
cc_1159 N_A_2360_115#_M1029_g N_A_3417_443#_c_2012_n 0.0156038f $X=17.62 $Y=2.59
+ $X2=0 $Y2=0
cc_1160 N_A_2360_115#_c_1784_n N_A_3417_443#_c_2012_n 0.0189679f $X=17.64
+ $Y=1.795 $X2=0 $Y2=0
cc_1161 N_A_2360_115#_M1005_g N_A_3417_443#_c_2014_n 5.26268e-19 $X=17.66
+ $Y=1.075 $X2=0 $Y2=0
cc_1162 N_A_2360_115#_c_1784_n N_A_3417_443#_c_2014_n 0.0103026f $X=17.64
+ $Y=1.795 $X2=0 $Y2=0
cc_1163 N_A_2360_115#_c_1799_n N_VPWR_M1039_d 0.00703438f $X=14.145 $Y=3.105
+ $X2=-0.33 $Y2=-0.265
cc_1164 N_A_2360_115#_c_1799_n N_VPWR_c_2211_n 0.0515564f $X=14.145 $Y=3.105
+ $X2=0 $Y2=0
cc_1165 N_A_2360_115#_c_1800_n N_VPWR_c_2211_n 0.0126631f $X=13.2 $Y=3.105 $X2=0
+ $Y2=0
cc_1166 N_A_2360_115#_c_1805_n N_VPWR_c_2211_n 0.0122871f $X=14.315 $Y=3.44
+ $X2=0 $Y2=0
cc_1167 N_A_2360_115#_M1028_g N_VPWR_c_2214_n 0.022391f $X=15.05 $Y=2.925 $X2=0
+ $Y2=0
cc_1168 N_A_2360_115#_c_1802_n N_VPWR_c_2214_n 0.0136633f $X=14.925 $Y=3.44
+ $X2=0 $Y2=0
cc_1169 N_A_2360_115#_c_1808_n N_VPWR_c_2214_n 0.0499617f $X=15.01 $Y=3.355
+ $X2=0 $Y2=0
cc_1170 N_A_2360_115#_M1029_g N_VPWR_c_2217_n 0.0493105f $X=17.62 $Y=2.59 $X2=0
+ $Y2=0
cc_1171 N_A_2360_115#_c_1784_n N_VPWR_c_2217_n 0.0013358f $X=17.64 $Y=1.795
+ $X2=0 $Y2=0
cc_1172 N_A_2360_115#_M1036_d N_VPWR_c_2220_n 0.00439715f $X=11.915 $Y=2.715
+ $X2=0 $Y2=0
cc_1173 N_A_2360_115#_M1028_g N_VPWR_c_2220_n 0.005707f $X=15.05 $Y=2.925 $X2=0
+ $Y2=0
cc_1174 N_A_2360_115#_M1029_g N_VPWR_c_2220_n 0.0102369f $X=17.62 $Y=2.59 $X2=0
+ $Y2=0
cc_1175 N_A_2360_115#_c_1799_n N_VPWR_c_2220_n 0.0123133f $X=14.145 $Y=3.105
+ $X2=0 $Y2=0
cc_1176 N_A_2360_115#_c_1800_n N_VPWR_c_2220_n 0.00111759f $X=13.2 $Y=3.105
+ $X2=0 $Y2=0
cc_1177 N_A_2360_115#_c_1802_n N_VPWR_c_2220_n 0.038308f $X=14.925 $Y=3.44 $X2=0
+ $Y2=0
cc_1178 N_A_2360_115#_c_1805_n N_VPWR_c_2220_n 0.00894946f $X=14.315 $Y=3.44
+ $X2=0 $Y2=0
cc_1179 N_A_2360_115#_M1005_g N_VGND_c_2404_n 0.00319778f $X=17.66 $Y=1.075
+ $X2=0 $Y2=0
cc_1180 N_A_2360_115#_M1005_g N_VGND_c_2406_n 0.0359877f $X=17.66 $Y=1.075 $X2=0
+ $Y2=0
cc_1181 N_A_2360_115#_M1005_g N_VGND_c_2408_n 0.0104851f $X=17.66 $Y=1.075 $X2=0
+ $Y2=0
cc_1182 N_A_2360_115#_c_1785_n N_VGND_c_2408_n 0.0307098f $X=11.94 $Y=0.7 $X2=0
+ $Y2=0
cc_1183 N_CLK_c_1958_n N_A_3417_443#_c_1997_n 0.00274083f $X=16.31 $Y=1.095
+ $X2=0 $Y2=0
cc_1184 N_CLK_c_1960_n N_VPWR_c_2214_n 0.0592969f $X=15.975 $Y=2.05 $X2=0 $Y2=0
cc_1185 N_CLK_c_1964_n N_VPWR_c_2214_n 0.0545199f $X=15.975 $Y=2.05 $X2=0 $Y2=0
cc_1186 N_CLK_c_1960_n N_VPWR_c_2220_n 0.00922818f $X=15.975 $Y=2.05 $X2=0 $Y2=0
cc_1187 N_CLK_c_1958_n N_VGND_c_2404_n 0.0369663f $X=16.31 $Y=1.095 $X2=0 $Y2=0
cc_1188 N_CLK_c_1958_n N_VGND_c_2408_n 0.0128107f $X=16.31 $Y=1.095 $X2=0 $Y2=0
cc_1189 N_A_3417_443#_M1017_g N_VPWR_c_2217_n 0.0816444f $X=18.515 $Y=2.965
+ $X2=0 $Y2=0
cc_1190 N_A_3417_443#_c_1999_n N_VPWR_c_2217_n 0.0419017f $X=18.45 $Y=1.65 $X2=0
+ $Y2=0
cc_1191 N_A_3417_443#_c_2012_n N_VPWR_c_2217_n 0.0640256f $X=17.307 $Y=2.305
+ $X2=0 $Y2=0
cc_1192 N_A_3417_443#_M1017_g N_VPWR_c_2220_n 0.00915578f $X=18.515 $Y=2.965
+ $X2=0 $Y2=0
cc_1193 N_A_3417_443#_c_2005_n N_VPWR_c_2220_n 0.0206348f $X=17.23 $Y=2.39 $X2=0
+ $Y2=0
cc_1194 N_A_3417_443#_M1017_g N_Q_c_2350_n 0.00855732f $X=18.515 $Y=2.965 $X2=0
+ $Y2=0
cc_1195 N_A_3417_443#_M1034_g N_Q_c_2350_n 0.0343925f $X=18.535 $Y=0.91 $X2=0
+ $Y2=0
cc_1196 N_A_3417_443#_c_1999_n N_Q_c_2350_n 0.0234288f $X=18.45 $Y=1.65 $X2=0
+ $Y2=0
cc_1197 N_A_3417_443#_c_1997_n N_VGND_c_2404_n 0.0118649f $X=17.38 $Y=0.95 $X2=0
+ $Y2=0
cc_1198 N_A_3417_443#_M1034_g N_VGND_c_2406_n 0.054682f $X=18.535 $Y=0.91 $X2=0
+ $Y2=0
cc_1199 N_A_3417_443#_c_1997_n N_VGND_c_2406_n 0.0194896f $X=17.38 $Y=0.95 $X2=0
+ $Y2=0
cc_1200 N_A_3417_443#_c_1998_n N_VGND_c_2406_n 0.0166239f $X=17.465 $Y=1.485
+ $X2=0 $Y2=0
cc_1201 N_A_3417_443#_c_1999_n N_VGND_c_2406_n 0.0705716f $X=18.45 $Y=1.65 $X2=0
+ $Y2=0
cc_1202 N_A_3417_443#_c_2000_n N_VGND_c_2406_n 5.8898e-19 $X=18.45 $Y=1.65 $X2=0
+ $Y2=0
cc_1203 N_A_3417_443#_M1034_g N_VGND_c_2408_n 0.00982681f $X=18.535 $Y=0.91
+ $X2=0 $Y2=0
cc_1204 N_A_3417_443#_c_1997_n N_VGND_c_2408_n 0.0227043f $X=17.38 $Y=0.95 $X2=0
+ $Y2=0
cc_1205 N_A_65_649#_c_2058_n A_222_649# 0.00124452f $X=2.56 $Y=3.19 $X2=0 $Y2=0
cc_1206 N_A_65_649#_c_2058_n N_VPWR_M1011_d 0.00183917f $X=2.56 $Y=3.19 $X2=0
+ $Y2=0
cc_1207 N_A_65_649#_c_2058_n N_VPWR_c_2199_n 0.0497043f $X=2.56 $Y=3.19 $X2=0
+ $Y2=0
cc_1208 N_A_65_649#_c_2127_n N_VPWR_c_2199_n 0.00455517f $X=2.645 $Y=3.535 $X2=0
+ $Y2=0
cc_1209 N_A_65_649#_c_2062_n N_VPWR_c_2199_n 0.00992085f $X=2.73 $Y=3.62 $X2=0
+ $Y2=0
cc_1210 N_A_65_649#_c_2059_n N_VPWR_c_2202_n 0.00891252f $X=3.385 $Y=3.62 $X2=0
+ $Y2=0
cc_1211 N_A_65_649#_c_2065_n N_VPWR_c_2202_n 0.00584887f $X=3.47 $Y=3.455 $X2=0
+ $Y2=0
cc_1212 N_A_65_649#_c_2066_n N_VPWR_c_2202_n 0.055498f $X=4.805 $Y=3.14 $X2=0
+ $Y2=0
cc_1213 N_A_65_649#_c_2099_n N_VPWR_c_2202_n 0.0103831f $X=4.89 $Y=3.635 $X2=0
+ $Y2=0
cc_1214 N_A_65_649#_c_2071_n N_VPWR_c_2202_n 0.00403448f $X=4.975 $Y=3.72 $X2=0
+ $Y2=0
cc_1215 N_A_65_649#_M1037_d N_VPWR_c_2220_n 0.00269567f $X=3.33 $Y=3.245 $X2=0
+ $Y2=0
cc_1216 N_A_65_649#_M1026_s N_VPWR_c_2220_n 0.00221032f $X=5.775 $Y=3.205 $X2=0
+ $Y2=0
cc_1217 N_A_65_649#_c_2055_n N_VPWR_c_2220_n 0.044402f $X=0.47 $Y=3.455 $X2=0
+ $Y2=0
cc_1218 N_A_65_649#_c_2058_n N_VPWR_c_2220_n 0.0684221f $X=2.56 $Y=3.19 $X2=0
+ $Y2=0
cc_1219 N_A_65_649#_c_2127_n N_VPWR_c_2220_n 0.00819962f $X=2.645 $Y=3.535 $X2=0
+ $Y2=0
cc_1220 N_A_65_649#_c_2059_n N_VPWR_c_2220_n 0.0329925f $X=3.385 $Y=3.62 $X2=0
+ $Y2=0
cc_1221 N_A_65_649#_c_2062_n N_VPWR_c_2220_n 0.00636947f $X=2.73 $Y=3.62 $X2=0
+ $Y2=0
cc_1222 N_A_65_649#_c_2065_n N_VPWR_c_2220_n 0.00833922f $X=3.47 $Y=3.455 $X2=0
+ $Y2=0
cc_1223 N_A_65_649#_c_2066_n N_VPWR_c_2220_n 0.0208558f $X=4.805 $Y=3.14 $X2=0
+ $Y2=0
cc_1224 N_A_65_649#_c_2099_n N_VPWR_c_2220_n 0.0136995f $X=4.89 $Y=3.635 $X2=0
+ $Y2=0
cc_1225 N_A_65_649#_c_2068_n N_VPWR_c_2220_n 0.0370252f $X=5.755 $Y=3.72 $X2=0
+ $Y2=0
cc_1226 N_A_65_649#_c_2071_n N_VPWR_c_2220_n 0.00701739f $X=4.975 $Y=3.72 $X2=0
+ $Y2=0
cc_1227 N_A_65_649#_c_2075_n N_VPWR_c_2220_n 0.0273006f $X=5.92 $Y=3.415 $X2=0
+ $Y2=0
cc_1228 N_A_65_649#_c_2058_n A_524_649# 3.33862e-19 $X=2.56 $Y=3.19 $X2=0 $Y2=0
cc_1229 N_A_65_649#_c_2127_n A_524_649# 0.0034507f $X=2.645 $Y=3.535 $X2=0 $Y2=0
cc_1230 N_A_65_649#_c_2059_n A_524_649# 7.156e-19 $X=3.385 $Y=3.62 $X2=0 $Y2=0
cc_1231 N_A_65_649#_c_2091_n N_noxref_23_c_2364_n 0.00360596f $X=1.38 $Y=1.69
+ $X2=0 $Y2=0
cc_1232 N_A_65_649#_c_2122_n N_noxref_23_c_2364_n 0.0150102f $X=1.465 $Y=0.765
+ $X2=0 $Y2=0
cc_1233 N_A_65_649#_c_2122_n N_noxref_23_c_2365_n 0.0109639f $X=1.465 $Y=0.765
+ $X2=0.24 $Y2=0
cc_1234 N_A_65_649#_c_2049_n N_noxref_23_c_2365_n 0.0667869f $X=2.32 $Y=0.82
+ $X2=0.24 $Y2=0
cc_1235 N_A_65_649#_c_2049_n noxref_24 0.00392319f $X=2.32 $Y=0.82 $X2=0 $Y2=0
cc_1236 N_A_65_649#_c_2122_n N_VGND_c_2408_n 0.0117813f $X=1.465 $Y=0.765 $X2=0
+ $Y2=0
cc_1237 N_A_65_649#_c_2049_n N_VGND_c_2408_n 0.0356958f $X=2.32 $Y=0.82 $X2=0
+ $Y2=0
cc_1238 N_A_65_649#_c_2050_n N_VGND_c_2408_n 0.0234009f $X=5.88 $Y=0.88 $X2=0
+ $Y2=0
cc_1239 A_222_649# N_VPWR_c_2220_n 0.00203998f $X=1.11 $Y=3.245 $X2=0 $Y2=0
cc_1240 N_VPWR_c_2220_n A_524_649# 0.00421212f $X=18.545 $Y=3.59 $X2=0 $Y2=3.985
cc_1241 N_VPWR_c_2205_n A_1468_641# 0.00218426f $X=8.19 $Y=3.5 $X2=0 $Y2=3.985
cc_1242 N_VPWR_c_2220_n A_1468_641# 5.8829e-19 $X=18.545 $Y=3.59 $X2=0 $Y2=3.985
cc_1243 N_VPWR_c_2220_n N_Q_M1017_d 0.00221032f $X=18.545 $Y=3.59 $X2=0 $Y2=0
cc_1244 N_VPWR_c_2217_n N_Q_c_2350_n 0.0677949f $X=18.125 $Y=2.34 $X2=9.6
+ $Y2=4.07
cc_1245 N_VPWR_c_2220_n N_Q_c_2350_n 0.035852f $X=18.545 $Y=3.59 $X2=9.6
+ $Y2=4.07
cc_1246 N_Q_c_2350_n N_VGND_c_2406_n 0.0335266f $X=18.925 $Y=0.68 $X2=0 $Y2=0
cc_1247 N_Q_M1034_d N_VGND_c_2408_n 0.00137624f $X=18.785 $Y=0.535 $X2=0 $Y2=0
cc_1248 N_Q_c_2350_n N_VGND_c_2408_n 0.0257233f $X=18.925 $Y=0.68 $X2=0 $Y2=0
cc_1249 N_noxref_23_c_2365_n N_VGND_c_2396_n 0.00433879f $X=3.645 $Y=0.35 $X2=0
+ $Y2=0
cc_1250 N_noxref_23_c_2369_n N_VGND_c_2396_n 0.0397171f $X=3.81 $Y=0.84 $X2=0
+ $Y2=0
cc_1251 N_noxref_23_c_2364_n N_VGND_c_2408_n 0.0253432f $X=0.83 $Y=0.84 $X2=0
+ $Y2=0
cc_1252 N_noxref_23_c_2365_n N_VGND_c_2408_n 0.11466f $X=3.645 $Y=0.35 $X2=0
+ $Y2=0
cc_1253 N_noxref_23_c_2367_n N_VGND_c_2408_n 0.0125579f $X=0.995 $Y=0.35 $X2=0
+ $Y2=0
cc_1254 N_noxref_23_c_2369_n N_VGND_c_2408_n 0.0209762f $X=3.81 $Y=0.84 $X2=0
+ $Y2=0
cc_1255 N_VGND_c_2398_n A_1610_126# 0.00573988f $X=8.23 $Y=0.48 $X2=0 $Y2=0
cc_1256 N_VGND_c_2402_n A_2539_181# 0.00707963f $X=13.2 $Y=0.48 $X2=0 $Y2=0
