* File: sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1.spice
* Created: Wed Sep  2 09:07:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1.pex.spice"
.subckt sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1  VNB VPB LVPWR SLEEP_B A X
+ VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* SLEEP_B	SLEEP_B
* LVPWR	LVPWR
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_241_1225#_M1009_g N_A_553_1225#_M1009_s N_VNB_M1009_b
+ NSHORT L=0.15 W=0.74 AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=11.34 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1000 N_A_241_1225#_M1000_d N_A_M1000_g N_VGND_M1000_s N_VNB_M1009_b NSHORT
+ L=0.15 W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1
+ R=4.93333 SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_229_967#_M1010_g N_X_M1010_s N_VNB_M1009_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1001 N_A_188_1293#_M1001_d N_A_241_1225#_M1001_g N_A_176_993#_M1001_s
+ N_VNB_M1009_b NHV L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1
+ R=2 SA=250000 SB=250002 A=0.5 P=3 MULT=1
MM1005 N_A_188_1293#_M1005_d N_A_241_1225#_M1005_g N_A_176_993#_M1001_s
+ N_VNB_M1009_b NHV L=0.5 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1
+ R=2 SA=250001 SB=250002 A=0.5 P=3 MULT=1
MM1004 N_A_188_1293#_M1005_d N_A_553_1225#_M1004_g N_A_229_967#_M1004_s
+ N_VNB_M1009_b NHV L=0.5 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1
+ R=2 SA=250002 SB=250001 A=0.5 P=3 MULT=1
MM1008 N_VGND_M1008_d N_A_507_107#_M1008_g N_A_176_993#_M1008_s N_VNB_M1009_b
+ NHV L=0.8 W=1 AD=0.183571 AS=0.265 PD=1.53143 PS=2.53 NRD=0 NRS=0 M=1 R=1.25
+ SA=400000 SB=400000 A=0.8 P=3.6 MULT=1
MM1012 N_A_188_1293#_M1012_d N_A_553_1225#_M1012_g N_A_229_967#_M1004_s
+ N_VNB_M1009_b NHV L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1
+ R=2 SA=250002 SB=250000 A=0.5 P=3 MULT=1
MM1011 N_A_507_107#_M1011_d N_SLEEP_B_M1011_g N_VGND_M1008_d N_VNB_M1009_b NHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.137679 PD=2.03 PS=1.14857 NRD=0 NRS=9.3708 M=1
+ R=1.5 SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1003 N_A_188_1293#_M1003_d N_SLEEP_B_M1003_g N_VGND_M1003_s N_VNB_M1009_b NHV
+ L=0.6 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 M=1 R=8.33333 SA=300000
+ SB=300001 A=3 P=11.2 MULT=1
MM1016 N_A_188_1293#_M1016_d N_SLEEP_B_M1016_g N_VGND_M1003_s N_VNB_M1009_b NHV
+ L=0.6 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 M=1 R=8.33333 SA=300001
+ SB=300000 A=3 P=11.2 MULT=1
MM1002 N_LVPWR_M1002_d N_A_241_1225#_M1002_g N_A_553_1225#_M1002_s
+ N_LVPWR_M1002_b PHIGHVT L=0.15 W=1.12 AD=0.3864 AS=0.3304 PD=2.93 PS=2.83
+ NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75000.2 SB=75000.3 A=0.168 P=2.54
+ MULT=1
MM1013 N_A_241_1225#_M1013_d N_A_M1013_g N_LVPWR_M1013_s N_LVPWR_M1002_b PHIGHVT
+ L=0.15 W=1.12 AD=0.3304 AS=0.3864 PD=2.83 PS=2.93 NRD=1.7533 NRS=10.5395 M=1
+ R=7.46667 SA=75000.3 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1007_d N_A_229_967#_M1007_g N_X_M1007_s N_VPB_M1014_b PHV L=0.5
+ W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1014 N_VPWR_M1014_d N_A_229_967#_M1014_g N_A_176_993#_M1014_s N_VPB_M1014_b
+ PHV L=2 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.21
+ SA=999999 SB=1e+06 A=0.84 P=4.84 MULT=1
MM1015 N_A_507_107#_M1015_d N_SLEEP_B_M1015_g N_VPWR_M1015_s N_VPB_M1014_b PHV
+ L=0.5 W=1.5 AD=0.3975 AS=0.3975 PD=3.53 PS=3.53 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
MM1006 N_A_229_967#_M1006_d N_A_176_993#_M1006_g N_VPWR_M1014_d N_VPB_M1014_b
+ PHV L=2 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.21
+ SA=1e+06 SB=999999 A=0.84 P=4.84 MULT=1
DX17_noxref N_VNB_M1009_b N_VPB_M1014_b NWDIODE A=25.2149 P=21.44
DX18_noxref N_VNB_M1009_b N_LVPWR_M1002_b NWDIODE A=7.371 P=11.74
*
.include "sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1.pxi.spice"
*
.ends
*
*
