* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_2539_181# a_1212_100# a_2360_115# VNB nhv w=420000u l=500000u
+  ad=2.247e+11p pd=1.91e+06u as=2.5995e+11p ps=2.29e+06u
M1001 a_1468_126# a_1212_471# a_1312_126# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1002 a_294_126# SCD a_137_126# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=2.373e+11p ps=2.81e+06u
M1003 a_1468_641# a_1212_100# a_1312_126# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=2.373e+11p ps=2.81e+06u
M1004 a_137_126# D a_592_126# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1005 VGND a_2360_115# a_3417_443# VNB nhv w=420000u l=500000u
+  ad=9.8655e+11p pd=1.017e+07u as=1.197e+11p ps=1.41e+06u
M1006 a_2616_417# RESET_B VPWR VPB phv w=420000u l=500000u
+  ad=1.176e+11p pd=1.4e+06u as=1.9878e+12p ps=1.661e+07u
M1007 a_1510_100# a_1312_126# VGND VNB nhv w=750000u l=500000u
+  ad=2.1e+11p pd=2.06e+06u as=0p ps=0u
M1008 a_222_649# a_116_451# a_65_649# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=3.57e+11p ps=4.22e+06u
M1009 a_1510_100# a_1312_126# VPWR VPB phv w=1e+06u l=500000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1010 a_1610_126# a_1510_100# a_1468_126# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1011 VPWR SCD a_222_649# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_116_451# SCE VGND VNB nhv w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 VGND RESET_B a_1610_126# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_116_451# SCE VPWR VPB phv w=420000u l=500000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1015 VPWR a_1510_100# a_1468_641# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_65_649# SCE a_294_126# VNB nhv w=420000u l=500000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1017 Q a_3417_443# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=0p ps=0u
M1018 a_1212_100# CLK VPWR VPB phv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
M1019 VPWR RESET_B a_65_649# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_1212_100# a_1212_471# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u
M1021 VGND a_2616_417# a_2539_181# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1312_126# a_1212_100# a_65_649# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_2574_543# a_1212_471# a_2360_115# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=3.912e+11p ps=2.91e+06u
M1024 VGND RESET_B a_137_126# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_2904_181# RESET_B VGND VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1026 a_1312_126# a_1212_471# a_65_649# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1312_126# RESET_B VPWR VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_2360_115# a_2616_417# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_2360_115# a_3417_443# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=2.1375e+11p ps=2.07e+06u
M1030 a_2360_115# a_1212_471# a_1510_100# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_2616_417# a_2360_115# a_2904_181# VNB nhv w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1032 VGND a_1212_100# a_1212_471# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1033 VGND CLK a_1212_100# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1034 Q a_3417_443# VGND VNB nhv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
M1035 a_524_649# SCE VPWR VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1036 a_2360_115# a_1212_100# a_1510_100# VPB phv w=1e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_65_649# D a_524_649# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_592_126# a_116_451# a_65_649# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_2616_417# a_2574_543# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
