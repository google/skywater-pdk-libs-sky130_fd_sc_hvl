* File: sky130_fd_sc_hvl__diode_2.spice
* Created: Fri Aug 28 09:34:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__diode_2.pex.spice"
.subckt sky130_fd_sc_hvl__diode_2  VNB VPB DIODE VGND VPWR
* 
* DIODE	DIODE
* VPB	VPB
* VNB	VNB
D0_noxref N_VNB_D0_noxref_pos N_DIODE_D0_noxref_neg NDIODE_H  AREA=0.6072
+ PJ=3.16 M=1 AHFTEMPPERIM=3.16
DX1_noxref N_VNB_D0_noxref_pos N_VPB_X1_noxref_D1 NWDIODE A=4.212 P=8.44
*
.include "sky130_fd_sc_hvl__diode_2.pxi.spice"
*
.ends
*
*
