* File: sky130_fd_sc_hvl__nor2_1.pxi.spice
* Created: Fri Aug 28 09:38:11 2020
* 
x_PM_SKY130_FD_SC_HVL__NOR2_1%VNB N_VNB_M1002_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__NOR2_1%VNB
x_PM_SKY130_FD_SC_HVL__NOR2_1%VPB N_VPB_M1000_b VPB N_VPB_c_21_p VPB
+ PM_SKY130_FD_SC_HVL__NOR2_1%VPB
x_PM_SKY130_FD_SC_HVL__NOR2_1%A N_A_M1002_g N_A_M1000_g A A A N_A_c_39_n
+ PM_SKY130_FD_SC_HVL__NOR2_1%A
x_PM_SKY130_FD_SC_HVL__NOR2_1%B B N_B_M1003_g N_B_c_70_n N_B_M1001_g
+ PM_SKY130_FD_SC_HVL__NOR2_1%B
x_PM_SKY130_FD_SC_HVL__NOR2_1%VPWR N_VPWR_M1000_s VPWR N_VPWR_c_85_n
+ N_VPWR_c_88_n PM_SKY130_FD_SC_HVL__NOR2_1%VPWR
x_PM_SKY130_FD_SC_HVL__NOR2_1%Y N_Y_M1002_d N_Y_M1001_d N_Y_c_103_n N_Y_c_105_n
+ N_Y_c_106_n Y Y Y Y Y N_Y_c_107_n Y PM_SKY130_FD_SC_HVL__NOR2_1%Y
x_PM_SKY130_FD_SC_HVL__NOR2_1%VGND N_VGND_M1002_s N_VGND_M1003_d VGND
+ N_VGND_c_132_n N_VGND_c_134_n N_VGND_c_136_n PM_SKY130_FD_SC_HVL__NOR2_1%VGND
cc_1 N_VNB_M1002_b N_A_M1002_g 0.0481897f $X=-0.33 $Y=-0.265 $X2=0.935 $Y2=0.91
cc_2 N_VNB_c_2_p N_A_M1002_g 7.72665e-19 $X=0.24 $Y=0 $X2=0.935 $Y2=0.91
cc_3 N_VNB_M1002_b A 0.0150288f $X=-0.33 $Y=-0.265 $X2=1.115 $Y2=1.95
cc_4 N_VNB_M1002_b N_A_c_39_n 0.0594534f $X=-0.33 $Y=-0.265 $X2=0.91 $Y2=1.89
cc_5 N_VNB_M1002_b N_B_M1003_g 0.0941342f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_c_2_p N_B_M1003_g 0.00119158f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_7 N_VNB_M1002_b N_Y_c_103_n 0.0121798f $X=-0.33 $Y=-0.265 $X2=0.155 $Y2=1.95
cc_8 N_VNB_c_2_p N_Y_c_103_n 9.05583e-19 $X=0.24 $Y=0 $X2=0.155 $Y2=1.95
cc_9 N_VNB_M1002_b N_Y_c_105_n 0.00235986f $X=-0.33 $Y=-0.265 $X2=1.115 $Y2=1.95
cc_10 N_VNB_M1002_b N_Y_c_106_n 0.00668365f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_11 N_VNB_M1002_b N_Y_c_107_n 0.0101781f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_12 N_VNB_M1002_b Y 0.0147008f $X=-0.33 $Y=-0.265 $X2=1.2 $Y2=1.947
cc_13 N_VNB_M1002_b N_VGND_c_132_n 0.0984979f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.95
cc_14 N_VNB_c_2_p N_VGND_c_132_n 0.00263373f $X=0.24 $Y=0 $X2=0.635 $Y2=1.95
cc_15 N_VNB_M1002_b N_VGND_c_134_n 0.0614087f $X=-0.33 $Y=-0.265 $X2=0.97
+ $Y2=2.085
cc_16 N_VNB_c_2_p N_VGND_c_134_n 0.00166879f $X=0.24 $Y=0 $X2=0.97 $Y2=2.085
cc_17 N_VNB_M1002_b N_VGND_c_136_n 0.0590711f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=1.947
cc_18 N_VNB_c_2_p N_VGND_c_136_n 0.256627f $X=0.24 $Y=0 $X2=0.24 $Y2=1.947
cc_19 N_VPB_M1000_b N_A_M1000_g 0.0408865f $X=-0.33 $Y=1.885 $X2=1.005 $Y2=2.965
cc_20 VPB N_A_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=1.005 $Y2=2.965
cc_21 N_VPB_c_21_p N_A_M1000_g 0.0137101f $X=2.16 $Y=4.07 $X2=1.005 $Y2=2.965
cc_22 N_VPB_M1000_b A 0.0207981f $X=-0.33 $Y=1.885 $X2=1.115 $Y2=1.95
cc_23 N_VPB_M1000_b N_A_c_39_n 0.0218389f $X=-0.33 $Y=1.885 $X2=0.91 $Y2=1.89
cc_24 N_VPB_M1000_b N_B_M1003_g 0.0572902f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_25 VPB N_B_M1003_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_26 N_VPB_c_21_p N_B_M1003_g 0.0161677f $X=2.16 $Y=4.07 $X2=0 $Y2=0
cc_27 N_VPB_M1000_b N_VPWR_c_85_n 0.0797891f $X=-0.33 $Y=1.885 $X2=1.005
+ $Y2=2.965
cc_28 VPB N_VPWR_c_85_n 0.00648924f $X=0 $Y=3.955 $X2=1.005 $Y2=2.965
cc_29 N_VPB_c_21_p N_VPWR_c_85_n 0.0849988f $X=2.16 $Y=4.07 $X2=1.005 $Y2=2.965
cc_30 N_VPB_M1000_b N_VPWR_c_88_n 0.0435745f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_88_n 0.254862f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_32 N_VPB_c_21_p N_VPWR_c_88_n 0.0102076f $X=2.16 $Y=4.07 $X2=0 $Y2=0
cc_33 N_VPB_M1000_b Y 0.0687543f $X=-0.33 $Y=1.885 $X2=1.2 $Y2=1.947
cc_34 VPB Y 7.75439e-19 $X=0 $Y=3.955 $X2=1.2 $Y2=1.947
cc_35 N_VPB_c_21_p Y 0.0133691f $X=2.16 $Y=4.07 $X2=1.2 $Y2=1.947
cc_36 N_A_M1002_g N_B_M1003_g 0.0171153f $X=0.935 $Y=0.91 $X2=0 $Y2=0
cc_37 A N_B_M1003_g 0.00235781f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_38 N_A_c_39_n N_B_M1003_g 0.164107f $X=0.91 $Y=1.89 $X2=0 $Y2=0
cc_39 A N_B_c_70_n 0.0277063f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_40 N_A_c_39_n N_B_c_70_n 3.59121e-19 $X=0.91 $Y=1.89 $X2=0 $Y2=0
cc_41 N_A_M1000_g N_VPWR_c_85_n 0.0931099f $X=1.005 $Y=2.965 $X2=0 $Y2=0
cc_42 A N_VPWR_c_85_n 0.0914751f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_43 N_A_c_39_n N_VPWR_c_85_n 3.29134e-19 $X=0.91 $Y=1.89 $X2=0 $Y2=0
cc_44 N_A_M1000_g N_VPWR_c_88_n 0.00248085f $X=1.005 $Y=2.965 $X2=0 $Y2=0
cc_45 N_A_M1002_g N_Y_c_103_n 0.00418089f $X=0.935 $Y=0.91 $X2=0 $Y2=0
cc_46 N_A_c_39_n N_Y_c_103_n 0.00189139f $X=0.91 $Y=1.89 $X2=0 $Y2=0
cc_47 A N_Y_c_106_n 0.0092789f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_48 N_A_c_39_n N_Y_c_106_n 0.0115591f $X=0.91 $Y=1.89 $X2=0 $Y2=0
cc_49 N_A_M1002_g N_VGND_c_132_n 0.0575735f $X=0.935 $Y=0.91 $X2=0.24 $Y2=0
cc_50 A N_VGND_c_132_n 0.0374179f $X=1.115 $Y=1.95 $X2=0.24 $Y2=0
cc_51 N_A_M1002_g N_VGND_c_134_n 7.92123e-19 $X=0.935 $Y=0.91 $X2=0 $Y2=0
cc_52 N_A_M1002_g N_VGND_c_136_n 0.0100067f $X=0.935 $Y=0.91 $X2=0 $Y2=0
cc_53 N_B_M1003_g N_VPWR_c_85_n 0.077604f $X=1.715 $Y=0.91 $X2=0 $Y2=0
cc_54 N_B_c_70_n N_VPWR_c_85_n 0.0202115f $X=1.66 $Y=1.89 $X2=0 $Y2=0
cc_55 N_B_M1003_g N_VPWR_c_88_n 0.0130863f $X=1.715 $Y=0.91 $X2=0 $Y2=0
cc_56 N_B_M1003_g N_Y_c_103_n 0.0271578f $X=1.715 $Y=0.91 $X2=0 $Y2=0
cc_57 N_B_M1003_g N_Y_c_105_n 0.0324609f $X=1.715 $Y=0.91 $X2=0.24 $Y2=0
cc_58 N_B_c_70_n N_Y_c_105_n 0.0201936f $X=1.66 $Y=1.89 $X2=0.24 $Y2=0
cc_59 N_B_M1003_g N_Y_c_106_n 0.00470766f $X=1.715 $Y=0.91 $X2=0 $Y2=0
cc_60 N_B_c_70_n N_Y_c_106_n 0.00261289f $X=1.66 $Y=1.89 $X2=0 $Y2=0
cc_61 N_B_M1003_g Y 0.0261302f $X=1.715 $Y=0.91 $X2=0 $Y2=0
cc_62 N_B_c_70_n Y 0.024131f $X=1.66 $Y=1.89 $X2=0 $Y2=0
cc_63 N_B_M1003_g N_VGND_c_132_n 0.00104764f $X=1.715 $Y=0.91 $X2=0.24 $Y2=0
cc_64 N_B_M1003_g N_VGND_c_134_n 0.0435168f $X=1.715 $Y=0.91 $X2=0 $Y2=0
cc_65 N_B_M1003_g N_VGND_c_136_n 0.0119169f $X=1.715 $Y=0.91 $X2=0 $Y2=0
cc_66 N_VPWR_c_85_n A_251_443# 0.00419528f $X=0.615 $Y=2.385 $X2=0 $Y2=3.985
cc_67 N_VPWR_c_88_n N_Y_M1001_d 0.00221032f $X=1.645 $Y=3.59 $X2=0 $Y2=0
cc_68 N_VPWR_c_85_n Y 0.0446026f $X=0.615 $Y=2.385 $X2=0 $Y2=0
cc_69 N_VPWR_c_88_n Y 0.0369651f $X=1.645 $Y=3.59 $X2=0 $Y2=0
cc_70 N_Y_c_103_n N_VGND_c_132_n 0.0364699f $X=1.325 $Y=0.66 $X2=0.24 $Y2=0
cc_71 N_Y_c_103_n N_VGND_c_134_n 0.0520535f $X=1.325 $Y=0.66 $X2=0 $Y2=0
cc_72 N_Y_c_105_n N_VGND_c_134_n 0.0196695f $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_73 N_Y_c_107_n N_VGND_c_134_n 0.022439f $X=2.147 $Y=1.595 $X2=0 $Y2=0
cc_74 N_Y_M1002_d N_VGND_c_136_n 5.42154e-19 $X=1.185 $Y=0.535 $X2=0 $Y2=0
cc_75 N_Y_c_103_n N_VGND_c_136_n 0.0313616f $X=1.325 $Y=0.66 $X2=0 $Y2=0
