* File: sky130_fd_sc_hvl__or3_1.pxi.spice
* Created: Fri Aug 28 09:39:09 2020
* 
x_PM_SKY130_FD_SC_HVL__OR3_1%VNB N_VNB_M1007_b VNB N_VNB_c_4_p VNB
+ PM_SKY130_FD_SC_HVL__OR3_1%VNB
x_PM_SKY130_FD_SC_HVL__OR3_1%VPB N_VPB_M1002_b VPB N_VPB_c_40_p VPB
+ PM_SKY130_FD_SC_HVL__OR3_1%VPB
x_PM_SKY130_FD_SC_HVL__OR3_1%C N_C_M1002_g N_C_c_52_n C C N_C_M1007_g
+ PM_SKY130_FD_SC_HVL__OR3_1%C
x_PM_SKY130_FD_SC_HVL__OR3_1%B B B B B N_B_M1004_g N_B_c_80_n N_B_M1005_g
+ PM_SKY130_FD_SC_HVL__OR3_1%B
x_PM_SKY130_FD_SC_HVL__OR3_1%A N_A_M1006_g N_A_M1001_g A N_A_c_106_n
+ PM_SKY130_FD_SC_HVL__OR3_1%A
x_PM_SKY130_FD_SC_HVL__OR3_1%A_30_107# N_A_30_107#_M1007_s N_A_30_107#_M1004_d
+ N_A_30_107#_M1002_s N_A_30_107#_M1000_g N_A_30_107#_M1003_g
+ N_A_30_107#_c_135_n N_A_30_107#_c_137_n N_A_30_107#_c_138_n
+ N_A_30_107#_c_139_n N_A_30_107#_c_140_n N_A_30_107#_c_141_n
+ N_A_30_107#_c_142_n N_A_30_107#_c_144_n N_A_30_107#_c_177_n
+ N_A_30_107#_c_145_n PM_SKY130_FD_SC_HVL__OR3_1%A_30_107#
x_PM_SKY130_FD_SC_HVL__OR3_1%VPWR N_VPWR_M1006_d VPWR N_VPWR_c_202_n
+ N_VPWR_c_205_n PM_SKY130_FD_SC_HVL__OR3_1%VPWR
x_PM_SKY130_FD_SC_HVL__OR3_1%X N_X_M1003_d N_X_M1000_d X X X X X X X N_X_c_223_n
+ PM_SKY130_FD_SC_HVL__OR3_1%X
x_PM_SKY130_FD_SC_HVL__OR3_1%VGND N_VGND_M1007_d N_VGND_M1001_d VGND
+ N_VGND_c_237_n N_VGND_c_239_n N_VGND_c_241_n PM_SKY130_FD_SC_HVL__OR3_1%VGND
cc_1 N_VNB_M1007_b N_C_c_52_n 0.0203412f $X=-0.33 $Y=-0.265 $X2=0.682 $Y2=2.19
cc_2 N_VNB_M1007_b C 0.00505959f $X=-0.33 $Y=-0.265 $X2=1.115 $Y2=1.21
cc_3 N_VNB_M1007_b N_C_M1007_g 0.101691f $X=-0.33 $Y=-0.265 $X2=0.665 $Y2=0.745
cc_4 N_VNB_c_4_p N_C_M1007_g 5.39935e-19 $X=0.24 $Y=0 $X2=0.665 $Y2=0.745
cc_5 N_VNB_M1007_b N_B_M1004_g 0.109265f $X=-0.33 $Y=-0.265 $X2=0.695 $Y2=1.235
cc_6 N_VNB_c_4_p N_B_M1004_g 0.00149413f $X=0.24 $Y=0 $X2=0.695 $Y2=1.235
cc_7 N_VNB_M1007_b N_A_M1006_g 0.02702f $X=-0.33 $Y=-0.265 $X2=0.7 $Y2=2.53
cc_8 N_VNB_M1007_b N_A_M1001_g 0.0522359f $X=-0.33 $Y=-0.265 $X2=0.682 $Y2=2.19
cc_9 N_VNB_c_4_p N_A_M1001_g 0.0023273f $X=0.24 $Y=0 $X2=0.682 $Y2=2.19
cc_10 N_VNB_M1007_b A 0.00267816f $X=-0.33 $Y=-0.265 $X2=1.115 $Y2=1.21
cc_11 N_VNB_M1007_b N_A_c_106_n 0.0528401f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=0.745
cc_12 N_VNB_M1007_b N_A_30_107#_M1003_g 0.0465472f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=1.28
cc_13 N_VNB_c_4_p N_A_30_107#_M1003_g 6.33027e-19 $X=0.24 $Y=0 $X2=0.695
+ $Y2=1.28
cc_14 N_VNB_M1007_b N_A_30_107#_c_135_n 0.0510106f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_15 N_VNB_c_4_p N_A_30_107#_c_135_n 4.99172e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_16 N_VNB_M1007_b N_A_30_107#_c_137_n 0.00751173f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_17 N_VNB_M1007_b N_A_30_107#_c_138_n 0.00635317f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1007_b N_A_30_107#_c_139_n 0.004782f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_19 N_VNB_M1007_b N_A_30_107#_c_140_n 0.019791f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_20 N_VNB_M1007_b N_A_30_107#_c_141_n 0.00891503f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_21 N_VNB_M1007_b N_A_30_107#_c_142_n 0.0128585f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_22 N_VNB_c_4_p N_A_30_107#_c_142_n 0.00120764f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_23 N_VNB_M1007_b N_A_30_107#_c_144_n 4.21834e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_24 N_VNB_M1007_b N_A_30_107#_c_145_n 0.0489504f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_25 N_VNB_M1007_b N_X_c_223_n 0.0672092f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_26 N_VNB_c_4_p N_X_c_223_n 5.92913e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_27 N_VNB_M1007_b N_VGND_c_237_n 0.0422668f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_28 N_VNB_c_4_p N_VGND_c_237_n 0.00242936f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_29 N_VNB_M1007_b N_VGND_c_239_n 0.0420549f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=1.28
cc_30 N_VNB_c_4_p N_VGND_c_239_n 0.00189583f $X=0.24 $Y=0 $X2=0.695 $Y2=1.28
cc_31 N_VNB_M1007_b N_VGND_c_241_n 0.079922f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=1.235
cc_32 N_VNB_c_4_p N_VGND_c_241_n 0.41076f $X=0.24 $Y=0 $X2=0.695 $Y2=1.235
cc_33 N_VPB_M1002_b N_C_M1002_g 0.0420873f $X=-0.33 $Y=1.885 $X2=0.7 $Y2=2.53
cc_34 N_VPB_M1002_b N_C_c_52_n 0.0305047f $X=-0.33 $Y=1.885 $X2=0.682 $Y2=2.19
cc_35 N_VPB_M1002_b N_B_M1004_g 0.060615f $X=-0.33 $Y=1.885 $X2=0.695 $Y2=1.235
cc_36 N_VPB_M1002_b N_B_c_80_n 0.0414764f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_37 N_VPB_M1002_b N_A_M1006_g 0.0651284f $X=-0.33 $Y=1.885 $X2=0.7 $Y2=2.53
cc_38 N_VPB_M1002_b N_A_30_107#_M1000_g 0.042585f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=0.745
cc_39 VPB N_A_30_107#_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.665 $Y2=0.745
cc_40 N_VPB_c_40_p N_A_30_107#_M1000_g 0.0152014f $X=3.6 $Y=4.07 $X2=0.665
+ $Y2=0.745
cc_41 N_VPB_M1002_b N_A_30_107#_c_137_n 0.0498671f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_42 N_VPB_M1002_b N_A_30_107#_c_145_n 0.0223978f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_43 N_VPB_M1002_b N_VPWR_c_202_n 0.0577931f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_202_n 0.00574106f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_45 N_VPB_c_40_p N_VPWR_c_202_n 0.0861811f $X=3.6 $Y=4.07 $X2=0 $Y2=0
cc_46 N_VPB_M1002_b N_VPWR_c_205_n 0.0900811f $X=-0.33 $Y=1.885 $X2=0.665
+ $Y2=1.28
cc_47 VPB N_VPWR_c_205_n 0.409802f $X=0 $Y=3.955 $X2=0.665 $Y2=1.28
cc_48 N_VPB_c_40_p N_VPWR_c_205_n 0.0214854f $X=3.6 $Y=4.07 $X2=0.665 $Y2=1.28
cc_49 N_VPB_M1002_b N_X_c_223_n 0.0691995f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_50 VPB N_X_c_223_n 7.75439e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_51 N_VPB_c_40_p N_X_c_223_n 0.0133691f $X=3.6 $Y=4.07 $X2=0 $Y2=0
cc_52 N_C_c_52_n N_B_M1004_g 0.06324f $X=0.682 $Y=2.19 $X2=0 $Y2=0
cc_53 C N_B_M1004_g 0.0152432f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_54 N_C_M1007_g N_B_M1004_g 0.0426103f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_55 N_C_M1002_g N_B_c_80_n 0.0469063f $X=0.7 $Y=2.53 $X2=0 $Y2=0
cc_56 N_C_c_52_n N_B_c_80_n 0.0203766f $X=0.682 $Y=2.19 $X2=0 $Y2=0
cc_57 C N_A_30_107#_c_135_n 0.0250337f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_58 N_C_M1007_g N_A_30_107#_c_135_n 0.023906f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_59 N_C_M1002_g N_A_30_107#_c_137_n 0.00563475f $X=0.7 $Y=2.53 $X2=1.92
+ $Y2=0.058
cc_60 N_C_c_52_n N_A_30_107#_c_137_n 0.0173468f $X=0.682 $Y=2.19 $X2=1.92
+ $Y2=0.058
cc_61 N_C_c_52_n N_A_30_107#_c_138_n 0.0169369f $X=0.682 $Y=2.19 $X2=0 $Y2=0
cc_62 C N_A_30_107#_c_138_n 0.058014f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_63 N_C_M1007_g N_A_30_107#_c_138_n 0.020451f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_64 C N_A_30_107#_c_139_n 0.0172142f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_65 N_C_M1007_g N_A_30_107#_c_139_n 0.00137401f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_66 N_C_M1002_g N_VPWR_c_205_n 0.00388009f $X=0.7 $Y=2.53 $X2=0 $Y2=0
cc_67 C N_VGND_c_237_n 0.0556457f $X=1.115 $Y=1.21 $X2=0.24 $Y2=0
cc_68 N_C_M1007_g N_VGND_c_237_n 0.0358112f $X=0.665 $Y=0.745 $X2=0.24 $Y2=0
cc_69 C N_VGND_c_241_n 0.00315508f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_70 N_C_M1007_g N_VGND_c_241_n 0.00834095f $X=0.665 $Y=0.745 $X2=0 $Y2=0
cc_71 N_B_c_80_n N_A_M1006_g 0.00180227f $X=1.37 $Y=1.995 $X2=0 $Y2=0
cc_72 N_B_M1004_g N_A_M1001_g 0.0139339f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_73 N_B_M1004_g A 3.55802e-19 $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_74 N_B_M1004_g N_A_c_106_n 0.121226f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_75 N_B_c_80_n N_A_30_107#_c_137_n 0.0461722f $X=1.37 $Y=1.995 $X2=1.92
+ $Y2=0.058
cc_76 N_B_M1004_g N_A_30_107#_c_138_n 0.0250656f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_77 N_B_c_80_n N_A_30_107#_c_138_n 0.0696376f $X=1.37 $Y=1.995 $X2=0 $Y2=0
cc_78 N_B_M1004_g N_A_30_107#_c_139_n 0.0225469f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_79 N_B_M1004_g N_A_30_107#_c_142_n 0.0125287f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_80 N_B_M1004_g N_A_30_107#_c_144_n 0.0110608f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_81 N_B_M1004_g N_VPWR_c_202_n 0.00888458f $X=1.455 $Y=0.745 $X2=0.24 $Y2=0
cc_82 N_B_c_80_n N_VPWR_c_202_n 0.0949417f $X=1.37 $Y=1.995 $X2=0.24 $Y2=0
cc_83 N_B_M1004_g N_VPWR_c_205_n 0.00213903f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_84 N_B_c_80_n N_VPWR_c_205_n 0.0524081f $X=1.37 $Y=1.995 $X2=0 $Y2=0
cc_85 N_B_M1004_g N_VGND_c_237_n 0.0236369f $X=1.455 $Y=0.745 $X2=0.24 $Y2=0
cc_86 N_B_M1004_g N_VGND_c_241_n 0.0121164f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_87 N_A_M1001_g N_A_30_107#_M1003_g 0.0176474f $X=2.235 $Y=0.745 $X2=3.6 $Y2=0
cc_88 A N_A_30_107#_M1003_g 4.71551e-19 $X=2.075 $Y=1.21 $X2=3.6 $Y2=0
cc_89 N_A_M1001_g N_A_30_107#_c_139_n 0.00252073f $X=2.235 $Y=0.745 $X2=0 $Y2=0
cc_90 A N_A_30_107#_c_139_n 0.0231404f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A_c_106_n N_A_30_107#_c_139_n 0.00439954f $X=2.08 $Y=1.28 $X2=0 $Y2=0
cc_92 N_A_M1006_g N_A_30_107#_c_140_n 0.0221698f $X=2.165 $Y=2.53 $X2=0 $Y2=0
cc_93 A N_A_30_107#_c_140_n 0.0380144f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_94 N_A_c_106_n N_A_30_107#_c_140_n 0.0119727f $X=2.08 $Y=1.28 $X2=0 $Y2=0
cc_95 N_A_M1001_g N_A_30_107#_c_142_n 0.00100123f $X=2.235 $Y=0.745 $X2=0 $Y2=0
cc_96 A N_A_30_107#_c_142_n 0.00243027f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A_c_106_n N_A_30_107#_c_142_n 2.69323e-19 $X=2.08 $Y=1.28 $X2=0 $Y2=0
cc_98 N_A_M1006_g N_A_30_107#_c_177_n 0.00134711f $X=2.165 $Y=2.53 $X2=0 $Y2=0
cc_99 N_A_M1006_g N_A_30_107#_c_145_n 0.0255522f $X=2.165 $Y=2.53 $X2=0 $Y2=0
cc_100 N_A_c_106_n N_A_30_107#_c_145_n 0.00686574f $X=2.08 $Y=1.28 $X2=0 $Y2=0
cc_101 N_A_M1006_g N_VPWR_c_202_n 0.0762953f $X=2.165 $Y=2.53 $X2=0.24 $Y2=0
cc_102 N_A_c_106_n N_VPWR_c_202_n 3.75842e-19 $X=2.08 $Y=1.28 $X2=0.24 $Y2=0
cc_103 N_A_M1001_g N_VGND_c_237_n 6.41433e-19 $X=2.235 $Y=0.745 $X2=0.24 $Y2=0
cc_104 N_A_M1001_g N_VGND_c_239_n 0.0164219f $X=2.235 $Y=0.745 $X2=3.6 $Y2=0
cc_105 A N_VGND_c_239_n 0.0212163f $X=2.075 $Y=1.21 $X2=3.6 $Y2=0
cc_106 N_A_M1001_g N_VGND_c_241_n 0.0203243f $X=2.235 $Y=0.745 $X2=0 $Y2=0
cc_107 A N_VGND_c_241_n 0.0161687f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_108 N_A_30_107#_M1000_g N_VPWR_c_202_n 0.0809107f $X=3.155 $Y=2.965 $X2=0.24
+ $Y2=0
cc_109 N_A_30_107#_c_140_n N_VPWR_c_202_n 0.0471327f $X=2.925 $Y=1.645 $X2=0.24
+ $Y2=0
cc_110 N_A_30_107#_c_144_n N_VPWR_c_202_n 0.00143827f $X=1.65 $Y=1.645 $X2=0.24
+ $Y2=0
cc_111 N_A_30_107#_c_177_n N_VPWR_c_202_n 0.0201091f $X=3.09 $Y=1.645 $X2=0.24
+ $Y2=0
cc_112 N_A_30_107#_M1000_g N_VPWR_c_205_n 0.00911082f $X=3.155 $Y=2.965 $X2=0
+ $Y2=0
cc_113 N_A_30_107#_M1000_g N_X_c_223_n 0.00855437f $X=3.155 $Y=2.965 $X2=0 $Y2=0
cc_114 N_A_30_107#_M1003_g N_X_c_223_n 0.0335968f $X=3.175 $Y=0.91 $X2=0 $Y2=0
cc_115 N_A_30_107#_c_177_n N_X_c_223_n 0.0252666f $X=3.09 $Y=1.645 $X2=0 $Y2=0
cc_116 N_A_30_107#_c_135_n N_VGND_c_237_n 0.0192182f $X=0.275 $Y=0.745 $X2=0.24
+ $Y2=0
cc_117 N_A_30_107#_c_138_n N_VGND_c_237_n 0.00168196f $X=1.565 $Y=1.645 $X2=0.24
+ $Y2=0
cc_118 N_A_30_107#_c_142_n N_VGND_c_237_n 0.0299404f $X=1.845 $Y=0.745 $X2=0.24
+ $Y2=0
cc_119 N_A_30_107#_M1003_g N_VGND_c_239_n 0.0566305f $X=3.175 $Y=0.91 $X2=3.6
+ $Y2=0
cc_120 N_A_30_107#_c_140_n N_VGND_c_239_n 0.0203787f $X=2.925 $Y=1.645 $X2=3.6
+ $Y2=0
cc_121 N_A_30_107#_c_142_n N_VGND_c_239_n 0.00606729f $X=1.845 $Y=0.745 $X2=3.6
+ $Y2=0
cc_122 N_A_30_107#_c_177_n N_VGND_c_239_n 0.0204526f $X=3.09 $Y=1.645 $X2=3.6
+ $Y2=0
cc_123 N_A_30_107#_c_145_n N_VGND_c_239_n 6.24206e-19 $X=3.09 $Y=1.77 $X2=3.6
+ $Y2=0
cc_124 N_A_30_107#_M1007_s N_VGND_c_241_n 0.00221032f $X=0.15 $Y=0.535 $X2=0
+ $Y2=0
cc_125 N_A_30_107#_M1004_d N_VGND_c_241_n 2.20496e-19 $X=1.705 $Y=0.535 $X2=0
+ $Y2=0
cc_126 N_A_30_107#_M1003_g N_VGND_c_241_n 0.00925078f $X=3.175 $Y=0.91 $X2=0
+ $Y2=0
cc_127 N_A_30_107#_c_135_n N_VGND_c_241_n 0.0233307f $X=0.275 $Y=0.745 $X2=0
+ $Y2=0
cc_128 N_A_30_107#_c_139_n N_VGND_c_241_n 5.47712e-19 $X=1.65 $Y=1.56 $X2=0
+ $Y2=0
cc_129 N_A_30_107#_c_142_n N_VGND_c_241_n 0.0287622f $X=1.845 $Y=0.745 $X2=0
+ $Y2=0
cc_130 N_VPWR_c_205_n N_X_M1000_d 0.00221032f $X=3.195 $Y=3.59 $X2=0 $Y2=0
cc_131 N_VPWR_c_202_n N_X_c_223_n 0.0681201f $X=1.755 $Y=3.59 $X2=1.92 $Y2=4.07
cc_132 N_VPWR_c_205_n N_X_c_223_n 0.0358369f $X=3.195 $Y=3.59 $X2=1.92 $Y2=4.07
cc_133 N_X_c_223_n N_VGND_c_239_n 0.0381137f $X=3.565 $Y=0.68 $X2=3.6 $Y2=0
cc_134 N_X_M1003_d N_VGND_c_241_n 0.00137624f $X=3.425 $Y=0.535 $X2=0 $Y2=0
cc_135 N_X_c_223_n N_VGND_c_241_n 0.0267201f $X=3.565 $Y=0.68 $X2=0 $Y2=0
