* File: sky130_fd_sc_hvl__sdfstp_1.pex.spice
* Created: Fri Aug 28 09:40:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%VNB 5 7 11
c122 11 0 1.2102e-19 $X=0.24 $Y=0
r123 7 11 0.000380609 $w=1.872e-05 $l=5.7e-08 $layer=MET1_cond $X=9.36 $Y=0.057
+ $X2=9.36 $Y2=0
r124 5 11 0.476923 $w=1.7e-07 $l=3.315e-06 $layer=mcon $count=19 $X=18.48 $Y=0
+ $X2=18.48 $Y2=0
r125 5 11 0.476923 $w=1.7e-07 $l=3.315e-06 $layer=mcon $count=19 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%VPB 4 6 14
c162 4 0 1.02273e-19 $X=-0.33 $Y=1.885
r163 10 14 0.476923 $w=1.7e-07 $l=3.315e-06 $layer=mcon $count=19 $X=18.48
+ $Y=4.07 $X2=18.48 $Y2=4.07
r164 9 14 1189.99 $w=1.68e-07 $l=1.824e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=18.48 $Y2=4.07
r165 9 10 0.476923 $w=1.7e-07 $l=3.315e-06 $layer=mcon $count=19 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r166 6 10 0.000380609 $w=1.872e-05 $l=5.7e-08 $layer=MET1_cond $X=9.36 $Y=4.013
+ $X2=9.36 $Y2=4.07
r167 4 14 9.33333 $w=1.7e-07 $l=1.85225e-05 $layer=licon1_NTAP_notbjt $count=19
+ $X=0 $Y=3.985 $X2=18.48 $Y2=4.07
r168 4 9 9.33333 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=19
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%SCE 1 3 4 6 9 10 15 18 20 21 25 29 30 31
c65 29 0 1.88256e-19 $X=2.8 $Y=1.26
r66 29 31 18.3095 $w=5.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.9 $Y=1.26 $X2=2.9
+ $Y2=1.075
r67 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.8 $Y=1.26
+ $X2=2.8 $Y2=1.26
r68 20 33 6.31476 $w=3.63e-07 $l=2e-07 $layer=LI1_cond $X=2.707 $Y=1.295
+ $X2=2.707 $Y2=1.495
r69 20 30 1.10508 $w=3.63e-07 $l=3.5e-08 $layer=LI1_cond $X=2.707 $Y=1.295
+ $X2=2.707 $Y2=1.26
r70 19 25 97.9104 $w=5e-07 $l=9.15e-07 $layer=POLY_cond $X=0.665 $Y=1.66
+ $X2=0.665 $Y2=0.745
r71 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.73
+ $Y=1.66 $X2=0.73 $Y2=1.66
r72 16 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.73 $Y2=1.58
r73 15 21 2.68377 $w=3.63e-07 $l=8.5e-08 $layer=LI1_cond $X=2.707 $Y=1.58
+ $X2=2.707 $Y2=1.665
r74 15 33 2.68377 $w=3.63e-07 $l=8.5e-08 $layer=LI1_cond $X=2.707 $Y=1.58
+ $X2=2.707 $Y2=1.495
r75 15 16 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=2.525 $Y=1.58
+ $X2=0.895 $Y2=1.58
r76 11 19 61.5284 $w=5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.665 $Y=2.235
+ $X2=0.665 $Y2=1.66
r77 10 12 78.325 $w=4.8e-07 $l=7.8e-07 $layer=POLY_cond $X=0.665 $Y=2.485
+ $X2=1.445 $Y2=2.485
r78 10 11 1.84115 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.665 $Y=2.485
+ $X2=0.665 $Y2=2.235
r79 9 31 31.812 $w=5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.935 $Y=0.745 $X2=2.935
+ $Y2=1.075
r80 4 12 1.84115 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.445 $Y=2.735
+ $X2=1.445 $Y2=2.485
r81 4 6 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.445 $Y=2.735 $X2=1.445
+ $Y2=3.055
r82 1 10 1.84115 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.665 $Y=2.735
+ $X2=0.665 $Y2=2.485
r83 1 3 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.665 $Y=2.735 $X2=0.665
+ $Y2=3.055
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%A_30_107# 1 2 7 9 13 16 19 23 26 30 33 34
+ 36
c73 30 0 1.43057e-19 $X=2.8 $Y=2.18
c74 26 0 6.3458e-20 $X=2.635 $Y=2.62
c75 23 0 1.88256e-19 $X=2.09 $Y=1.23
c76 7 0 1.52716e-19 $X=2.935 $Y=2.715
r77 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.8 $Y=2.18
+ $X2=2.8 $Y2=2.18
r78 28 30 16.0438 $w=2.53e-07 $l=3.55e-07 $layer=LI1_cond $X=2.762 $Y=2.535
+ $X2=2.762 $Y2=2.18
r79 27 34 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.44 $Y=2.62
+ $X2=0.275 $Y2=2.62
r80 26 28 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=2.635 $Y=2.62
+ $X2=2.762 $Y2=2.535
r81 26 27 143.203 $w=1.68e-07 $l=2.195e-06 $layer=LI1_cond $X=2.635 $Y=2.62
+ $X2=0.44 $Y2=2.62
r82 24 36 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.155 $Y=1.23
+ $X2=2.155 $Y2=0.745
r83 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.09
+ $Y=1.23 $X2=2.09 $Y2=1.23
r84 21 33 1.80668 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.44 $Y=1.205
+ $X2=0.275 $Y2=1.205
r85 21 23 86.4332 $w=2.18e-07 $l=1.65e-06 $layer=LI1_cond $X=0.44 $Y=1.205
+ $X2=2.09 $Y2=1.205
r86 17 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.275 $Y=2.705
+ $X2=0.275 $Y2=2.62
r87 17 19 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.275 $Y=2.705
+ $X2=0.275 $Y2=3.055
r88 16 34 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.195 $Y=2.535
+ $X2=0.275 $Y2=2.62
r89 15 33 4.63873 $w=2.5e-07 $l=1.44568e-07 $layer=LI1_cond $X=0.195 $Y=1.315
+ $X2=0.275 $Y2=1.205
r90 15 16 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=0.195 $Y=1.315
+ $X2=0.195 $Y2=2.535
r91 11 33 4.63873 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=0.275 $Y=1.095
+ $X2=0.275 $Y2=1.205
r92 11 13 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.275 $Y=1.095
+ $X2=0.275 $Y2=0.745
r93 7 31 47.5188 $w=5.48e-07 $l=5.52223e-07 $layer=POLY_cond $X=2.935 $Y=2.715
+ $X2=2.9 $Y2=2.18
r94 7 9 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.935 $Y=2.715 $X2=2.935
+ $Y2=3.055
r95 2 19 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.845 $X2=0.275 $Y2=3.055
r96 1 13 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.535 $X2=0.275 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%D 3 7 9 13 14
c34 7 0 4.41352e-20 $X=2.155 $Y=3.055
r35 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.11
+ $Y=1.93 $X2=2.11 $Y2=1.93
r36 9 14 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.11 $Y=2.035
+ $X2=2.11 $Y2=1.93
r37 5 13 5.92623 $w=3.66e-07 $l=4.5e-08 $layer=POLY_cond $X=2.155 $Y=1.875
+ $X2=2.11 $Y2=1.875
r38 5 7 104.866 $w=5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.155 $Y=2.075 $X2=2.155
+ $Y2=3.055
r39 1 13 87.5765 $w=3.66e-07 $l=6.65e-07 $layer=POLY_cond $X=1.445 $Y=1.875
+ $X2=2.11 $Y2=1.875
r40 1 3 99.5155 $w=5e-07 $l=9.3e-07 $layer=POLY_cond $X=1.445 $Y=1.675 $X2=1.445
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%SCD 1 2 3 8 14
c25 8 0 3.27535e-19 $X=3.645 $Y=0.745
c26 1 0 1.52716e-19 $X=3.6 $Y=1.295
r27 11 14 183.515 $w=5e-07 $l=1.715e-06 $layer=POLY_cond $X=3.645 $Y=1.34
+ $X2=3.645 $Y2=3.055
r28 8 11 63.6685 $w=5e-07 $l=5.95e-07 $layer=POLY_cond $X=3.645 $Y=0.745
+ $X2=3.645 $Y2=1.34
r29 2 3 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.585 $Y=1.665
+ $X2=3.585 $Y2=2.035
r30 1 2 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.585 $Y=1.295
+ $X2=3.585 $Y2=1.665
r31 1 11 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.585
+ $Y=1.34 $X2=3.585 $Y2=1.34
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%CLK 3 6 9 10 11 12 13 18
r39 18 20 24.2123 $w=6.15e-07 $l=2.55e-07 $layer=POLY_cond $X=4.482 $Y=1.34
+ $X2=4.482 $Y2=1.085
r40 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.36
+ $Y=1.34 $X2=4.36 $Y2=1.34
r41 12 13 7.90266 $w=5.58e-07 $l=3.7e-07 $layer=LI1_cond $X=4.245 $Y=1.665
+ $X2=4.245 $Y2=2.035
r42 12 19 6.94153 $w=5.58e-07 $l=3.25e-07 $layer=LI1_cond $X=4.245 $Y=1.665
+ $X2=4.245 $Y2=1.34
r43 11 19 0.961134 $w=5.58e-07 $l=4.5e-08 $layer=LI1_cond $X=4.245 $Y=1.295
+ $X2=4.245 $Y2=1.34
r44 9 10 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.54 $Y=3.22 $X2=4.54
+ $Y2=2.735
r45 6 10 28.7361 $w=6.15e-07 $l=3.07e-07 $layer=POLY_cond $X=4.482 $Y=2.428
+ $X2=4.482 $Y2=2.735
r46 5 18 4.52383 $w=6.15e-07 $l=5.2e-08 $layer=POLY_cond $X=4.482 $Y=1.392
+ $X2=4.482 $Y2=1.34
r47 5 6 90.1285 $w=6.15e-07 $l=1.036e-06 $layer=POLY_cond $X=4.482 $Y=1.392
+ $X2=4.482 $Y2=2.428
r48 3 20 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.425 $Y=0.745 $X2=4.425
+ $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%A_935_107# 1 2 7 9 10 12 14 16 24 28 31 33
+ 36 38 42 43 47 50 51 52 55 56 59 60 63 64 65 66 68 69 71 72 74 75 77 80 84 87
+ 88 91 93 94 103 106 110
c268 110 0 1.31759e-20 $X=7.105 $Y=0.775
c269 93 0 1.17996e-19 $X=8.272 $Y=2.66
c270 80 0 1.31874e-19 $X=13.185 $Y=1.58
c271 69 0 1.77953e-19 $X=12.042 $Y=2.935
c272 65 0 9.67046e-20 $X=9.795 $Y=3.19
c273 60 0 9.02861e-20 $X=9.625 $Y=2.66
c274 56 0 1.81757e-19 $X=8.245 $Y=2.39
c275 33 0 1.50078e-19 $X=5.505 $Y=1.82
c276 7 0 1.19183e-19 $X=6.03 $Y=2.555
r277 101 103 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=12.18 $Y=1.42
+ $X2=12.485 $Y2=1.42
r278 99 100 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.07
+ $Y=2.39 $X2=12.07 $Y2=2.39
r279 94 96 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.57 $Y=3.02
+ $X2=10.57 $Y2=3.19
r280 89 91 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.145 $Y=1.69
+ $X2=7.36 $Y2=1.69
r281 84 86 10.5766 $w=3.63e-07 $l=2.3e-07 $layer=LI1_cond $X=4.832 $Y=0.745
+ $X2=4.832 $Y2=0.975
r282 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.185
+ $Y=1.58 $X2=13.185 $Y2=1.58
r283 78 80 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=13.225 $Y=0.785
+ $X2=13.225 $Y2=1.58
r284 76 103 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.485 $Y=1.505
+ $X2=12.485 $Y2=1.42
r285 76 77 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=12.485 $Y=1.505
+ $X2=12.485 $Y2=2.225
r286 74 78 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=13.1 $Y=0.7
+ $X2=13.225 $Y2=0.785
r287 74 75 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=13.1 $Y=0.7
+ $X2=12.265 $Y2=0.7
r288 73 99 4.53113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=12.18 $Y=2.31
+ $X2=12.042 $Y2=2.31
r289 72 77 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.4 $Y=2.31
+ $X2=12.485 $Y2=2.225
r290 72 73 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=12.4 $Y=2.31
+ $X2=12.18 $Y2=2.31
r291 71 101 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.18 $Y=1.335
+ $X2=12.18 $Y2=1.42
r292 70 75 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.18 $Y=0.785
+ $X2=12.265 $Y2=0.7
r293 70 71 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=12.18 $Y=0.785
+ $X2=12.18 $Y2=1.335
r294 68 99 2.79091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=12.042 $Y=2.395
+ $X2=12.042 $Y2=2.31
r295 68 69 22.6298 $w=2.73e-07 $l=5.4e-07 $layer=LI1_cond $X=12.042 $Y=2.395
+ $X2=12.042 $Y2=2.935
r296 67 94 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.655 $Y=3.02
+ $X2=10.57 $Y2=3.02
r297 66 69 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=11.905 $Y=3.02
+ $X2=12.042 $Y2=2.935
r298 66 67 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=11.905 $Y=3.02
+ $X2=10.655 $Y2=3.02
r299 64 96 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.485 $Y=3.19
+ $X2=10.57 $Y2=3.19
r300 64 65 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.485 $Y=3.19
+ $X2=9.795 $Y2=3.19
r301 63 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.71 $Y=3.105
+ $X2=9.795 $Y2=3.19
r302 62 63 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.71 $Y=2.745
+ $X2=9.71 $Y2=3.105
r303 61 93 2.32734 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=8.41 $Y=2.66
+ $X2=8.272 $Y2=2.66
r304 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.625 $Y=2.66
+ $X2=9.71 $Y2=2.745
r305 60 61 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=9.625 $Y=2.66
+ $X2=8.41 $Y2=2.66
r306 58 93 4.10697 $w=2.22e-07 $l=1.07912e-07 $layer=LI1_cond $X=8.22 $Y=2.745
+ $X2=8.272 $Y2=2.66
r307 58 59 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=8.22 $Y=2.745
+ $X2=8.22 $Y2=3.355
r308 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.245
+ $Y=2.39 $X2=8.245 $Y2=2.39
r309 53 93 4.10697 $w=2.22e-07 $l=8.5e-08 $layer=LI1_cond $X=8.272 $Y=2.575
+ $X2=8.272 $Y2=2.66
r310 53 55 7.7528 $w=2.73e-07 $l=1.85e-07 $layer=LI1_cond $X=8.272 $Y=2.575
+ $X2=8.272 $Y2=2.39
r311 51 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.135 $Y=3.44
+ $X2=8.22 $Y2=3.355
r312 51 52 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.135 $Y=3.44
+ $X2=7.445 $Y2=3.44
r313 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.36 $Y=3.355
+ $X2=7.445 $Y2=3.44
r314 49 91 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=1.775
+ $X2=7.36 $Y2=1.69
r315 49 50 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=7.36 $Y=1.775
+ $X2=7.36 $Y2=3.355
r316 48 110 52.9679 $w=5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.105 $Y=1.27
+ $X2=7.105 $Y2=0.775
r317 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.145
+ $Y=1.27 $X2=7.145 $Y2=1.27
r318 45 89 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.145 $Y=1.605
+ $X2=7.145 $Y2=1.69
r319 45 47 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.145 $Y=1.605
+ $X2=7.145 $Y2=1.27
r320 44 47 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=7.145 $Y=0.435
+ $X2=7.145 $Y2=1.27
r321 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.06 $Y=0.35
+ $X2=7.145 $Y2=0.435
r322 42 43 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=7.06 $Y=0.35
+ $X2=5.8 $Y2=0.35
r323 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.715 $Y=0.435
+ $X2=5.8 $Y2=0.35
r324 40 88 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=5.715 $Y=0.435
+ $X2=5.715 $Y2=1.235
r325 39 106 61.5284 $w=5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.755 $Y=1.4
+ $X2=5.755 $Y2=0.825
r326 38 88 7.64045 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.67 $Y=1.4
+ $X2=5.67 $Y2=1.235
r327 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.67
+ $Y=1.4 $X2=5.67 $Y2=1.4
r328 36 38 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.67 $Y=1.735
+ $X2=5.67 $Y2=1.4
r329 34 87 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.015 $Y=1.82
+ $X2=4.93 $Y2=1.82
r330 33 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.505 $Y=1.82
+ $X2=5.67 $Y2=1.735
r331 33 34 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=5.505 $Y=1.82
+ $X2=5.015 $Y2=1.82
r332 29 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=1.905
+ $X2=4.93 $Y2=1.82
r333 29 31 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=4.93 $Y=1.905
+ $X2=4.93 $Y2=3.13
r334 28 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=1.735
+ $X2=4.93 $Y2=1.82
r335 28 86 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.93 $Y=1.735
+ $X2=4.93 $Y2=0.975
r336 25 56 32.1495 $w=3.5e-07 $l=1.95e-07 $layer=POLY_cond $X=8.255 $Y=2.585
+ $X2=8.255 $Y2=2.39
r337 24 25 41.2577 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=8.18 $Y=2.925
+ $X2=8.18 $Y2=2.585
r338 18 39 105.401 $w=5e-07 $l=9.85e-07 $layer=POLY_cond $X=5.755 $Y=2.385
+ $X2=5.755 $Y2=1.4
r339 14 81 19.4359 $w=5e-07 $l=1.85997e-07 $layer=POLY_cond $X=13.095 $Y=1.395
+ $X2=13.097 $Y2=1.58
r340 14 16 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=13.095 $Y=1.395
+ $X2=13.095 $Y2=1.075
r341 10 100 17.1785 $w=5e-07 $l=1.75e-07 $layer=POLY_cond $X=12.135 $Y=2.565
+ $X2=12.135 $Y2=2.39
r342 10 12 69.5538 $w=5e-07 $l=6.5e-07 $layer=POLY_cond $X=12.135 $Y=2.565
+ $X2=12.135 $Y2=3.215
r343 7 18 116.272 $w=1.7e-07 $l=2.75e-07 $layer=POLY_cond $X=6.03 $Y=2.47
+ $X2=5.755 $Y2=2.47
r344 7 9 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.03 $Y=2.555 $X2=6.03
+ $Y2=3.04
r345 2 31 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=4.79
+ $Y=2.845 $X2=4.93 $Y2=3.13
r346 1 84 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.675
+ $Y=0.535 $X2=4.815 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%A_1201_123# 1 2 9 13 17 19 21 25 28 30 33
+ 37 38 39 40 42 48 49 58
c159 58 0 2.04378e-19 $X=7.885 $Y=1.985
c160 49 0 1.31874e-19 $X=12.135 $Y=1.85
c161 48 0 1.61924e-19 $X=12.135 $Y=1.85
c162 39 0 1.31759e-20 $X=6.335 $Y=1.425
c163 38 0 1.50078e-19 $X=6.4 $Y=1.59
c164 25 0 1.02273e-19 $X=6.335 $Y=1.9
c165 19 0 1.77953e-19 $X=13.03 $Y=2.605
c166 17 0 1.43632e-19 $X=12.22 $Y=0.91
r167 57 58 35.2594 $w=6.63e-07 $l=4.85e-07 $layer=POLY_cond $X=7.4 $Y=1.985
+ $X2=7.885 $Y2=1.985
r168 53 57 70.5189 $w=6.63e-07 $l=9.7e-07 $layer=POLY_cond $X=6.43 $Y=1.985
+ $X2=7.4 $Y2=1.985
r169 48 51 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=12.095 $Y=1.85
+ $X2=12.095 $Y2=1.96
r170 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.135
+ $Y=1.85 $X2=12.135 $Y2=1.85
r171 43 58 18.5385 $w=6.63e-07 $l=2.55e-07 $layer=POLY_cond $X=8.14 $Y=1.985
+ $X2=7.885 $Y2=1.985
r172 42 45 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=8.14 $Y=1.815
+ $X2=8.14 $Y2=1.96
r173 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.14
+ $Y=1.815 $X2=8.14 $Y2=1.815
r174 38 53 51.0886 $w=4.3e-07 $l=3.95e-07 $layer=POLY_cond $X=6.43 $Y=1.59
+ $X2=6.43 $Y2=1.985
r175 37 39 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=6.335 $Y=1.59
+ $X2=6.335 $Y2=1.425
r176 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.4
+ $Y=1.59 $X2=6.4 $Y2=1.59
r177 35 39 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.225 $Y=1.055
+ $X2=6.225 $Y2=1.425
r178 33 35 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=6.145 $Y=0.825
+ $X2=6.145 $Y2=1.055
r179 31 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.305 $Y=1.96
+ $X2=8.14 $Y2=1.96
r180 30 51 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.97 $Y=1.96
+ $X2=12.095 $Y2=1.96
r181 30 31 239.107 $w=1.68e-07 $l=3.665e-06 $layer=LI1_cond $X=11.97 $Y=1.96
+ $X2=8.305 $Y2=1.96
r182 28 40 29.1254 $w=2.73e-07 $l=6.95e-07 $layer=LI1_cond $X=6.392 $Y=2.79
+ $X2=6.392 $Y2=2.095
r183 25 40 6.77877 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=6.335 $Y=1.9
+ $X2=6.335 $Y2=2.095
r184 24 37 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=6.335 $Y=1.62
+ $X2=6.335 $Y2=1.59
r185 24 25 8.27395 $w=3.88e-07 $l=2.8e-07 $layer=LI1_cond $X=6.335 $Y=1.62
+ $X2=6.335 $Y2=1.9
r186 19 49 104.706 $w=4.12e-07 $l=1.05856e-06 $layer=POLY_cond $X=13.03 $Y=2.207
+ $X2=12.135 $Y2=1.85
r187 19 21 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=13.03 $Y=2.605
+ $X2=13.03 $Y2=2.925
r188 17 49 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=12.22 $Y=0.91 $X2=12.22
+ $Y2=1.81
r189 11 58 9.44957 $w=5e-07 $l=8.7e-07 $layer=POLY_cond $X=7.885 $Y=1.115
+ $X2=7.885 $Y2=1.985
r190 11 13 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.885 $Y=1.115
+ $X2=7.885 $Y2=0.775
r191 7 57 9.44957 $w=5e-07 $l=6e-07 $layer=POLY_cond $X=7.4 $Y=2.585 $X2=7.4
+ $Y2=1.985
r192 7 9 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.4 $Y=2.585 $X2=7.4
+ $Y2=2.925
r193 2 28 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=6.28
+ $Y=2.665 $X2=6.42 $Y2=2.79
r194 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.005
+ $Y=0.615 $X2=6.145 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%A_1669_87# 1 2 7 9 10 13 15 19 23 29 30 33
c61 13 0 1.48209e-19 $X=8.955 $Y=2.31
r62 27 30 12.105 $w=4.38e-07 $l=1.1e-07 $layer=POLY_cond $X=9 $Y=1.345 $X2=8.89
+ $Y2=1.345
r63 26 29 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=9 $Y=1.225
+ $X2=9.165 $Y2=1.225
r64 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9 $Y=1.26
+ $X2=9 $Y2=1.26
r65 21 23 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=10.14 $Y=2.395
+ $X2=10.14 $Y2=2.84
r66 17 19 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=9.535 $Y=1.105
+ $X2=9.535 $Y2=0.745
r67 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.37 $Y=1.19
+ $X2=9.535 $Y2=1.105
r68 15 29 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=9.37 $Y=1.19
+ $X2=9.165 $Y2=1.19
r69 13 33 65.8086 $w=5e-07 $l=6.15e-07 $layer=POLY_cond $X=8.89 $Y=2.31 $X2=8.89
+ $Y2=2.925
r70 13 30 76.5092 $w=5e-07 $l=7.15e-07 $layer=POLY_cond $X=8.89 $Y=2.31 $X2=8.89
+ $Y2=1.595
r71 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.955
+ $Y=2.31 $X2=8.955 $Y2=2.31
r72 10 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.975 $Y=2.31
+ $X2=10.14 $Y2=2.395
r73 10 12 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=9.975 $Y=2.31
+ $X2=8.955 $Y2=2.31
r74 7 30 32.4635 $w=4.38e-07 $l=2.95e-07 $layer=POLY_cond $X=8.595 $Y=1.345
+ $X2=8.89 $Y2=1.345
r75 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.595 $Y=1.095 $X2=8.595
+ $Y2=0.775
r76 2 23 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=10
+ $Y=2.715 $X2=10.14 $Y2=2.84
r77 1 19 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.41
+ $Y=0.535 $X2=9.535 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%A_1471_113# 1 2 9 12 16 19 20 22 25 27 29
+ 35 36 41 43 44 45 51 52 53 56
c137 29 0 1.81757e-19 $X=8.485 $Y=1.44
c138 25 0 5.1504e-20 $X=7.79 $Y=2.84
c139 12 0 1.61924e-19 $X=11.425 $Y=3.215
r140 51 56 144.458 $w=5e-07 $l=1.35e-06 $layer=POLY_cond $X=9.75 $Y=1.575
+ $X2=9.75 $Y2=2.925
r141 50 53 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=9.685 $Y=1.575
+ $X2=9.85 $Y2=1.575
r142 50 52 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=9.685 $Y=1.575
+ $X2=9.52 $Y2=1.575
r143 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.685
+ $Y=1.575 $X2=9.685 $Y2=1.575
r144 45 47 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.57 $Y=1.44
+ $X2=8.57 $Y2=1.61
r145 39 41 5.14314 $w=4.98e-07 $l=2.15e-07 $layer=LI1_cond $X=7.495 $Y=0.775
+ $X2=7.71 $Y2=0.775
r146 36 60 29.1757 $w=5.85e-07 $l=3.05e-07 $layer=POLY_cond $X=11.467 $Y=1.61
+ $X2=11.467 $Y2=1.915
r147 36 59 19.1153 $w=5.85e-07 $l=1.95e-07 $layer=POLY_cond $X=11.467 $Y=1.61
+ $X2=11.467 $Y2=1.415
r148 35 53 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=11.36 $Y=1.61
+ $X2=9.85 $Y2=1.61
r149 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.36
+ $Y=1.61 $X2=11.36 $Y2=1.61
r150 32 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.655 $Y=1.61
+ $X2=8.57 $Y2=1.61
r151 32 52 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=8.655 $Y=1.61
+ $X2=9.52 $Y2=1.61
r152 30 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.795 $Y=1.44
+ $X2=7.71 $Y2=1.44
r153 29 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.485 $Y=1.44
+ $X2=8.57 $Y2=1.44
r154 29 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.485 $Y=1.44
+ $X2=7.795 $Y2=1.44
r155 25 44 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.79 $Y=2.84
+ $X2=7.79 $Y2=2.675
r156 25 27 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.79 $Y=2.84
+ $X2=7.79 $Y2=2.925
r157 23 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.71 $Y=1.525
+ $X2=7.71 $Y2=1.44
r158 23 44 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=7.71 $Y=1.525
+ $X2=7.71 $Y2=2.675
r159 22 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.71 $Y=1.355
+ $X2=7.71 $Y2=1.44
r160 21 41 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=7.71 $Y=1.025
+ $X2=7.71 $Y2=0.775
r161 21 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.71 $Y=1.025
+ $X2=7.71 $Y2=1.355
r162 20 51 1.07006 $w=5e-07 $l=1e-08 $layer=POLY_cond $X=9.75 $Y=1.565 $X2=9.75
+ $Y2=1.575
r163 19 20 39.6318 $w=6.75e-07 $l=5e-07 $layer=POLY_cond $X=9.837 $Y=1.065
+ $X2=9.837 $Y2=1.565
r164 16 59 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=11.51 $Y=0.91
+ $X2=11.51 $Y2=1.415
r165 12 60 139.108 $w=5e-07 $l=1.3e-06 $layer=POLY_cond $X=11.425 $Y=3.215
+ $X2=11.425 $Y2=1.915
r166 9 19 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.925 $Y=0.745
+ $X2=9.925 $Y2=1.065
r167 2 27 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.65
+ $Y=2.715 $X2=7.79 $Y2=2.925
r168 1 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.355
+ $Y=0.565 $X2=7.495 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%SET_B 3 6 7 13 14 15 18 19 20 25 29 35 45
c88 6 0 9.02861e-20 $X=10.582 $Y=2.605
r89 32 35 143.923 $w=5e-07 $l=1.345e-06 $layer=POLY_cond $X=14.52 $Y=1.58
+ $X2=14.52 $Y2=2.925
r90 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.435
+ $Y=1.58 $X2=14.435 $Y2=1.58
r91 29 32 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=14.52 $Y=1.075
+ $X2=14.52 $Y2=1.58
r92 20 33 2.14035 $w=4.73e-07 $l=8.5e-08 $layer=LI1_cond $X=14.282 $Y=1.665
+ $X2=14.282 $Y2=1.58
r93 19 33 7.17647 $w=4.73e-07 $l=2.85e-07 $layer=LI1_cond $X=14.282 $Y=1.295
+ $X2=14.282 $Y2=1.58
r94 19 37 6.24479 $w=4.73e-07 $l=2.48e-07 $layer=LI1_cond $X=14.282 $Y=1.295
+ $X2=14.282 $Y2=1.047
r95 18 37 3.07203 $w=4.73e-07 $l=1.22e-07 $layer=LI1_cond $X=14.282 $Y=0.925
+ $X2=14.282 $Y2=1.047
r96 18 45 8.10777 $w=4.73e-07 $l=1.15e-07 $layer=LI1_cond $X=14.282 $Y=0.925
+ $X2=14.282 $Y2=0.81
r97 16 45 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=14.13 $Y=0.435
+ $X2=14.13 $Y2=0.81
r98 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.045 $Y=0.35
+ $X2=14.13 $Y2=0.435
r99 14 15 157.23 $w=1.68e-07 $l=2.41e-06 $layer=LI1_cond $X=14.045 $Y=0.35
+ $X2=11.635 $Y2=0.35
r100 12 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.55 $Y=0.435
+ $X2=11.635 $Y2=0.35
r101 12 13 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=11.55 $Y=0.435
+ $X2=11.55 $Y2=1.175
r102 10 25 55.108 $w=5e-07 $l=5.15e-07 $layer=POLY_cond $X=10.635 $Y=1.26
+ $X2=10.635 $Y2=0.745
r103 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.7
+ $Y=1.26 $X2=10.7 $Y2=1.26
r104 7 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.465 $Y=1.26
+ $X2=11.55 $Y2=1.175
r105 7 9 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=11.465 $Y=1.26
+ $X2=10.7 $Y2=1.26
r106 5 10 90.42 $w=5e-07 $l=8.45e-07 $layer=POLY_cond $X=10.635 $Y=2.105
+ $X2=10.635 $Y2=1.26
r107 5 6 44.2173 $w=6.05e-07 $l=5e-07 $layer=POLY_cond $X=10.582 $Y=2.105
+ $X2=10.582 $Y2=2.605
r108 3 6 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.53 $Y=2.925 $X2=10.53
+ $Y2=2.605
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%A_2698_421# 1 2 9 12 14 17 20 21 22 26 27
+ 29 37
c72 37 0 9.75335e-20 $X=13.775 $Y=2.605
c73 17 0 1.96117e-19 $X=13.875 $Y=2.39
r74 27 29 74.6783 $w=2.48e-07 $l=1.62e-06 $layer=LI1_cond $X=15.895 $Y=2.695
+ $X2=15.895 $Y2=1.075
r75 24 26 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=15.46 $Y=3.335
+ $X2=15.46 $Y2=3.275
r76 23 27 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=15.46 $Y=2.78
+ $X2=15.895 $Y2=2.78
r77 23 26 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=15.46 $Y=2.865
+ $X2=15.46 $Y2=3.275
r78 21 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=15.295 $Y=3.42
+ $X2=15.46 $Y2=3.335
r79 21 22 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=15.295 $Y=3.42
+ $X2=14.565 $Y2=3.42
r80 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.48 $Y=3.335
+ $X2=14.565 $Y2=3.42
r81 19 20 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=14.48 $Y=2.495
+ $X2=14.48 $Y2=3.335
r82 17 37 21.1255 $w=5.7e-07 $l=2.15e-07 $layer=POLY_cond $X=13.775 $Y=2.39
+ $X2=13.775 $Y2=2.605
r83 17 36 27.696 $w=5.7e-07 $l=2.85e-07 $layer=POLY_cond $X=13.775 $Y=2.39
+ $X2=13.775 $Y2=2.105
r84 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.875
+ $Y=2.39 $X2=13.875 $Y2=2.39
r85 14 19 6.89401 $w=2.05e-07 $l=1.39155e-07 $layer=LI1_cond $X=14.395 $Y=2.392
+ $X2=14.48 $Y2=2.495
r86 14 16 28.133 $w=2.03e-07 $l=5.2e-07 $layer=LI1_cond $X=14.395 $Y=2.392
+ $X2=13.875 $Y2=2.392
r87 12 36 110.216 $w=5e-07 $l=1.03e-06 $layer=POLY_cond $X=13.81 $Y=1.075
+ $X2=13.81 $Y2=2.105
r88 9 37 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=13.74 $Y=2.925 $X2=13.74
+ $Y2=2.605
r89 2 26 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=15.335
+ $Y=3.065 $X2=15.46 $Y2=3.275
r90 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=15.715
+ $Y=0.865 $X2=15.855 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%A_2477_543# 1 2 3 12 16 18 22 26 28 31 33
+ 38 40 45 47 49 55 57 59 66
c124 55 0 9.75335e-20 $X=12.835 $Y=2.76
c125 47 0 1.96117e-19 $X=15.42 $Y=1.94
r126 65 66 23.0853 $w=7.8e-07 $l=2.5e-07 $layer=POLY_cond $X=15.85 $Y=1.805
+ $X2=16.1 $Y2=1.805
r127 64 65 25.379 $w=7.8e-07 $l=3.85e-07 $layer=POLY_cond $X=15.465 $Y=1.805
+ $X2=15.85 $Y2=1.805
r128 53 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=12.525 $Y=2.76
+ $X2=12.835 $Y2=2.76
r129 50 64 2.96637 $w=7.8e-07 $l=4.5e-08 $layer=POLY_cond $X=15.42 $Y=1.805
+ $X2=15.465 $Y2=1.805
r130 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=15.42
+ $Y=1.67 $X2=15.42 $Y2=1.67
r131 47 49 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=15.42 $Y=1.94
+ $X2=15.42 $Y2=1.67
r132 43 47 25.0105 $w=2.33e-07 $l=5.1e-07 $layer=LI1_cond $X=14.91 $Y=2.057
+ $X2=15.42 $Y2=2.057
r133 43 59 8.99284 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=14.91 $Y=2.057
+ $X2=14.745 $Y2=2.057
r134 43 45 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=14.91 $Y=2.175
+ $X2=14.91 $Y2=2.925
r135 42 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.92 $Y=2.025
+ $X2=12.835 $Y2=2.025
r136 42 59 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=12.92 $Y=2.025
+ $X2=14.745 $Y2=2.025
r137 40 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.835 $Y=2.675
+ $X2=12.835 $Y2=2.76
r138 39 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.835 $Y=2.11
+ $X2=12.835 $Y2=2.025
r139 39 40 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=12.835 $Y=2.11
+ $X2=12.835 $Y2=2.675
r140 38 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.835 $Y=1.94
+ $X2=12.835 $Y2=2.025
r141 37 38 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=12.835 $Y=1.155
+ $X2=12.835 $Y2=1.94
r142 33 37 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=12.75 $Y=1.06
+ $X2=12.835 $Y2=1.155
r143 33 35 8.17225 $w=1.88e-07 $l=1.4e-07 $layer=LI1_cond $X=12.75 $Y=1.06
+ $X2=12.61 $Y2=1.06
r144 31 53 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.525 $Y=3.215
+ $X2=12.525 $Y2=2.845
r145 24 28 20.4101 $w=5e-07 $l=2.59808e-07 $layer=POLY_cond $X=17.18 $Y=1.915
+ $X2=17.16 $Y2=1.665
r146 24 26 89.3499 $w=5e-07 $l=8.35e-07 $layer=POLY_cond $X=17.18 $Y=1.915
+ $X2=17.18 $Y2=2.75
r147 20 28 20.4101 $w=5e-07 $l=2.59808e-07 $layer=POLY_cond $X=17.14 $Y=1.415
+ $X2=17.16 $Y2=1.665
r148 20 22 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=17.14 $Y=1.415
+ $X2=17.14 $Y2=1.075
r149 18 28 5.30422 $w=5e-07 $l=2.7e-07 $layer=POLY_cond $X=16.89 $Y=1.665
+ $X2=17.16 $Y2=1.665
r150 18 66 84.5347 $w=5e-07 $l=7.9e-07 $layer=POLY_cond $X=16.89 $Y=1.665
+ $X2=16.1 $Y2=1.665
r151 14 65 13.1928 $w=5e-07 $l=3.9e-07 $layer=POLY_cond $X=15.85 $Y=2.195
+ $X2=15.85 $Y2=1.805
r152 14 16 115.566 $w=5e-07 $l=1.08e-06 $layer=POLY_cond $X=15.85 $Y=2.195
+ $X2=15.85 $Y2=3.275
r153 10 64 13.1928 $w=5e-07 $l=3.9e-07 $layer=POLY_cond $X=15.465 $Y=1.415
+ $X2=15.465 $Y2=1.805
r154 10 12 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=15.465 $Y=1.415
+ $X2=15.465 $Y2=1.075
r155 3 45 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=14.77
+ $Y=2.715 $X2=14.91 $Y2=2.925
r156 2 53 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=12.385
+ $Y=2.715 $X2=12.525 $Y2=2.84
r157 2 31 300 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_PDIFF $count=2 $X=12.385
+ $Y=2.715 $X2=12.525 $Y2=3.215
r158 1 35 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=12.47
+ $Y=0.535 $X2=12.61 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%A_3321_173# 1 2 9 13 17 23 27 29 30 32 33
r49 33 36 54.5563 $w=5.75e-07 $l=5.75e-07 $layer=POLY_cond $X=18.017 $Y=1.67
+ $X2=18.017 $Y2=2.245
r50 33 35 24.7808 $w=5.75e-07 $l=2.55e-07 $layer=POLY_cond $X=18.017 $Y=1.67
+ $X2=18.017 $Y2=1.415
r51 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=17.915
+ $Y=1.67 $X2=17.915 $Y2=1.67
r52 29 30 5.30085 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=16.77 $Y=2.52
+ $X2=16.77 $Y2=2.355
r53 24 27 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.915 $Y=1.59
+ $X2=16.75 $Y2=1.59
r54 23 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.75 $Y=1.59
+ $X2=17.915 $Y2=1.59
r55 23 24 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=17.75 $Y=1.59
+ $X2=16.915 $Y2=1.59
r56 19 27 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=16.75 $Y=1.675
+ $X2=16.75 $Y2=1.59
r57 19 30 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=16.75 $Y=1.675
+ $X2=16.75 $Y2=2.355
r58 15 27 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=16.75 $Y=1.505
+ $X2=16.75 $Y2=1.59
r59 15 17 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=16.75 $Y=1.505
+ $X2=16.75 $Y2=1.075
r60 13 36 67.4137 $w=5e-07 $l=6.3e-07 $layer=POLY_cond $X=18.055 $Y=2.875
+ $X2=18.055 $Y2=2.245
r61 9 35 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=18.035 $Y=0.91
+ $X2=18.035 $Y2=1.415
r62 2 29 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=16.665
+ $Y=2.375 $X2=16.79 $Y2=2.52
r63 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=16.605
+ $Y=0.865 $X2=16.75 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%VPWR 1 2 3 4 5 6 7 8 25 28 37 48 55 69 73
+ 82 89 97
r131 95 97 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=17.245 $Y=3.63
+ $X2=17.965 $Y2=3.63
r132 94 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.965 $Y=3.59
+ $X2=17.965 $Y2=3.59
r133 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.245 $Y=3.59
+ $X2=17.245 $Y2=3.59
r134 92 94 4.64762 $w=9.43e-07 $l=3.6e-07 $layer=LI1_cond $X=17.607 $Y=3.23
+ $X2=17.607 $Y2=3.59
r135 89 92 9.16614 $w=9.43e-07 $l=7.1e-07 $layer=LI1_cond $X=17.607 $Y=2.52
+ $X2=17.607 $Y2=3.23
r136 86 95 0.36663 $w=3.7e-07 $l=9.55e-07 $layer=MET1_cond $X=16.29 $Y=3.63
+ $X2=17.245 $Y2=3.63
r137 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.29 $Y=3.59
+ $X2=16.29 $Y2=3.59
r138 82 85 6.38584 $w=5.88e-07 $l=3.15e-07 $layer=LI1_cond $X=16.11 $Y=3.275
+ $X2=16.11 $Y2=3.59
r139 79 86 0.840753 $w=3.7e-07 $l=2.19e-06 $layer=MET1_cond $X=14.1 $Y=3.63
+ $X2=16.29 $Y2=3.63
r140 77 79 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=13.38 $Y=3.63
+ $X2=14.1 $Y2=3.63
r141 76 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.1 $Y=3.59
+ $X2=14.1 $Y2=3.59
r142 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.38 $Y=3.59
+ $X2=13.38 $Y2=3.59
r143 73 76 8.54 $w=9.48e-07 $l=6.65e-07 $layer=LI1_cond $X=13.74 $Y=2.925
+ $X2=13.74 $Y2=3.59
r144 70 77 0.656478 $w=3.7e-07 $l=1.71e-06 $layer=MET1_cond $X=11.67 $Y=3.63
+ $X2=13.38 $Y2=3.63
r145 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.67 $Y=3.59
+ $X2=11.67 $Y2=3.59
r146 65 70 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.95 $Y=3.63
+ $X2=11.67 $Y2=3.63
r147 64 69 18.3229 $w=4.68e-07 $l=7.2e-07 $layer=LI1_cond $X=10.95 $Y=3.52
+ $X2=11.67 $Y2=3.52
r148 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.95 $Y=3.59
+ $X2=10.95 $Y2=3.59
r149 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.61 $Y=3.59
+ $X2=8.61 $Y2=3.59
r150 55 58 7.44842 $w=9.48e-07 $l=5.8e-07 $layer=LI1_cond $X=8.97 $Y=3.01
+ $X2=8.97 $Y2=3.59
r151 52 59 1.14212 $w=3.7e-07 $l=2.975e-06 $layer=MET1_cond $X=5.635 $Y=3.63
+ $X2=8.61 $Y2=3.63
r152 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.635 $Y=3.59
+ $X2=5.635 $Y2=3.59
r153 48 51 49.2929 $w=1.78e-07 $l=8e-07 $layer=LI1_cond $X=5.635 $Y=2.79
+ $X2=5.635 $Y2=3.59
r154 45 52 0.541307 $w=3.7e-07 $l=1.41e-06 $layer=MET1_cond $X=4.225 $Y=3.63
+ $X2=5.635 $Y2=3.63
r155 43 45 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.505 $Y=3.63
+ $X2=4.225 $Y2=3.63
r156 42 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.225 $Y=3.59
+ $X2=4.225 $Y2=3.59
r157 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.505 $Y=3.59
+ $X2=3.505 $Y2=3.59
r158 40 42 1.63575 $w=8.93e-07 $l=1.2e-07 $layer=LI1_cond $X=3.867 $Y=3.47
+ $X2=3.867 $Y2=3.59
r159 37 40 6.81564 $w=8.93e-07 $l=5e-07 $layer=LI1_cond $X=3.867 $Y=2.97
+ $X2=3.867 $Y2=3.47
r160 34 43 0.787006 $w=3.7e-07 $l=2.05e-06 $layer=MET1_cond $X=1.455 $Y=3.63
+ $X2=3.505 $Y2=3.63
r161 32 34 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.735 $Y=3.63
+ $X2=1.455 $Y2=3.63
r162 31 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.455 $Y=3.59
+ $X2=1.455 $Y2=3.59
r163 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.735 $Y=3.59
+ $X2=0.735 $Y2=3.59
r164 28 31 6.87053 $w=9.48e-07 $l=5.35e-07 $layer=LI1_cond $X=1.095 $Y=3.055
+ $X2=1.095 $Y2=3.59
r165 25 65 0.621927 $w=3.7e-07 $l=1.62e-06 $layer=MET1_cond $X=9.33 $Y=3.63
+ $X2=10.95 $Y2=3.63
r166 25 59 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=9.33 $Y=3.63
+ $X2=8.61 $Y2=3.63
r167 25 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.33 $Y=3.59
+ $X2=9.33 $Y2=3.59
r168 8 92 600 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=17.43
+ $Y=2.375 $X2=17.665 $Y2=3.23
r169 8 89 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=17.43
+ $Y=2.375 $X2=17.665 $Y2=2.52
r170 7 82 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=16.1
+ $Y=3.065 $X2=16.24 $Y2=3.275
r171 6 73 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=13.99
+ $Y=2.715 $X2=14.13 $Y2=2.925
r172 5 64 600 $w=1.7e-07 $l=8.83346e-07 $layer=licon1_PDIFF $count=1 $X=10.78
+ $Y=2.715 $X2=11.035 $Y2=3.48
r173 4 55 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=9.14
+ $Y=2.715 $X2=9.28 $Y2=3.01
r174 3 48 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=5.495
+ $Y=2.665 $X2=5.64 $Y2=2.79
r175 2 40 600 $w=1.7e-07 $l=7.4162e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=2.845 $X2=4.15 $Y2=3.47
r176 2 37 600 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=2.845 $X2=4.15 $Y2=2.97
r177 1 28 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.915
+ $Y=2.845 $X2=1.055 $Y2=3.055
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%A_481_107# 1 2 3 4 13 15 18 20 21 24 25 26
+ 28 29 30 32 33 34 37 40 42 46 51 53 56
c133 56 0 1.19183e-19 $X=6.902 $Y=2.675
c134 51 0 4.41352e-20 $X=3.155 $Y=2.54
c135 32 0 8.63818e-20 $X=5.99 $Y=3.635
r136 55 56 107.647 $w=1.68e-07 $l=1.65e-06 $layer=LI1_cond $X=6.795 $Y=1.025
+ $X2=6.795 $Y2=2.675
r137 53 55 11.256 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6.715 $Y=0.78
+ $X2=6.715 $Y2=1.025
r138 46 49 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=2.97
+ $X2=2.545 $Y2=3.055
r139 42 44 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=0.745
+ $X2=2.545 $Y2=0.83
r140 38 40 21.2528 $w=3.83e-07 $l=7.1e-07 $layer=LI1_cond $X=6.902 $Y=3.635
+ $X2=6.902 $Y2=2.925
r141 37 56 9.39714 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=6.902 $Y=2.867
+ $X2=6.902 $Y2=2.675
r142 37 40 1.73615 $w=3.83e-07 $l=5.8e-08 $layer=LI1_cond $X=6.902 $Y=2.867
+ $X2=6.902 $Y2=2.925
r143 33 38 8.24022 $w=1.7e-07 $l=2.30617e-07 $layer=LI1_cond $X=6.71 $Y=3.72
+ $X2=6.902 $Y2=3.635
r144 33 34 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.71 $Y=3.72
+ $X2=6.075 $Y2=3.72
r145 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.99 $Y=3.635
+ $X2=6.075 $Y2=3.72
r146 31 32 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=5.99 $Y=2.445
+ $X2=5.99 $Y2=3.635
r147 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.905 $Y=2.36
+ $X2=5.99 $Y2=2.445
r148 29 30 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.905 $Y=2.36
+ $X2=5.365 $Y2=2.36
r149 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.28 $Y=2.445
+ $X2=5.365 $Y2=2.36
r150 27 28 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=5.28 $Y=2.445
+ $X2=5.28 $Y2=3.635
r151 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.195 $Y=3.72
+ $X2=5.28 $Y2=3.635
r152 25 26 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.195 $Y=3.72
+ $X2=4.665 $Y2=3.72
r153 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.58 $Y=3.635
+ $X2=4.665 $Y2=3.72
r154 23 24 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=4.58 $Y=2.625
+ $X2=4.58 $Y2=3.635
r155 22 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.24 $Y=2.54
+ $X2=3.155 $Y2=2.54
r156 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.495 $Y=2.54
+ $X2=4.58 $Y2=2.625
r157 21 22 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=4.495 $Y=2.54
+ $X2=3.24 $Y2=2.54
r158 19 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=2.625
+ $X2=3.155 $Y2=2.54
r159 19 20 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.155 $Y=2.625
+ $X2=3.155 $Y2=2.885
r160 18 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=2.455
+ $X2=3.155 $Y2=2.54
r161 17 18 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=3.155 $Y=0.915
+ $X2=3.155 $Y2=2.455
r162 16 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=2.97
+ $X2=2.545 $Y2=2.97
r163 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.07 $Y=2.97
+ $X2=3.155 $Y2=2.885
r164 15 16 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.07 $Y=2.97
+ $X2=2.71 $Y2=2.97
r165 14 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0.83
+ $X2=2.545 $Y2=0.83
r166 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.07 $Y=0.83
+ $X2=3.155 $Y2=0.915
r167 13 14 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.07 $Y=0.83
+ $X2=2.71 $Y2=0.83
r168 4 40 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=6.865
+ $Y=2.715 $X2=7.01 $Y2=2.925
r169 3 49 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=2.845 $X2=2.545 $Y2=3.055
r170 2 53 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=6.57
+ $Y=0.565 $X2=6.715 $Y2=0.78
r171 1 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.405
+ $Y=0.535 $X2=2.545 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%Q 1 2 7 8 9 10 11 12 13 22
r12 12 13 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=18.435 $Y=2.775
+ $X2=18.435 $Y2=3.145
r13 12 35 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=18.435 $Y=2.775
+ $X2=18.435 $Y2=2.52
r14 11 35 3.7866 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=18.435 $Y=2.405
+ $X2=18.435 $Y2=2.52
r15 10 11 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=18.435 $Y=2.035
+ $X2=18.435 $Y2=2.405
r16 9 10 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=18.435 $Y=1.665
+ $X2=18.435 $Y2=2.035
r17 8 9 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=18.435 $Y=1.295
+ $X2=18.435 $Y2=1.665
r18 7 8 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=18.435 $Y=0.925
+ $X2=18.435 $Y2=1.295
r19 7 22 8.72564 $w=3.48e-07 $l=2.65e-07 $layer=LI1_cond $X=18.435 $Y=0.925
+ $X2=18.435 $Y2=0.66
r20 2 13 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=18.305
+ $Y=2.375 $X2=18.445 $Y2=3.23
r21 2 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=18.305
+ $Y=2.375 $X2=18.445 $Y2=2.52
r22 1 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=18.285
+ $Y=0.535 $X2=18.425 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFSTP_1%VGND 1 2 3 4 5 6 7 22 25 34 43 56 60 69 78
+ 82
c127 60 0 1.43632e-19 $X=10.45 $Y=0.48
r128 84 86 6.42105 $w=9.48e-07 $l=5e-07 $layer=LI1_cond $X=17.57 $Y=0.66
+ $X2=17.57 $Y2=1.16
r129 79 82 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=17.21 $Y=0.44
+ $X2=17.93 $Y2=0.44
r130 78 84 2.31158 $w=9.48e-07 $l=1.8e-07 $layer=LI1_cond $X=17.57 $Y=0.48
+ $X2=17.57 $Y2=0.66
r131 78 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.93 $Y=0.48
+ $X2=17.93 $Y2=0.48
r132 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.21 $Y=0.48
+ $X2=17.21 $Y2=0.48
r133 73 79 0.654559 $w=3.7e-07 $l=1.705e-06 $layer=MET1_cond $X=15.505 $Y=0.44
+ $X2=17.21 $Y2=0.44
r134 70 73 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=14.785 $Y=0.44
+ $X2=15.505 $Y2=0.44
r135 69 75 8.15618 $w=8.88e-07 $l=5.95e-07 $layer=LI1_cond $X=15.145 $Y=0.48
+ $X2=15.145 $Y2=1.075
r136 69 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.505 $Y=0.48
+ $X2=15.505 $Y2=0.48
r137 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.785 $Y=0.48
+ $X2=14.785 $Y2=0.48
r138 64 70 1.38782 $w=3.7e-07 $l=3.615e-06 $layer=MET1_cond $X=11.17 $Y=0.44
+ $X2=14.785 $Y2=0.44
r139 61 64 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.45 $Y=0.44
+ $X2=11.17 $Y2=0.44
r140 60 66 4.04526 $w=9.48e-07 $l=3.15e-07 $layer=LI1_cond $X=10.81 $Y=0.48
+ $X2=10.81 $Y2=0.795
r141 60 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.17 $Y=0.48
+ $X2=11.17 $Y2=0.48
r142 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.45 $Y=0.48
+ $X2=10.45 $Y2=0.48
r143 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.035 $Y=0.48
+ $X2=9.035 $Y2=0.48
r144 54 56 1.06793 $w=5.58e-07 $l=5e-08 $layer=LI1_cond $X=8.985 $Y=0.645
+ $X2=9.035 $Y2=0.645
r145 51 57 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.315 $Y=0.44
+ $X2=9.035 $Y2=0.44
r146 50 54 14.3102 $w=5.58e-07 $l=6.7e-07 $layer=LI1_cond $X=8.315 $Y=0.645
+ $X2=8.985 $Y2=0.645
r147 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.315 $Y=0.48
+ $X2=8.315 $Y2=0.48
r148 44 51 1.15172 $w=3.7e-07 $l=3e-06 $layer=MET1_cond $X=5.315 $Y=0.44
+ $X2=8.315 $Y2=0.44
r149 43 47 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=5.325 $Y=0.48
+ $X2=5.325 $Y2=0.825
r150 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.315 $Y=0.48
+ $X2=5.315 $Y2=0.48
r151 38 44 0.40694 $w=3.7e-07 $l=1.06e-06 $layer=MET1_cond $X=4.255 $Y=0.44
+ $X2=5.315 $Y2=0.44
r152 35 38 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.535 $Y=0.44
+ $X2=4.255 $Y2=0.44
r153 34 40 3.40316 $w=9.48e-07 $l=2.65e-07 $layer=LI1_cond $X=3.895 $Y=0.48
+ $X2=3.895 $Y2=0.745
r154 34 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.255 $Y=0.48
+ $X2=4.255 $Y2=0.48
r155 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.535 $Y=0.48
+ $X2=3.535 $Y2=0.48
r156 29 35 0.798523 $w=3.7e-07 $l=2.08e-06 $layer=MET1_cond $X=1.455 $Y=0.44
+ $X2=3.535 $Y2=0.44
r157 26 29 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.735 $Y=0.44
+ $X2=1.455 $Y2=0.44
r158 25 31 3.40316 $w=9.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.095 $Y=0.48
+ $X2=1.095 $Y2=0.745
r159 25 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.455 $Y=0.48
+ $X2=1.455 $Y2=0.48
r160 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.735 $Y=0.48
+ $X2=0.735 $Y2=0.48
r161 22 61 0.418457 $w=3.7e-07 $l=1.09e-06 $layer=MET1_cond $X=9.36 $Y=0.44
+ $X2=10.45 $Y2=0.44
r162 22 57 0.124769 $w=3.7e-07 $l=3.25e-07 $layer=MET1_cond $X=9.36 $Y=0.44
+ $X2=9.035 $Y2=0.44
r163 7 86 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=17.39
+ $Y=0.865 $X2=17.645 $Y2=1.16
r164 7 84 182 $w=1.7e-07 $l=3.42491e-07 $layer=licon1_NDIFF $count=1 $X=17.39
+ $Y=0.865 $X2=17.645 $Y2=0.66
r165 6 75 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=14.77
+ $Y=0.865 $X2=14.91 $Y2=1.075
r166 5 66 182 $w=1.7e-07 $l=3.58748e-07 $layer=licon1_NDIFF $count=1 $X=10.885
+ $Y=0.535 $X2=11.12 $Y2=0.795
r167 4 54 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.845
+ $Y=0.565 $X2=8.985 $Y2=0.775
r168 3 47 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.24
+ $Y=0.615 $X2=5.365 $Y2=0.825
r169 2 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.895
+ $Y=0.535 $X2=4.035 $Y2=0.745
r170 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.915
+ $Y=0.535 $X2=1.055 $Y2=0.745
.ends

