* NGSPICE file created from sky130_fd_sc_hvl__conb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__conb_1 VGND VNB VPB VPWR HI LO
R0 HI VPWR short w=510000u l=45000u
R1 VGND LO short w=510000u l=45000u
.ends

