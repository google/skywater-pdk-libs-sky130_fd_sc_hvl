# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__nand2_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__nand2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.525000 2.275000 1.855000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.550000 1.015000 1.935000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.633750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.220000 1.525000 1.795000 1.695000 ;
        RECT 1.220000 1.695000 1.470000 3.755000 ;
        RECT 1.580000 1.175000 2.180000 1.345000 ;
        RECT 1.580000 1.345000 1.795000 1.525000 ;
        RECT 1.850000 0.515000 2.180000 1.175000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 2.400000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 2.400000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 2.400000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 2.400000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.985000 2.400000 4.155000 ;
      RECT 0.090000  0.365000 1.400000 1.345000 ;
      RECT 0.090000  2.175000 1.040000 3.755000 ;
      RECT 1.660000  2.175000 2.250000 3.755000 ;
    LAYER mcon ;
      RECT 0.120000  0.395000 0.290000 0.565000 ;
      RECT 0.120000  3.505000 0.290000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.480000  0.395000 0.650000 0.565000 ;
      RECT 0.480000  3.505000 0.650000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.840000  0.395000 1.010000 0.565000 ;
      RECT 0.840000  3.505000 1.010000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.200000  0.395000 1.370000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.690000  3.505000 1.860000 3.675000 ;
      RECT 2.050000  3.505000 2.220000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
  END
END sky130_fd_sc_hvl__nand2_1
