* NGSPICE file created from sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3 A SLEEP_B LVPWR VGND VNB VPB VPWR
+ X
M1000 a_362_1243# VGND VGND VNB nhv w=420000u l=500000u
+  ad=6.713e+11p pd=6.49e+06u as=1.79135e+12p ps=1.751e+07u
M1001 VGND a_1472_1171# a_840_107# VNB nhvnative w=1e+06u l=900000u
+  ad=0p pd=0u as=6.713e+11p ps=6.49e+06u
M1002 VGND a_2092_381# a_840_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_1472_1171# a_528_1171# LVPWR LVPWR phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=2.632e+12p ps=2.262e+07u
M1004 VGND a_528_1171# a_362_1243# VNB nhvnative w=1e+06u l=900000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_262_107# X VPB phv w=3e+06u l=500000u
+  ad=1.83375e+12p pd=1.512e+07u as=1.635e+12p ps=1.309e+07u
M1006 a_528_1171# a_3617_1198# LVPWR LVPWR phighvt w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1007 a_362_133# a_528_1171# a_1472_1171# VNB nshort w=740000u l=150000u
+  ad=6.882e+11p pd=6.3e+06u as=4.44e+11p ps=4.16e+06u
M1008 a_362_133# a_262_107# X VNB nhv w=1e+06u l=500000u
+  ad=8.25e+11p pd=7.65e+06u as=5.45e+11p ps=5.09e+06u
M1009 a_1472_1171# a_528_1171# a_362_133# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_362_1243# a_528_1171# VGND VNB nhvnative w=1e+06u l=900000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_262_107# X VPB phv w=3e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_362_133# a_840_107# a_262_107# VNB nhv w=1e+06u l=500000u
+  ad=0p pd=0u as=5.3e+11p ps=5.06e+06u
M1013 LVPWR a_3617_1198# a_528_1171# LVPWR phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1472_1171# a_528_1171# a_362_133# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 LVPWR a_3617_1198# a_528_1171# LVPWR phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_362_133# a_528_1171# a_1472_1171# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1410_571# a_2092_381# a_940_485# VPB phv w=3e+06u l=500000u
+  ad=2.1e+12p pd=1.668e+07u as=2.85e+12p ps=2.318e+07u
M1018 VGND a_3617_1198# a_528_1171# VNB nshort w=740000u l=150000u
+  ad=1.11e+12p pd=1.04e+07u as=4.44e+11p ps=4.16e+06u
M1019 VGND a_3617_1198# a_528_1171# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR SLEEP_B a_2092_381# VPB phv w=750000u l=500000u
+  ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u
M1021 a_940_485# a_840_107# a_262_107# VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=7.95e+11p ps=7.06e+06u
M1022 a_1410_571# a_840_107# a_362_1243# VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=3.975e+11p ps=3.53e+06u
M1023 a_362_1243# a_528_1171# VGND VNB nhvnative w=1e+06u l=900000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND A a_3617_1198# VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1025 a_528_1171# a_3617_1198# LVPWR LVPWR phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1472_1171# a_528_1171# LVPWR LVPWR phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_528_1171# a_3617_1198# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_940_485# a_2092_381# a_1410_571# VPB phv w=3e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_840_107# a_1472_1171# VGND VNB nhvnative w=1e+06u l=900000u
+  ad=0p pd=0u as=0p ps=0u
M1030 X a_262_107# a_362_133# VNB nhv w=1e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_3617_1198# A LVPWR LVPWR phighvt w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1032 a_840_107# a_1472_1171# VGND VNB nhvnative w=1e+06u l=900000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_528_1171# a_3617_1198# VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_262_107# a_840_107# a_362_133# VNB nhv w=1e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1035 LVPWR a_528_1171# a_1472_1171# LVPWR phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 X a_262_107# VPWR VPB phv w=3e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_940_485# a_2092_381# a_1410_571# VPB phv w=3e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1038 LVPWR a_528_1171# a_1472_1171# LVPWR phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1410_571# a_2092_381# a_940_485# VPB phv w=3e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND a_528_1171# a_362_1243# VNB nhvnative w=1e+06u l=900000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND a_1472_1171# a_840_107# VNB nhvnative w=1e+06u l=900000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_262_107# a_840_107# a_940_485# VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_840_107# a_362_1243# a_1410_571# VPB phv w=1.5e+06u l=500000u
+  ad=3.975e+11p pd=3.53e+06u as=0p ps=0u
M1044 LVPWR A a_3617_1198# LVPWR phighvt w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND SLEEP_B a_2092_381# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u
M1046 a_3617_1198# A VGND VNB nshort w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_362_133# a_262_107# X VNB nhv w=1e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends

