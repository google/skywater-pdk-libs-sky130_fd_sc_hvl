* File: sky130_fd_sc_hvl__o22a_1.pex.spice
* Created: Fri Aug 28 09:38:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__O22A_1%VNB 5 7 11 25
r35 7 25 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=0.057
+ $X2=2.64 $Y2=0.058
r36 7 11 0.00134943 $w=5.28e-06 $l=5.7e-08 $layer=MET1_cond $X=2.64 $Y=0.057
+ $X2=2.64 $Y2=0
r37 5 11 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r38 5 11 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__O22A_1%VPB 4 6 14 21
r37 10 21 0.00134943 $w=5.28e-06 $l=5.7e-08 $layer=MET1_cond $X=2.64 $Y=4.07
+ $X2=2.64 $Y2=4.013
r38 10 14 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=4.07
+ $X2=5.04 $Y2=4.07
r39 9 14 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=5.04
+ $Y2=4.07
r40 9 10 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r41 6 21 2.36742e-05 $w=5.28e-06 $l=1e-09 $layer=MET1_cond $X=2.64 $Y=4.012
+ $X2=2.64 $Y2=4.013
r42 4 14 33.0909 $w=1.7e-07 $l=5.08232e-06 $layer=licon1_NTAP_notbjt $count=5
+ $X=0 $Y=3.985 $X2=5.04 $Y2=4.07
r43 4 9 33.0909 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=5
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__O22A_1%A_87_81# 1 2 7 8 9 11 12 14 15 16 17 19 31
+ 35
c77 17 0 1.50932e-19 $X=3.555 $Y=2.47
r78 25 35 147.133 $w=5e-07 $l=1.375e-06 $layer=POLY_cond $X=0.685 $Y=1.59
+ $X2=0.685 $Y2=2.965
r79 25 31 72.764 $w=5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.685 $Y=1.59 $X2=0.685
+ $Y2=0.91
r80 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.59 $X2=0.75 $Y2=1.59
r81 19 21 38.4916 $w=2.48e-07 $l=8.35e-07 $layer=LI1_cond $X=3.555 $Y=2.755
+ $X2=3.555 $Y2=3.59
r82 17 29 3.14639 $w=2.5e-07 $l=1.48e-07 $layer=LI1_cond $X=3.555 $Y=2.47
+ $X2=3.555 $Y2=2.322
r83 17 19 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=3.555 $Y=2.47
+ $X2=3.555 $Y2=2.755
r84 15 27 18.0926 $w=3.63e-07 $l=5.32968e-07 $layer=LI1_cond $X=2.255 $Y=1.135
+ $X2=2.69 $Y2=0.917
r85 15 16 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.255 $Y=1.135
+ $X2=1.8 $Y2=1.135
r86 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.715 $Y=1.22
+ $X2=1.8 $Y2=1.135
r87 13 14 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.715 $Y=1.22
+ $X2=1.715 $Y2=1.425
r88 11 29 3.99677 $w=1.7e-07 $l=1.53297e-07 $layer=LI1_cond $X=3.43 $Y=2.385
+ $X2=3.555 $Y2=2.322
r89 11 12 164.08 $w=1.68e-07 $l=2.515e-06 $layer=LI1_cond $X=3.43 $Y=2.385
+ $X2=0.915 $Y2=2.385
r90 10 24 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=1.51
+ $X2=0.75 $Y2=1.51
r91 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.63 $Y=1.51
+ $X2=1.715 $Y2=1.425
r92 9 10 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.63 $Y=1.51
+ $X2=0.915 $Y2=1.51
r93 8 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.75 $Y=2.3
+ $X2=0.915 $Y2=2.385
r94 7 24 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.595 $X2=0.75
+ $Y2=1.51
r95 7 8 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=0.75 $Y=1.595
+ $X2=0.75 $Y2=2.3
r96 2 29 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.375
+ $Y=2.215 $X2=3.515 $Y2=2.34
r97 2 21 400 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=1 $X=3.375
+ $Y=2.215 $X2=3.515 $Y2=3.59
r98 2 19 400 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=3.375
+ $Y=2.215 $X2=3.515 $Y2=2.755
r99 1 27 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.55
+ $Y=0.535 $X2=2.69 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_HVL__O22A_1%A1 3 5 11 12 13 14 18 19 21 26 27 34 41 42
+ 46 52 54
c86 42 0 8.33675e-20 $X=3.13 $Y=1.305
c87 3 0 1.50932e-19 $X=4.615 $Y=2.965
r88 42 52 0.583732 $w=1.88e-07 $l=1e-08 $layer=LI1_cond $X=3.13 $Y=1.305
+ $X2=3.12 $Y2=1.305
r89 41 46 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=3.615 $Y=1.305
+ $X2=3.6 $Y2=1.305
r90 27 54 3.65058 $w=1.88e-07 $l=6e-08 $layer=LI1_cond $X=3.65 $Y=1.305 $X2=3.71
+ $Y2=1.305
r91 27 41 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=3.65 $Y=1.305
+ $X2=3.615 $Y2=1.305
r92 27 46 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=3.565 $Y=1.305
+ $X2=3.6 $Y2=1.305
r93 26 52 2.21818 $w=1.88e-07 $l=3.8e-08 $layer=LI1_cond $X=3.082 $Y=1.305
+ $X2=3.12 $Y2=1.305
r94 26 27 23.2325 $w=1.88e-07 $l=3.98e-07 $layer=LI1_cond $X=3.167 $Y=1.305
+ $X2=3.565 $Y2=1.305
r95 26 42 2.15981 $w=1.88e-07 $l=3.7e-08 $layer=LI1_cond $X=3.167 $Y=1.305
+ $X2=3.13 $Y2=1.305
r96 22 26 10.7125 $w=3.18e-07 $l=2.6e-07 $layer=LI1_cond $X=2.775 $Y=1.315
+ $X2=3.035 $Y2=1.315
r97 21 24 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.69 $Y=1.315
+ $X2=2.69 $Y2=1.485
r98 21 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.69 $Y=1.315
+ $X2=2.775 $Y2=1.315
r99 19 40 54.3061 $w=5.35e-07 $l=5.4e-07 $layer=POLY_cond $X=4.632 $Y=1.545
+ $X2=4.632 $Y2=2.085
r100 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.715
+ $Y=1.545 $X2=4.715 $Y2=1.545
r101 16 18 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=4.715 $Y=1.4
+ $X2=4.715 $Y2=1.545
r102 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.55 $Y=1.315
+ $X2=4.715 $Y2=1.4
r103 14 54 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.55 $Y=1.315
+ $X2=3.71 $Y2=1.315
r104 12 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=1.485
+ $X2=2.69 $Y2=1.485
r105 12 13 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.605 $Y=1.485
+ $X2=2.15 $Y2=1.485
r106 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.065 $Y=1.57
+ $X2=2.15 $Y2=1.485
r107 10 11 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.065 $Y=1.57
+ $X2=2.065 $Y2=1.775
r108 8 34 104.866 $w=5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.52 $Y=1.89 $X2=1.52
+ $Y2=0.91
r109 7 8 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.585
+ $Y=1.89 $X2=1.585 $Y2=1.89
r110 5 11 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.98 $Y=1.915
+ $X2=2.065 $Y2=1.775
r111 5 7 16.2577 $w=2.78e-07 $l=3.95e-07 $layer=LI1_cond $X=1.98 $Y=1.915
+ $X2=1.585 $Y2=1.915
r112 3 40 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=4.615 $Y=2.965
+ $X2=4.615 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_HVL__O22A_1%B1 3 7 9 12
c41 3 0 8.33675e-20 $X=2.3 $Y=0.91
r42 12 15 18.9925 $w=6.15e-07 $l=1.95e-07 $layer=POLY_cond $X=2.357 $Y=1.89
+ $X2=2.357 $Y2=2.085
r43 12 14 43.3516 $w=6.15e-07 $l=4.75e-07 $layer=POLY_cond $X=2.357 $Y=1.89
+ $X2=2.357 $Y2=1.415
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.495
+ $Y=1.89 $X2=2.495 $Y2=1.89
r45 9 13 4.51633 $w=3.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.64 $Y=1.935
+ $X2=2.495 $Y2=1.935
r46 7 15 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.415 $Y=2.965
+ $X2=2.415 $Y2=2.085
r47 3 14 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.3 $Y=0.91 $X2=2.3
+ $Y2=1.415
.ends

.subckt PM_SKY130_FD_SC_HVL__O22A_1%B2 1 2 6 12
r29 9 12 130.547 $w=5e-07 $l=1.22e-06 $layer=POLY_cond $X=3.125 $Y=1.745
+ $X2=3.125 $Y2=2.965
r30 6 9 89.3499 $w=5e-07 $l=8.35e-07 $layer=POLY_cond $X=3.125 $Y=0.91 $X2=3.125
+ $Y2=1.745
r31 1 2 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=3.102 $Y=1.665
+ $X2=3.102 $Y2=2.035
r32 1 9 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.1 $Y=1.745
+ $X2=3.1 $Y2=1.745
.ends

.subckt PM_SKY130_FD_SC_HVL__O22A_1%A2 1 2 6 12
r29 9 12 130.547 $w=5e-07 $l=1.22e-06 $layer=POLY_cond $X=3.905 $Y=1.745
+ $X2=3.905 $Y2=2.965
r30 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.84
+ $Y=1.745 $X2=3.84 $Y2=1.745
r31 6 9 89.3499 $w=5e-07 $l=8.35e-07 $layer=POLY_cond $X=3.905 $Y=0.91 $X2=3.905
+ $Y2=1.745
r32 2 10 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.08 $Y=1.745 $X2=3.84
+ $Y2=1.745
r33 1 10 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.6 $Y=1.745 $X2=3.84
+ $Y2=1.745
.ends

.subckt PM_SKY130_FD_SC_HVL__O22A_1%X 1 2 7 8 9 10 11 12 13 22
r14 13 40 20.1113 $w=2.53e-07 $l=4.45e-07 $layer=LI1_cond $X=0.252 $Y=3.145
+ $X2=0.252 $Y2=3.59
r15 12 13 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=2.775
+ $X2=0.252 $Y2=3.145
r16 11 12 19.6593 $w=2.53e-07 $l=4.35e-07 $layer=LI1_cond $X=0.252 $Y=2.34
+ $X2=0.252 $Y2=2.775
r17 10 11 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=0.252 $Y=2.035
+ $X2=0.252 $Y2=2.34
r18 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=1.665
+ $X2=0.252 $Y2=2.035
r19 8 9 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=1.295
+ $X2=0.252 $Y2=1.665
r20 7 8 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=0.925
+ $X2=0.252 $Y2=1.295
r21 7 22 11.9764 $w=2.53e-07 $l=2.65e-07 $layer=LI1_cond $X=0.252 $Y=0.925
+ $X2=0.252 $Y2=0.66
r22 2 40 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.215 $X2=0.295 $Y2=3.59
r23 2 11 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.215 $X2=0.295 $Y2=2.34
r24 1 22 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.535 $X2=0.295 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__O22A_1%VPWR 1 2 7 17 21 29
r35 27 29 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=3.975 $Y=3.63
+ $X2=5.055 $Y2=3.63
r36 26 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.055 $Y=3.59
+ $X2=5.055 $Y2=3.59
r37 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.975 $Y=3.59
+ $X2=3.975 $Y2=3.59
r38 24 26 0.18626 $w=1.308e-06 $l=2e-08 $layer=LI1_cond $X=4.515 $Y=3.57
+ $X2=4.515 $Y2=3.59
r39 21 24 11.2687 $w=1.308e-06 $l=1.21e-06 $layer=LI1_cond $X=4.515 $Y=2.36
+ $X2=4.515 $Y2=3.57
r40 18 27 0.310963 $w=3.7e-07 $l=8.1e-07 $layer=MET1_cond $X=3.165 $Y=3.63
+ $X2=3.975 $Y2=3.63
r41 17 18 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.165 $Y=3.59
+ $X2=3.165 $Y2=3.59
r42 14 17 23.0751 $w=1.103e-06 $l=2.09e-06 $layer=LI1_cond $X=1.075 $Y=3.202
+ $X2=3.165 $Y2=3.202
r43 10 14 4.74751 $w=1.103e-06 $l=4.3e-07 $layer=LI1_cond $X=0.645 $Y=3.202
+ $X2=1.075 $Y2=3.202
r44 10 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.645 $Y=3.59
+ $X2=0.645 $Y2=3.59
r45 7 18 0.20155 $w=3.7e-07 $l=5.25e-07 $layer=MET1_cond $X=2.64 $Y=3.63
+ $X2=3.165 $Y2=3.63
r46 7 11 0.765891 $w=3.7e-07 $l=1.995e-06 $layer=MET1_cond $X=2.64 $Y=3.63
+ $X2=0.645 $Y2=3.63
r47 2 24 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=2.215 $X2=5.005 $Y2=3.57
r48 2 21 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=2.215 $X2=5.005 $Y2=2.36
r49 1 14 400 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=2.215 $X2=1.075 $Y2=3.59
r50 1 14 400 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=2.215 $X2=1.075 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_HVL__O22A_1%VGND 1 2 7 10 19 23
r43 20 23 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=4 $Y=0.44 $X2=5.08
+ $Y2=0.44
r44 19 25 3.09692 $w=1.298e-06 $l=3.3e-07 $layer=LI1_cond $X=4.54 $Y=0.48
+ $X2=4.54 $Y2=0.81
r45 19 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.08 $Y=0.48
+ $X2=5.08 $Y2=0.48
r46 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4 $Y=0.48 $X2=4
+ $Y2=0.48
r47 11 14 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.645 $Y=0.44
+ $X2=1.365 $Y2=0.44
r48 10 16 2.46742 $w=8.88e-07 $l=1.8e-07 $layer=LI1_cond $X=1.005 $Y=0.48
+ $X2=1.005 $Y2=0.66
r49 10 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.365 $Y=0.48
+ $X2=1.365 $Y2=0.48
r50 10 11 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.645 $Y=0.48
+ $X2=0.645 $Y2=0.48
r51 7 20 0.522111 $w=3.7e-07 $l=1.36e-06 $layer=MET1_cond $X=2.64 $Y=0.44 $X2=4
+ $Y2=0.44
r52 7 14 0.489479 $w=3.7e-07 $l=1.275e-06 $layer=MET1_cond $X=2.64 $Y=0.44
+ $X2=1.365 $Y2=0.44
r53 2 25 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.155
+ $Y=0.535 $X2=4.295 $Y2=0.81
r54 1 16 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.935
+ $Y=0.535 $X2=1.075 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__O22A_1%A_354_107# 1 2 9 11 12 15
r28 13 15 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.515 $Y=0.435
+ $X2=3.515 $Y2=0.8
r29 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.35 $Y=0.35
+ $X2=3.515 $Y2=0.435
r30 11 12 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=3.35 $Y=0.35
+ $X2=2.075 $Y2=0.35
r31 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.91 $Y=0.435
+ $X2=2.075 $Y2=0.35
r32 7 9 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.91 $Y=0.435
+ $X2=1.91 $Y2=0.72
r33 2 15 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=3.375
+ $Y=0.535 $X2=3.515 $Y2=0.8
r34 1 9 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.77
+ $Y=0.535 $X2=1.91 $Y2=0.72
.ends

