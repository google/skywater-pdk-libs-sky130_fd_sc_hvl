* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbufhv2hv_hl_1 A LOWHVPWR VGND VNB VPB VPWR X
X0 X a_662_81# LOWHVPWR LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 LOWHVPWR A a_662_81# LOWHVPWR sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 X a_662_81# a_762_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X3 a_762_107# A a_662_81# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends
