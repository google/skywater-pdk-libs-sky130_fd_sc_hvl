* File: sky130_fd_sc_hvl__mux4_1.spice
* Created: Wed Sep  2 09:08:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__mux4_1.pex.spice"
.subckt sky130_fd_sc_hvl__mux4_1  VNB VPB S0 A2 A3 A1 A0 S1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S1	S1
* A0	A0
* A1	A1
* A3	A3
* A2	A2
* S0	S0
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_S0_M1020_g N_A_30_107#_M1020_s N_VNB_M1020_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250006 A=0.21 P=1.84 MULT=1
MM1006 A_339_107# N_A2_M1006_g N_VGND_M1020_d N_VNB_M1020_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84 SA=250001
+ SB=250005 A=0.21 P=1.84 MULT=1
MM1007 N_A_481_107#_M1007_d N_A_30_107#_M1007_g A_339_107# N_VNB_M1020_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1025 A_637_107# N_S0_M1025_g N_A_481_107#_M1007_d N_VNB_M1020_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250004 A=0.21 P=1.84 MULT=1
MM1002 N_VGND_M1002_d N_A3_M1002_g A_637_107# N_VNB_M1020_b NHV L=0.5 W=0.42
+ AD=0.1092 AS=0.0441 PD=0.94 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250003
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1004 A_983_107# N_A1_M1004_g N_VGND_M1002_d N_VNB_M1020_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=0.94 NRD=13.566 NRS=65.1396 M=1 R=0.84
+ SA=250004 SB=250002 A=0.21 P=1.84 MULT=1
MM1012 N_A_1097_627#_M1012_d N_S0_M1012_g A_983_107# N_VNB_M1020_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250005 SB=250002 A=0.21 P=1.84 MULT=1
MM1021 A_1281_107# N_A_30_107#_M1021_g N_A_1097_627#_M1012_d N_VNB_M1020_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250006 SB=250001 A=0.21 P=1.84 MULT=1
MM1008 N_VGND_M1008_d N_A0_M1008_g A_1281_107# N_VNB_M1020_b NHV L=0.5 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250006
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1011 N_A_1669_615#_M1011_d N_A_1681_89#_M1011_g N_A_1097_627#_M1011_s
+ N_VNB_M1020_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1005 N_A_481_107#_M1005_d N_S1_M1005_g N_A_1669_615#_M1011_d N_VNB_M1020_b NHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1010 N_VGND_M1010_d N_S1_M1010_g N_A_1681_89#_M1010_s N_VNB_M1020_b NHV L=0.5
+ W=0.42 AD=0.107638 AS=0.1197 PD=0.890256 PS=1.41 NRD=56.9886 NRS=0 M=1 R=0.84
+ SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1022 N_X_M1022_d N_A_1669_615#_M1022_g N_VGND_M1010_d N_VNB_M1020_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.192212 PD=2.03 PS=1.58974 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1013 N_VPWR_M1013_d N_S0_M1013_g N_A_30_107#_M1013_s N_VPB_M1013_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250006 A=0.21 P=1.84 MULT=1
MM1000 A_339_627# N_A2_M1000_g N_VPWR_M1013_d N_VPB_M1013_b PHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84 SA=250001
+ SB=250005 A=0.21 P=1.84 MULT=1
MM1023 N_A_481_107#_M1023_d N_S0_M1023_g A_339_627# N_VPB_M1013_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1016 A_637_627# N_A_30_107#_M1016_g N_A_481_107#_M1023_d N_VPB_M1013_b PHV
+ L=0.5 W=0.42 AD=0.0651 AS=0.0588 PD=0.73 PS=0.7 NRD=45.458 NRS=0 M=1 R=0.84
+ SA=250002 SB=250004 A=0.21 P=1.84 MULT=1
MM1009 N_VPWR_M1009_d N_A3_M1009_g A_637_627# N_VPB_M1013_b PHV L=0.5 W=0.42
+ AD=0.0588 AS=0.0651 PD=0.7 PS=0.73 NRD=0 NRS=45.458 M=1 R=0.84 SA=250003
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1024 A_955_627# N_A1_M1024_g N_VPWR_M1009_d N_VPB_M1013_b PHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84 SA=250004
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1001 N_A_1097_627#_M1001_d N_A_30_107#_M1001_g A_955_627# N_VPB_M1013_b PHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250005 SB=250002 A=0.21 P=1.84 MULT=1
MM1018 A_1253_627# N_S0_M1018_g N_A_1097_627#_M1001_d N_VPB_M1013_b PHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250005 SB=250001 A=0.21 P=1.84 MULT=1
MM1019 N_VPWR_M1019_d N_A0_M1019_g A_1253_627# N_VPB_M1013_b PHV L=0.5 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84 SA=250006
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1003 N_A_1669_615#_M1003_d N_S1_M1003_g N_A_1097_627#_M1003_s N_VPB_M1013_b
+ PHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1017 N_A_481_107#_M1017_d N_A_1681_89#_M1017_g N_A_1669_615#_M1003_d
+ N_VPB_M1013_b PHV L=0.5 W=0.42 AD=0.2751 AS=0.0588 PD=2.15 PS=0.7 NRD=168.252
+ NRS=0 M=1 R=0.84 SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1014 N_VPWR_M1014_d N_S1_M1014_g N_A_1681_89#_M1014_s N_VPB_M1013_b PHV L=0.5
+ W=0.42 AD=0.134794 AS=0.1113 PD=0.870625 PS=1.37 NRD=52.2958 NRS=0 M=1 R=0.84
+ SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1015 N_X_M1015_d N_A_1669_615#_M1015_g N_VPWR_M1014_d N_VPB_M1013_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.481406 PD=3.53 PS=3.10937 NRD=0 NRS=12.0903 M=1 R=3
+ SA=250000 SB=250000 A=0.75 P=4 MULT=1
DX26_noxref N_VNB_M1020_b N_VPB_M1013_b NWDIODE A=34.164 P=31.48
*
.include "sky130_fd_sc_hvl__mux4_1.pxi.spice"
*
.ends
*
*
