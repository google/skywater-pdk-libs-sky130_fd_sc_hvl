# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  8.140000 ;
  SYMMETRY X Y R90 ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.495000 1.530000 2.805000 2.200000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.600000 4.405000 10.930000 6.055000 ;
        RECT 10.600000 6.725000 10.930000 7.625000 ;
        RECT 10.690000 6.055000 10.930000 6.725000 ;
    END
  END X
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 10.970000 3.305000 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 11.040000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 11.040000 8.255000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 11.040000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 11.040000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.985000  0.800000 4.155000 ;
      RECT  0.000000  8.055000 11.040000 8.225000 ;
      RECT  2.885000  2.765000  3.265000 3.055000 ;
      RECT  2.885000  3.055000  3.175000 5.495000 ;
      RECT  2.975000  0.735000  3.265000 1.745000 ;
      RECT  2.975000  1.745000  4.310000 1.995000 ;
      RECT  2.975000  1.995000  3.265000 2.765000 ;
      RECT  3.095000  0.335000  4.045000 0.565000 ;
      RECT  3.145000  6.165000  3.735000 7.715000 ;
      RECT  3.145000  7.715000  5.295000 7.885000 ;
      RECT  3.345000  3.225000  4.115000 4.200000 ;
      RECT  3.435000  0.565000  3.705000 1.575000 ;
      RECT  3.435000  2.165000  3.705000 3.075000 ;
      RECT  3.435000  3.075000  4.115000 3.225000 ;
      RECT  3.875000  0.735000  4.185000 1.245000 ;
      RECT  3.875000  1.245000  4.810000 1.575000 ;
      RECT  3.875000  2.165000  5.790000 2.475000 ;
      RECT  3.875000  2.475000  4.185000 2.905000 ;
      RECT  4.055000  5.665000  7.025000 5.995000 ;
      RECT  4.055000  5.995000  4.385000 7.545000 ;
      RECT  4.480000  1.575000  4.810000 2.145000 ;
      RECT  4.480000  2.145000  5.790000 2.165000 ;
      RECT  4.705000  6.165000  5.295000 7.715000 ;
      RECT  5.050000  0.255000  7.200000 0.425000 ;
      RECT  5.050000  0.425000  5.640000 1.975000 ;
      RECT  5.960000  0.595000  6.290000 2.145000 ;
      RECT  5.960000  2.145000  7.850000 2.325000 ;
      RECT  6.565000  2.795000  6.895000 4.405000 ;
      RECT  6.565000  4.405000  7.025000 4.735000 ;
      RECT  6.610000  0.425000  7.200000 1.975000 ;
      RECT  6.695000  4.735000  7.025000 5.665000 ;
      RECT  6.695000  5.995000  7.025000 6.285000 ;
      RECT  6.695000  6.285000  8.815000 6.615000 ;
      RECT  7.095000  2.495000  9.835000 2.705000 ;
      RECT  7.095000  2.705000  7.765000 4.215000 ;
      RECT  7.390000  4.405000  7.980000 5.945000 ;
      RECT  7.520000  0.255000  9.410000 0.425000 ;
      RECT  7.520000  0.425000  7.850000 2.145000 ;
      RECT  7.955000  2.875000  8.545000 3.705000 ;
      RECT  8.170000  0.595000  8.760000 2.495000 ;
      RECT  8.235000  3.985000 11.040000 4.155000 ;
      RECT  8.300000  4.405000  8.630000 6.285000 ;
      RECT  8.535000  6.615000  8.815000 6.955000 ;
      RECT  8.915000  2.705000  9.835000 3.465000 ;
      RECT  8.995000  4.405000  9.325000 6.225000 ;
      RECT  8.995000  6.225000 10.520000 6.555000 ;
      RECT  8.995000  6.555000  9.325000 7.625000 ;
      RECT  9.080000  0.425000  9.410000 2.055000 ;
      RECT  9.690000  4.405000 10.280000 5.945000 ;
      RECT  9.690000  6.835000 10.280000 7.745000 ;
      RECT 10.125000  2.795000 10.715000 3.705000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.155000  8.055000  0.325000 8.225000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  8.055000  0.805000 8.225000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  8.055000  1.285000 8.225000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  8.055000  1.765000 8.225000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  8.055000  2.245000 8.225000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  8.055000  2.725000 8.225000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  8.055000  3.205000 8.225000 ;
      RECT  3.125000  0.365000  3.295000 0.535000 ;
      RECT  3.175000  7.545000  3.345000 7.715000 ;
      RECT  3.485000  0.425000  3.655000 0.595000 ;
      RECT  3.485000  3.050000  3.655000 3.220000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  8.055000  3.685000 8.225000 ;
      RECT  3.535000  7.545000  3.705000 7.715000 ;
      RECT  3.845000  0.365000  4.015000 0.535000 ;
      RECT  3.845000  3.105000  4.015000 3.275000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  8.055000  4.165000 8.225000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  8.055000  4.645000 8.225000 ;
      RECT  4.735000  7.545000  4.905000 7.715000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  8.055000  5.125000 8.225000 ;
      RECT  5.080000  0.425000  5.250000 0.595000 ;
      RECT  5.095000  7.545000  5.265000 7.715000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  8.055000  5.605000 8.225000 ;
      RECT  5.440000  0.425000  5.610000 0.595000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  8.055000  6.085000 8.225000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  8.055000  6.565000 8.225000 ;
      RECT  6.640000  0.425000  6.810000 0.595000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  8.055000  7.045000 8.225000 ;
      RECT  7.000000  0.425000  7.170000 0.595000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  8.055000  7.525000 8.225000 ;
      RECT  7.420000  4.495000  7.590000 4.665000 ;
      RECT  7.780000  4.495000  7.950000 4.665000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  8.055000  8.005000 8.225000 ;
      RECT  7.985000  3.475000  8.155000 3.645000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.315000  8.055000  8.485000 8.225000 ;
      RECT  8.345000  3.475000  8.515000 3.645000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.795000  8.055000  8.965000 8.225000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.275000  8.055000  9.445000 8.225000 ;
      RECT  9.720000  4.495000  9.890000 4.665000 ;
      RECT  9.720000  7.545000  9.890000 7.715000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.755000  8.055000  9.925000 8.225000 ;
      RECT 10.080000  4.495000 10.250000 4.665000 ;
      RECT 10.080000  7.545000 10.250000 7.715000 ;
      RECT 10.155000  3.475000 10.325000 3.645000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.235000  8.055000 10.405000 8.225000 ;
      RECT 10.515000  3.475000 10.685000 3.645000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.715000  8.055000 10.885000 8.225000 ;
    LAYER met1 ;
      RECT 0.000000 -0.115000 11.040000 0.115000 ;
      RECT 0.000000  0.255000 11.040000 0.625000 ;
      RECT 0.000000  3.445000 11.040000 3.815000 ;
  END
END sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1
END LIBRARY
