* File: sky130_fd_sc_hvl__a22oi_1.pxi.spice
* Created: Wed Sep  2 09:03:30 2020
* 
x_PM_SKY130_FD_SC_HVL__A22OI_1%VNB N_VNB_M1003_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__A22OI_1%VNB
x_PM_SKY130_FD_SC_HVL__A22OI_1%VPB N_VPB_M1004_b VPB N_VPB_c_26_p VPB
+ PM_SKY130_FD_SC_HVL__A22OI_1%VPB
x_PM_SKY130_FD_SC_HVL__A22OI_1%B2 N_B2_M1004_g N_B2_M1003_g B2 B2 N_B2_c_63_n
+ PM_SKY130_FD_SC_HVL__A22OI_1%B2
x_PM_SKY130_FD_SC_HVL__A22OI_1%B1 N_B1_M1005_g N_B1_M1007_g B1 N_B1_c_91_n
+ PM_SKY130_FD_SC_HVL__A22OI_1%B1
x_PM_SKY130_FD_SC_HVL__A22OI_1%A1 A1 A1 N_A1_M1001_g N_A1_M1006_g
+ PM_SKY130_FD_SC_HVL__A22OI_1%A1
x_PM_SKY130_FD_SC_HVL__A22OI_1%A2 N_A2_M1002_g N_A2_M1000_g A2 A2 N_A2_c_158_n
+ PM_SKY130_FD_SC_HVL__A22OI_1%A2
x_PM_SKY130_FD_SC_HVL__A22OI_1%A_33_443# N_A_33_443#_M1004_s N_A_33_443#_M1007_d
+ N_A_33_443#_M1000_d N_A_33_443#_c_177_n N_A_33_443#_c_178_n
+ N_A_33_443#_c_181_n N_A_33_443#_c_184_n N_A_33_443#_c_185_n
+ N_A_33_443#_c_186_n N_A_33_443#_c_187_n PM_SKY130_FD_SC_HVL__A22OI_1%A_33_443#
x_PM_SKY130_FD_SC_HVL__A22OI_1%Y N_Y_M1005_d N_Y_M1004_d N_Y_c_224_n N_Y_c_239_n
+ N_Y_c_226_n Y Y Y Y Y Y Y N_Y_c_236_n Y PM_SKY130_FD_SC_HVL__A22OI_1%Y
x_PM_SKY130_FD_SC_HVL__A22OI_1%VPWR N_VPWR_M1006_d VPWR N_VPWR_c_270_n
+ N_VPWR_c_273_n PM_SKY130_FD_SC_HVL__A22OI_1%VPWR
x_PM_SKY130_FD_SC_HVL__A22OI_1%VGND N_VGND_M1003_s N_VGND_M1002_d VGND
+ N_VGND_c_295_n N_VGND_c_297_n N_VGND_c_299_n PM_SKY130_FD_SC_HVL__A22OI_1%VGND
cc_1 N_VNB_M1003_b N_B2_M1003_g 0.0515897f $X=-0.33 $Y=-0.265 $X2=0.77 $Y2=0.91
cc_2 N_VNB_c_2_p N_B2_M1003_g 0.00158722f $X=0.24 $Y=0 $X2=0.77 $Y2=0.91
cc_3 N_VNB_M1003_b B2 0.0227556f $X=-0.33 $Y=-0.265 $X2=0.635 $Y2=1.58
cc_4 N_VNB_M1003_b N_B2_c_63_n 0.0551137f $X=-0.33 $Y=-0.265 $X2=0.635 $Y2=1.67
cc_5 N_VNB_M1003_b N_B1_M1005_g 0.0488073f $X=-0.33 $Y=-0.265 $X2=0.7 $Y2=2.965
cc_6 N_VNB_c_2_p N_B1_M1005_g 0.0023273f $X=0.24 $Y=0 $X2=0.7 $Y2=2.965
cc_7 N_VNB_M1003_b N_B1_c_91_n 0.0428652f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_8 N_VNB_M1003_b A1 0.00395482f $X=-0.33 $Y=-0.265 $X2=0.7 $Y2=2.965
cc_9 N_VNB_M1003_b N_A1_M1001_g 0.0802199f $X=-0.33 $Y=-0.265 $X2=0.77 $Y2=0.91
cc_10 N_VNB_c_2_p N_A1_M1001_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.77 $Y2=0.91
cc_11 N_VNB_M1003_b N_A2_M1002_g 0.0431665f $X=-0.33 $Y=-0.265 $X2=0.7 $Y2=2.965
cc_12 N_VNB_M1003_b A2 0.0232779f $X=-0.33 $Y=-0.265 $X2=0.635 $Y2=1.58
cc_13 N_VNB_M1003_b N_A2_c_158_n 0.0557118f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.67
cc_14 N_VNB_M1003_b N_Y_c_224_n 0.00864253f $X=-0.33 $Y=-0.265 $X2=0.155
+ $Y2=1.58
cc_15 N_VNB_c_2_p N_Y_c_224_n 6.32535e-19 $X=0.24 $Y=0 $X2=0.155 $Y2=1.58
cc_16 N_VNB_M1003_b N_Y_c_226_n 0.00326934f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.67
cc_17 N_VNB_M1003_b Y 0.00462661f $X=-0.33 $Y=-0.265 $X2=0.635 $Y2=1.67
cc_18 N_VNB_M1003_b N_VGND_c_295_n 0.0712556f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.58
cc_19 N_VNB_c_2_p N_VGND_c_295_n 0.00166879f $X=0.24 $Y=0 $X2=0.635 $Y2=1.58
cc_20 N_VNB_M1003_b N_VGND_c_297_n 0.12799f $X=-0.33 $Y=-0.265 $X2=0.735
+ $Y2=2.085
cc_21 N_VNB_c_2_p N_VGND_c_297_n 0.00457781f $X=0.24 $Y=0 $X2=0.735 $Y2=2.085
cc_22 N_VNB_M1003_b N_VGND_c_299_n 0.0719343f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.67
cc_23 N_VNB_c_2_p N_VGND_c_299_n 0.410664f $X=0.24 $Y=0 $X2=0.635 $Y2=1.67
cc_24 N_VPB_M1004_b N_B2_M1004_g 0.0410728f $X=-0.33 $Y=1.885 $X2=0.7 $Y2=2.965
cc_25 VPB N_B2_M1004_g 0.00970178f $X=0 $Y=3.955 $X2=0.7 $Y2=2.965
cc_26 N_VPB_c_26_p N_B2_M1004_g 0.0134683f $X=3.6 $Y=4.07 $X2=0.7 $Y2=2.965
cc_27 N_VPB_M1004_b N_B2_c_63_n 0.0280136f $X=-0.33 $Y=1.885 $X2=0.635 $Y2=1.67
cc_28 N_VPB_M1004_b N_B1_M1007_g 0.0468862f $X=-0.33 $Y=1.885 $X2=0.77 $Y2=0.91
cc_29 VPB N_B1_M1007_g 0.00970178f $X=0 $Y=3.955 $X2=0.77 $Y2=0.91
cc_30 N_VPB_c_26_p N_B1_M1007_g 0.0134683f $X=3.6 $Y=4.07 $X2=0.77 $Y2=0.91
cc_31 N_VPB_M1004_b N_B1_c_91_n 0.00430391f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_32 N_VPB_M1004_b N_A1_M1001_g 0.0513018f $X=-0.33 $Y=1.885 $X2=0.77 $Y2=0.91
cc_33 VPB N_A1_M1001_g 0.00970178f $X=0 $Y=3.955 $X2=0.77 $Y2=0.91
cc_34 N_VPB_c_26_p N_A1_M1001_g 0.0152133f $X=3.6 $Y=4.07 $X2=0.77 $Y2=0.91
cc_35 N_VPB_M1004_b N_A2_M1000_g 0.0393796f $X=-0.33 $Y=1.885 $X2=0.77 $Y2=0.91
cc_36 VPB N_A2_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.77 $Y2=0.91
cc_37 N_VPB_c_26_p N_A2_M1000_g 0.0158814f $X=3.6 $Y=4.07 $X2=0.77 $Y2=0.91
cc_38 N_VPB_M1004_b N_A2_c_158_n 0.0232969f $X=-0.33 $Y=1.885 $X2=0.635 $Y2=1.67
cc_39 N_VPB_M1004_b N_A_33_443#_c_177_n 0.054709f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_40 N_VPB_M1004_b N_A_33_443#_c_178_n 0.00275086f $X=-0.33 $Y=1.885 $X2=0.735
+ $Y2=1.415
cc_41 VPB N_A_33_443#_c_178_n 0.00596296f $X=0 $Y=3.955 $X2=0.735 $Y2=1.415
cc_42 N_VPB_c_26_p N_A_33_443#_c_178_n 0.0949207f $X=3.6 $Y=4.07 $X2=0.735
+ $Y2=1.415
cc_43 N_VPB_M1004_b N_A_33_443#_c_181_n 0.00377064f $X=-0.33 $Y=1.885 $X2=0.735
+ $Y2=2.085
cc_44 VPB N_A_33_443#_c_181_n 0.00113681f $X=0 $Y=3.955 $X2=0.735 $Y2=2.085
cc_45 N_VPB_c_26_p N_A_33_443#_c_181_n 0.0222211f $X=3.6 $Y=4.07 $X2=0.735
+ $Y2=2.085
cc_46 N_VPB_M1004_b N_A_33_443#_c_184_n 0.00107607f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.67
cc_47 N_VPB_M1004_b N_A_33_443#_c_185_n 0.0189244f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_48 N_VPB_M1004_b N_A_33_443#_c_186_n 0.00296772f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_49 N_VPB_M1004_b N_A_33_443#_c_187_n 0.0571973f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_50 VPB N_A_33_443#_c_187_n 0.00104693f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_51 N_VPB_c_26_p N_A_33_443#_c_187_n 0.0172373f $X=3.6 $Y=4.07 $X2=0 $Y2=0
cc_52 N_VPB_M1004_b Y 0.00271084f $X=-0.33 $Y=1.885 $X2=0.635 $Y2=1.67
cc_53 N_VPB_M1004_b Y 0.00340939f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_54 N_VPB_M1004_b N_VPWR_c_270_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0.77
+ $Y2=0.91
cc_55 VPB N_VPWR_c_270_n 0.00406397f $X=0 $Y=3.955 $X2=0.77 $Y2=0.91
cc_56 N_VPB_c_26_p N_VPWR_c_270_n 0.047451f $X=3.6 $Y=4.07 $X2=0.77 $Y2=0.91
cc_57 N_VPB_M1004_b N_VPWR_c_273_n 0.0534948f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.67
cc_58 VPB N_VPWR_c_273_n 0.406982f $X=0 $Y=3.955 $X2=0.635 $Y2=1.67
cc_59 N_VPB_c_26_p N_VPWR_c_273_n 0.0158275f $X=3.6 $Y=4.07 $X2=0.635 $Y2=1.67
cc_60 N_B2_M1003_g N_B1_M1005_g 0.0555749f $X=0.77 $Y=0.91 $X2=0 $Y2=0
cc_61 N_B2_M1004_g N_B1_M1007_g 0.0195539f $X=0.7 $Y=2.965 $X2=0 $Y2=0
cc_62 B2 N_B1_c_91_n 2.47254e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_63 N_B2_c_63_n N_B1_c_91_n 0.0555749f $X=0.635 $Y=1.67 $X2=0 $Y2=0
cc_64 N_B2_M1004_g N_A_33_443#_c_177_n 0.0409222f $X=0.7 $Y=2.965 $X2=0 $Y2=0
cc_65 B2 N_A_33_443#_c_177_n 0.01771f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_66 N_B2_M1004_g N_A_33_443#_c_178_n 0.0214561f $X=0.7 $Y=2.965 $X2=3.6 $Y2=0
cc_67 N_B2_M1004_g N_A_33_443#_c_181_n 0.00223748f $X=0.7 $Y=2.965 $X2=3.6 $Y2=0
cc_68 N_B2_M1003_g N_Y_c_224_n 0.00113617f $X=0.77 $Y=0.91 $X2=0 $Y2=0
cc_69 N_B2_M1004_g Y 0.00208322f $X=0.7 $Y=2.965 $X2=0 $Y2=0
cc_70 N_B2_M1003_g Y 0.0168225f $X=0.77 $Y=0.91 $X2=0 $Y2=0
cc_71 B2 Y 0.0198905f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_72 N_B2_M1004_g Y 0.00645595f $X=0.7 $Y=2.965 $X2=0 $Y2=0
cc_73 N_B2_c_63_n Y 0.00369494f $X=0.635 $Y=1.67 $X2=0 $Y2=0
cc_74 N_B2_M1003_g N_Y_c_236_n 0.00209596f $X=0.77 $Y=0.91 $X2=0 $Y2=0
cc_75 N_B2_M1004_g Y 0.0290626f $X=0.7 $Y=2.965 $X2=0 $Y2=0
cc_76 N_B2_M1004_g N_VPWR_c_273_n 0.0231873f $X=0.7 $Y=2.965 $X2=0 $Y2=0
cc_77 N_B2_M1003_g N_VGND_c_295_n 0.0421303f $X=0.77 $Y=0.91 $X2=0.24 $Y2=0
cc_78 B2 N_VGND_c_295_n 0.0453819f $X=0.635 $Y=1.58 $X2=0.24 $Y2=0
cc_79 N_B2_c_63_n N_VGND_c_295_n 0.00211209f $X=0.635 $Y=1.67 $X2=0.24 $Y2=0
cc_80 N_B2_M1003_g N_VGND_c_299_n 0.0224116f $X=0.77 $Y=0.91 $X2=1.92 $Y2=0
cc_81 B1 A1 0.0143333f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_82 N_B1_c_91_n A1 8.89781e-19 $X=1.63 $Y=1.625 $X2=0 $Y2=0
cc_83 N_B1_M1005_g N_A1_M1001_g 0.0186731f $X=1.48 $Y=0.91 $X2=0 $Y2=0
cc_84 N_B1_M1007_g N_A1_M1001_g 0.0239388f $X=1.48 $Y=2.965 $X2=0 $Y2=0
cc_85 B1 N_A1_M1001_g 9.317e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_86 N_B1_c_91_n N_A1_M1001_g 0.0365739f $X=1.63 $Y=1.625 $X2=0 $Y2=0
cc_87 N_B1_M1007_g N_A_33_443#_c_178_n 0.0222208f $X=1.48 $Y=2.965 $X2=3.6 $Y2=0
cc_88 N_B1_M1007_g N_A_33_443#_c_184_n 0.0400904f $X=1.48 $Y=2.965 $X2=1.92
+ $Y2=0
cc_89 N_B1_M1007_g N_A_33_443#_c_186_n 0.00668511f $X=1.48 $Y=2.965 $X2=1.92
+ $Y2=0.058
cc_90 B1 N_A_33_443#_c_186_n 0.00701076f $X=1.595 $Y=1.58 $X2=1.92 $Y2=0.058
cc_91 N_B1_c_91_n N_A_33_443#_c_186_n 0.002196f $X=1.63 $Y=1.625 $X2=1.92
+ $Y2=0.058
cc_92 N_B1_M1005_g N_Y_c_224_n 0.00812791f $X=1.48 $Y=0.91 $X2=0 $Y2=0
cc_93 N_B1_M1005_g N_Y_c_239_n 0.0267476f $X=1.48 $Y=0.91 $X2=0 $Y2=0
cc_94 B1 N_Y_c_239_n 0.00663973f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_95 N_B1_M1005_g N_Y_c_226_n 0.0099212f $X=1.48 $Y=0.91 $X2=0 $Y2=0
cc_96 B1 N_Y_c_226_n 0.00693648f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_97 N_B1_c_91_n N_Y_c_226_n 0.00199898f $X=1.63 $Y=1.625 $X2=0 $Y2=0
cc_98 N_B1_M1005_g Y 0.0157222f $X=1.48 $Y=0.91 $X2=0 $Y2=0
cc_99 N_B1_M1007_g Y 0.00900347f $X=1.48 $Y=2.965 $X2=0 $Y2=0
cc_100 B1 Y 0.0168581f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_101 N_B1_c_91_n Y 0.0196976f $X=1.63 $Y=1.625 $X2=0 $Y2=0
cc_102 N_B1_M1007_g Y 0.00555411f $X=1.48 $Y=2.965 $X2=0 $Y2=0
cc_103 N_B1_M1005_g N_Y_c_236_n 0.00276601f $X=1.48 $Y=0.91 $X2=0 $Y2=0
cc_104 N_B1_M1007_g Y 0.031404f $X=1.48 $Y=2.965 $X2=0 $Y2=0
cc_105 N_B1_M1007_g N_VPWR_c_270_n 6.22341e-19 $X=1.48 $Y=2.965 $X2=0 $Y2=0
cc_106 N_B1_M1007_g N_VPWR_c_273_n 0.0216437f $X=1.48 $Y=2.965 $X2=0 $Y2=0
cc_107 N_B1_M1005_g N_VGND_c_295_n 0.00236145f $X=1.48 $Y=0.91 $X2=0.24 $Y2=0
cc_108 N_B1_M1005_g N_VGND_c_297_n 0.00114166f $X=1.48 $Y=0.91 $X2=3.6 $Y2=0
cc_109 N_B1_M1005_g N_VGND_c_299_n 0.01539f $X=1.48 $Y=0.91 $X2=1.92 $Y2=0
cc_110 N_A1_M1001_g N_A2_M1002_g 0.114738f $X=2.26 $Y=0.91 $X2=0 $Y2=0
cc_111 N_A1_M1001_g N_A2_M1000_g 0.0169765f $X=2.26 $Y=0.91 $X2=0 $Y2=0
cc_112 A1 A2 0.0192701f $X=2.555 $Y=1.58 $X2=0.24 $Y2=0
cc_113 A1 N_A2_c_158_n 0.00770185f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A1_M1001_g N_A_33_443#_c_178_n 0.00161577f $X=2.26 $Y=0.91 $X2=3.6
+ $Y2=0
cc_115 N_A1_M1001_g N_A_33_443#_c_184_n 0.00375436f $X=2.26 $Y=0.91 $X2=1.92
+ $Y2=0
cc_116 A1 N_A_33_443#_c_185_n 0.0489292f $X=2.555 $Y=1.58 $X2=1.92 $Y2=0.058
cc_117 N_A1_M1001_g N_A_33_443#_c_185_n 0.0304124f $X=2.26 $Y=0.91 $X2=1.92
+ $Y2=0.058
cc_118 N_A1_M1001_g N_Y_c_224_n 3.88512e-19 $X=2.26 $Y=0.91 $X2=0 $Y2=0
cc_119 N_A1_M1001_g N_Y_c_226_n 3.46334e-19 $X=2.26 $Y=0.91 $X2=0 $Y2=0
cc_120 N_A1_M1001_g N_VPWR_c_270_n 0.0712157f $X=2.26 $Y=0.91 $X2=0 $Y2=0
cc_121 N_A1_M1001_g N_VPWR_c_273_n 0.00783253f $X=2.26 $Y=0.91 $X2=0 $Y2=0
cc_122 A1 N_VGND_c_297_n 0.0479872f $X=2.555 $Y=1.58 $X2=3.6 $Y2=0
cc_123 N_A1_M1001_g N_VGND_c_297_n 0.0599913f $X=2.26 $Y=0.91 $X2=3.6 $Y2=0
cc_124 N_A1_M1001_g N_VGND_c_299_n 0.00778503f $X=2.26 $Y=0.91 $X2=1.92 $Y2=0
cc_125 N_A2_M1000_g N_A_33_443#_c_185_n 0.0131445f $X=3.04 $Y=2.965 $X2=1.92
+ $Y2=0.058
cc_126 A2 N_A_33_443#_c_185_n 0.0488517f $X=3.515 $Y=1.58 $X2=1.92 $Y2=0.058
cc_127 N_A2_c_158_n N_A_33_443#_c_185_n 0.024281f $X=3.105 $Y=1.63 $X2=1.92
+ $Y2=0.058
cc_128 N_A2_M1000_g N_A_33_443#_c_187_n 0.0357986f $X=3.04 $Y=2.965 $X2=0 $Y2=0
cc_129 N_A2_M1000_g N_VPWR_c_270_n 0.0674428f $X=3.04 $Y=2.965 $X2=0 $Y2=0
cc_130 N_A2_c_158_n N_VPWR_c_270_n 3.48699e-19 $X=3.105 $Y=1.63 $X2=0 $Y2=0
cc_131 N_A2_M1000_g N_VPWR_c_273_n 0.010606f $X=3.04 $Y=2.965 $X2=0 $Y2=0
cc_132 N_A2_M1002_g N_VGND_c_297_n 0.0754742f $X=2.97 $Y=0.91 $X2=3.6 $Y2=0
cc_133 A2 N_VGND_c_297_n 0.0617855f $X=3.515 $Y=1.58 $X2=3.6 $Y2=0
cc_134 N_A2_c_158_n N_VGND_c_297_n 0.00211209f $X=3.105 $Y=1.63 $X2=3.6 $Y2=0
cc_135 N_A_33_443#_c_178_n N_Y_M1004_d 8.28689e-19 $X=1.705 $Y=3.72 $X2=0 $Y2=0
cc_136 N_A_33_443#_c_186_n N_Y_c_226_n 0.00612234f $X=1.955 $Y=2.015 $X2=3.6
+ $Y2=4.07
cc_137 N_A_33_443#_c_184_n Y 0.047981f $X=1.87 $Y=2.34 $X2=3.6 $Y2=4.07
cc_138 N_A_33_443#_c_186_n Y 0.00629234f $X=1.955 $Y=2.015 $X2=3.6 $Y2=4.07
cc_139 N_A_33_443#_c_177_n Y 0.0437718f $X=0.31 $Y=2.34 $X2=0 $Y2=0
cc_140 N_A_33_443#_c_178_n Y 0.0197284f $X=1.705 $Y=3.72 $X2=0 $Y2=0
cc_141 N_A_33_443#_c_178_n N_VPWR_c_270_n 0.00650116f $X=1.705 $Y=3.72 $X2=0
+ $Y2=0
cc_142 N_A_33_443#_c_184_n N_VPWR_c_270_n 0.0556936f $X=1.87 $Y=2.34 $X2=0 $Y2=0
cc_143 N_A_33_443#_c_185_n N_VPWR_c_270_n 0.0658158f $X=3.265 $Y=2.015 $X2=0
+ $Y2=0
cc_144 N_A_33_443#_c_187_n N_VPWR_c_270_n 0.107449f $X=3.43 $Y=2.34 $X2=0 $Y2=0
cc_145 N_A_33_443#_M1007_d N_VPWR_c_273_n 0.00221032f $X=1.73 $Y=2.215 $X2=3.6
+ $Y2=4.07
cc_146 N_A_33_443#_c_177_n N_VPWR_c_273_n 0.035897f $X=0.31 $Y=2.34 $X2=3.6
+ $Y2=4.07
cc_147 N_A_33_443#_c_178_n N_VPWR_c_273_n 0.0522119f $X=1.705 $Y=3.72 $X2=3.6
+ $Y2=4.07
cc_148 N_A_33_443#_c_181_n N_VPWR_c_273_n 0.0113189f $X=0.475 $Y=3.72 $X2=3.6
+ $Y2=4.07
cc_149 N_A_33_443#_c_184_n N_VPWR_c_273_n 0.0265865f $X=1.87 $Y=2.34 $X2=3.6
+ $Y2=4.07
cc_150 N_A_33_443#_c_187_n N_VPWR_c_273_n 0.0442247f $X=3.43 $Y=2.34 $X2=3.6
+ $Y2=4.07
cc_151 N_A_33_443#_c_185_n N_VGND_c_297_n 0.00491237f $X=3.265 $Y=2.015 $X2=0
+ $Y2=0
cc_152 Y N_VPWR_c_273_n 0.0249982f $X=1.2 $Y=2.405 $X2=0 $Y2=0
cc_153 Y N_VGND_c_295_n 0.0138271f $X=1.115 $Y=0.84 $X2=0.24 $Y2=0
cc_154 N_Y_c_236_n N_VGND_c_295_n 0.00747777f $X=1.185 $Y=0.98 $X2=0.24 $Y2=0
cc_155 N_Y_c_224_n N_VGND_c_297_n 0.0142624f $X=1.87 $Y=0.66 $X2=3.6 $Y2=0
cc_156 N_Y_c_226_n N_VGND_c_297_n 0.0153104f $X=1.83 $Y=0.895 $X2=3.6 $Y2=0
cc_157 N_Y_M1005_d N_VGND_c_299_n 0.00221032f $X=1.73 $Y=0.535 $X2=1.92 $Y2=0
cc_158 N_Y_c_224_n N_VGND_c_299_n 0.0265242f $X=1.87 $Y=0.66 $X2=1.92 $Y2=0
cc_159 N_Y_c_239_n N_VGND_c_299_n 0.0174486f $X=1.705 $Y=0.895 $X2=1.92 $Y2=0
cc_160 N_Y_c_236_n N_VGND_c_299_n 0.0108538f $X=1.185 $Y=0.98 $X2=1.92 $Y2=0
cc_161 Y A_204_107# 0.00356248f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_162 N_Y_c_236_n A_204_107# 0.00343956f $X=1.185 $Y=0.98 $X2=0 $Y2=0
cc_163 N_VGND_c_299_n A_204_107# 0.0039851f $X=3.66 $Y=0.48 $X2=0 $Y2=0
