* NGSPICE file created from sky130_fd_sc_hvl__inv_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__inv_1 A VGND VNB VPB VPWR Y
M1000 Y A VPWR VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=4.275e+11p ps=3.57e+06u
M1001 Y A VGND VNB nhv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=2.1375e+11p ps=2.07e+06u
.ends

