* File: sky130_fd_sc_hvl__inv_8.pex.spice
* Created: Fri Aug 28 09:36:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__INV_8%VNB 5 7 11 25
c27 11 0 3.8543e-21 $X=0.24 $Y=0
r28 7 25 1.73611e-05 $w=7.2e-06 $l=1e-09 $layer=MET1_cond $X=3.6 $Y=0.057
+ $X2=3.6 $Y2=0.058
r29 7 11 0.000989583 $w=7.2e-06 $l=5.7e-08 $layer=MET1_cond $X=3.6 $Y=0.057
+ $X2=3.6 $Y2=0
r30 5 11 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r31 5 11 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_8%VPB 4 6 14 21
r58 10 21 0.000989583 $w=7.2e-06 $l=5.7e-08 $layer=MET1_cond $X=3.6 $Y=4.07
+ $X2=3.6 $Y2=4.013
r59 10 14 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=6.96 $Y=4.07
+ $X2=6.96 $Y2=4.07
r60 9 14 438.417 $w=1.68e-07 $l=6.72e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=6.96 $Y2=4.07
r61 9 10 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r62 6 21 1.73611e-05 $w=7.2e-06 $l=1e-09 $layer=MET1_cond $X=3.6 $Y=4.012
+ $X2=3.6 $Y2=4.013
r63 4 14 24.2667 $w=1.7e-07 $l=7.00237e-06 $layer=licon1_NTAP_notbjt $count=7
+ $X=0 $Y=3.985 $X2=6.96 $Y2=4.07
r64 4 9 24.2667 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=7
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_8%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34 36
+ 38 41 43 45 48 50 52 55 57 58 59 60 61 62 63 90 91
c178 1 0 3.8543e-21 $X=0.91 $Y=1.565
r179 90 91 15.2926 $w=1.7e-07 $l=1.615e-06 $layer=licon1_POLY $count=9 $X=6.595
+ $Y=1.73 $X2=6.595 $Y2=1.73
r180 88 90 9.0955 $w=5e-07 $l=8.5e-08 $layer=POLY_cond $X=6.51 $Y=1.815
+ $X2=6.595 $Y2=1.815
r181 87 88 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=5.73 $Y=1.815
+ $X2=6.51 $Y2=1.815
r182 86 87 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=4.95 $Y=1.815
+ $X2=5.73 $Y2=1.815
r183 85 86 14.9808 $w=5e-07 $l=1.4e-07 $layer=POLY_cond $X=4.81 $Y=1.815
+ $X2=4.95 $Y2=1.815
r184 84 85 68.4838 $w=5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.17 $Y=1.815
+ $X2=4.81 $Y2=1.815
r185 83 84 14.9808 $w=5e-07 $l=1.4e-07 $layer=POLY_cond $X=4.03 $Y=1.815
+ $X2=4.17 $Y2=1.815
r186 82 83 68.4838 $w=5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.39 $Y=1.815
+ $X2=4.03 $Y2=1.815
r187 81 82 14.9808 $w=5e-07 $l=1.4e-07 $layer=POLY_cond $X=3.25 $Y=1.815
+ $X2=3.39 $Y2=1.815
r188 80 81 68.4838 $w=5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.61 $Y=1.815
+ $X2=3.25 $Y2=1.815
r189 79 80 14.9808 $w=5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.47 $Y=1.815
+ $X2=2.61 $Y2=1.815
r190 78 79 68.4838 $w=5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.83 $Y=1.815
+ $X2=2.47 $Y2=1.815
r191 77 78 14.9808 $w=5e-07 $l=1.4e-07 $layer=POLY_cond $X=1.69 $Y=1.815
+ $X2=1.83 $Y2=1.815
r192 76 77 68.4838 $w=5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.05 $Y=1.815
+ $X2=1.69 $Y2=1.815
r193 75 76 14.9808 $w=5e-07 $l=1.4e-07 $layer=POLY_cond $X=0.91 $Y=1.815
+ $X2=1.05 $Y2=1.815
r194 72 75 46.5476 $w=5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=1.815
+ $X2=0.91 $Y2=1.815
r195 72 73 15.2926 $w=1.7e-07 $l=1.615e-06 $layer=licon1_POLY $count=9 $X=0.475
+ $Y=1.73 $X2=0.475 $Y2=1.73
r196 63 91 99.7967 $w=2.33e-07 $l=2.035e-06 $layer=LI1_cond $X=4.56 $Y=1.697
+ $X2=6.595 $Y2=1.697
r197 62 63 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.697
+ $X2=4.56 $Y2=1.697
r198 61 62 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.697
+ $X2=4.08 $Y2=1.697
r199 60 61 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.697
+ $X2=3.6 $Y2=1.697
r200 59 60 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.697
+ $X2=3.12 $Y2=1.697
r201 58 59 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.697
+ $X2=2.64 $Y2=1.697
r202 57 58 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.697
+ $X2=2.16 $Y2=1.697
r203 57 73 59.0934 $w=2.33e-07 $l=1.205e-06 $layer=LI1_cond $X=1.68 $Y=1.697
+ $X2=0.475 $Y2=1.697
r204 53 88 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.51 $Y=2.065
+ $X2=6.51 $Y2=1.815
r205 53 55 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=6.51 $Y=2.065 $X2=6.51
+ $Y2=2.965
r206 50 88 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.51 $Y=1.565
+ $X2=6.51 $Y2=1.815
r207 50 52 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.51 $Y=1.565
+ $X2=6.51 $Y2=1.08
r208 46 87 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.73 $Y=2.065
+ $X2=5.73 $Y2=1.815
r209 46 48 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=5.73 $Y=2.065 $X2=5.73
+ $Y2=2.965
r210 43 87 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.73 $Y=1.565
+ $X2=5.73 $Y2=1.815
r211 43 45 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=5.73 $Y=1.565
+ $X2=5.73 $Y2=1.08
r212 39 86 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.95 $Y=2.065
+ $X2=4.95 $Y2=1.815
r213 39 41 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=4.95 $Y=2.065 $X2=4.95
+ $Y2=2.965
r214 36 85 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.81 $Y=1.565
+ $X2=4.81 $Y2=1.815
r215 36 38 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.81 $Y=1.565
+ $X2=4.81 $Y2=1.08
r216 32 84 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.17 $Y=2.065
+ $X2=4.17 $Y2=1.815
r217 32 34 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=4.17 $Y=2.065 $X2=4.17
+ $Y2=2.965
r218 29 83 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.03 $Y=1.565
+ $X2=4.03 $Y2=1.815
r219 29 31 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.03 $Y=1.565
+ $X2=4.03 $Y2=1.08
r220 25 82 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.39 $Y=2.065
+ $X2=3.39 $Y2=1.815
r221 25 27 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=3.39 $Y=2.065 $X2=3.39
+ $Y2=2.965
r222 22 81 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.25 $Y=1.565
+ $X2=3.25 $Y2=1.815
r223 22 24 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.25 $Y=1.565
+ $X2=3.25 $Y2=1.08
r224 18 80 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.61 $Y=2.065
+ $X2=2.61 $Y2=1.815
r225 18 20 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=2.61 $Y=2.065 $X2=2.61
+ $Y2=2.965
r226 15 79 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.47 $Y=1.565
+ $X2=2.47 $Y2=1.815
r227 15 17 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.47 $Y=1.565
+ $X2=2.47 $Y2=1.08
r228 11 78 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.83 $Y=2.065
+ $X2=1.83 $Y2=1.815
r229 11 13 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=1.83 $Y=2.065 $X2=1.83
+ $Y2=2.965
r230 8 77 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.69 $Y=1.565 $X2=1.69
+ $Y2=1.815
r231 8 10 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.69 $Y=1.565 $X2=1.69
+ $Y2=1.08
r232 4 76 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.05 $Y=2.065 $X2=1.05
+ $Y2=1.815
r233 4 6 96.3053 $w=5e-07 $l=9e-07 $layer=POLY_cond $X=1.05 $Y=2.065 $X2=1.05
+ $Y2=2.965
r234 1 75 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.91 $Y=1.565 $X2=0.91
+ $Y2=1.815
r235 1 3 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.91 $Y=1.565 $X2=0.91
+ $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_8%VPWR 1 2 3 4 5 16 17 18 20 22 26 28 30 32 35
+ 45 57 69 81 87
r96 85 87 0.153562 $w=3.7e-07 $l=4e-07 $layer=MET1_cond $X=6.54 $Y=3.63 $X2=6.94
+ $Y2=3.63
r97 84 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.94 $Y=3.56
+ $X2=6.94 $Y2=3.56
r98 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.54 $Y=3.56
+ $X2=6.54 $Y2=3.56
r99 81 84 21.1937 $w=5.68e-07 $l=1.01e-06 $layer=LI1_cond $X=6.74 $Y=2.55
+ $X2=6.74 $Y2=3.56
r100 77 85 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=5.7 $Y=3.63
+ $X2=6.54 $Y2=3.63
r101 75 77 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=5.34 $Y=3.63
+ $X2=5.7 $Y2=3.63
r102 73 75 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=4.98 $Y=3.63
+ $X2=5.34 $Y2=3.63
r103 72 79 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=5.34 $Y=3.56
+ $X2=5.34 $Y2=3.57
r104 72 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.7 $Y=3.56 $X2=5.7
+ $Y2=3.56
r105 72 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.34 $Y=3.56
+ $X2=5.34 $Y2=3.56
r106 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.98 $Y=3.56
+ $X2=4.98 $Y2=3.56
r107 69 72 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=5.34 $Y=2.55
+ $X2=5.34 $Y2=3.56
r108 65 73 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=4.14 $Y=3.63
+ $X2=4.98 $Y2=3.63
r109 63 65 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=3.78 $Y=3.63
+ $X2=4.14 $Y2=3.63
r110 60 67 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=3.78 $Y=3.56
+ $X2=3.78 $Y2=3.57
r111 60 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.14 $Y=3.56
+ $X2=4.14 $Y2=3.56
r112 60 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.78 $Y=3.56
+ $X2=3.78 $Y2=3.56
r113 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.42 $Y=3.56
+ $X2=3.42 $Y2=3.56
r114 57 60 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=3.78 $Y=2.55
+ $X2=3.78 $Y2=3.56
r115 53 61 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=2.58 $Y=3.63
+ $X2=3.42 $Y2=3.63
r116 51 53 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=2.22 $Y=3.63
+ $X2=2.58 $Y2=3.63
r117 49 51 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=1.86 $Y=3.63
+ $X2=2.22 $Y2=3.63
r118 48 55 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=2.22 $Y=3.56
+ $X2=2.22 $Y2=3.57
r119 48 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.58 $Y=3.56
+ $X2=2.58 $Y2=3.56
r120 48 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.22 $Y=3.56
+ $X2=2.22 $Y2=3.56
r121 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.86 $Y=3.56
+ $X2=1.86 $Y2=3.56
r122 45 48 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=2.22 $Y=2.55
+ $X2=2.22 $Y2=3.56
r123 41 49 0.368549 $w=3.7e-07 $l=9.6e-07 $layer=MET1_cond $X=0.9 $Y=3.63
+ $X2=1.86 $Y2=3.63
r124 39 41 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=0.54 $Y=3.63
+ $X2=0.9 $Y2=3.63
r125 38 43 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=0.54 $Y=3.56
+ $X2=0.54 $Y2=3.57
r126 38 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.9 $Y=3.56 $X2=0.9
+ $Y2=3.56
r127 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.54 $Y=3.56
+ $X2=0.54 $Y2=3.56
r128 35 38 13.8449 $w=8.88e-07 $l=1.01e-06 $layer=LI1_cond $X=0.54 $Y=2.55
+ $X2=0.54 $Y2=3.56
r129 32 63 0.069103 $w=3.7e-07 $l=1.8e-07 $layer=MET1_cond $X=3.6 $Y=3.63
+ $X2=3.78 $Y2=3.63
r130 32 61 0.069103 $w=3.7e-07 $l=1.8e-07 $layer=MET1_cond $X=3.6 $Y=3.63
+ $X2=3.42 $Y2=3.63
r131 31 84 1.36395 $w=5.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.74 $Y=3.625
+ $X2=6.74 $Y2=3.56
r132 29 79 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=5.34 $Y=3.625
+ $X2=5.34 $Y2=3.57
r133 29 30 3.33002 $w=8.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=3.625
+ $X2=5.34 $Y2=3.71
r134 27 67 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=3.78 $Y=3.625
+ $X2=3.78 $Y2=3.57
r135 27 28 3.33002 $w=8.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=3.625
+ $X2=3.78 $Y2=3.71
r136 25 55 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=2.22 $Y=3.625
+ $X2=2.22 $Y2=3.57
r137 25 26 3.33002 $w=8.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=3.625
+ $X2=2.22 $Y2=3.71
r138 24 43 0.753933 $w=8.88e-07 $l=5.5e-08 $layer=LI1_cond $X=0.54 $Y=3.625
+ $X2=0.54 $Y2=3.57
r139 23 30 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=5.785 $Y=3.71
+ $X2=5.34 $Y2=3.71
r140 22 31 9.80657 $w=1.7e-07 $l=3.24731e-07 $layer=LI1_cond $X=6.455 $Y=3.71
+ $X2=6.74 $Y2=3.625
r141 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.455 $Y=3.71
+ $X2=5.785 $Y2=3.71
r142 21 28 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=4.225 $Y=3.71
+ $X2=3.78 $Y2=3.71
r143 20 30 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=4.895 $Y=3.71
+ $X2=5.34 $Y2=3.71
r144 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.895 $Y=3.71
+ $X2=4.225 $Y2=3.71
r145 19 26 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=2.665 $Y=3.71
+ $X2=2.22 $Y2=3.71
r146 18 28 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=3.335 $Y=3.71
+ $X2=3.78 $Y2=3.71
r147 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.335 $Y=3.71
+ $X2=2.665 $Y2=3.71
r148 17 24 12.0932 $w=1.7e-07 $l=4.85644e-07 $layer=LI1_cond $X=0.985 $Y=3.71
+ $X2=0.54 $Y2=3.625
r149 16 26 15.4217 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=1.775 $Y=3.71
+ $X2=2.22 $Y2=3.71
r150 16 17 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.775 $Y=3.71
+ $X2=0.985 $Y2=3.71
r151 5 84 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=6.76
+ $Y=2.215 $X2=6.9 $Y2=3.57
r152 5 81 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=6.76
+ $Y=2.215 $X2=6.9 $Y2=2.55
r153 4 79 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=5.2
+ $Y=2.215 $X2=5.34 $Y2=3.57
r154 4 69 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=5.2
+ $Y=2.215 $X2=5.34 $Y2=2.55
r155 3 67 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=3.64
+ $Y=2.215 $X2=3.78 $Y2=3.57
r156 3 57 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=3.64
+ $Y=2.215 $X2=3.78 $Y2=2.55
r157 2 55 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=2.08
+ $Y=2.215 $X2=2.22 $Y2=3.57
r158 2 45 300 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=2 $X=2.08
+ $Y=2.215 $X2=2.22 $Y2=2.55
r159 1 43 300 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_PDIFF $count=2 $X=0.535
+ $Y=2.215 $X2=0.66 $Y2=3.57
r160 1 35 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=0.535
+ $Y=2.215 $X2=0.66 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_8%Y 1 2 3 4 5 6 7 8 27 31 35 36 37 38 41 45 49
+ 51 55 59 63 65 69 73 75 78 79 80 81 82 83 84 93
r121 93 94 0.0942813 $w=6.47e-07 $l=5e-09 $layer=LI1_cond $X=6.24 $Y=1.31
+ $X2=6.24 $Y2=1.315
r122 84 93 7.25966 $w=6.47e-07 $l=3.85e-07 $layer=LI1_cond $X=6.24 $Y=0.925
+ $X2=6.24 $Y2=1.31
r123 84 89 0.565688 $w=6.47e-07 $l=3e-08 $layer=LI1_cond $X=6.24 $Y=0.925
+ $X2=6.24 $Y2=0.895
r124 77 78 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=7.025 $Y=1.395
+ $X2=7.025 $Y2=2.035
r125 76 93 8.80565 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=6.565 $Y=1.31
+ $X2=6.24 $Y2=1.31
r126 75 77 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.94 $Y=1.31
+ $X2=7.025 $Y2=1.395
r127 75 76 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.94 $Y=1.31
+ $X2=6.565 $Y2=1.31
r128 74 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.285 $Y=2.12
+ $X2=6.12 $Y2=2.12
r129 73 78 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.94 $Y=2.12
+ $X2=7.025 $Y2=2.035
r130 73 74 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=6.94 $Y=2.12
+ $X2=6.285 $Y2=2.12
r131 69 71 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=6.12 $Y=2.34
+ $X2=6.12 $Y2=3.36
r132 67 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.12 $Y=2.205
+ $X2=6.12 $Y2=2.12
r133 67 69 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.12 $Y=2.205
+ $X2=6.12 $Y2=2.34
r134 66 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=2.12
+ $X2=4.56 $Y2=2.12
r135 65 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.955 $Y=2.12
+ $X2=6.12 $Y2=2.12
r136 65 66 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=5.955 $Y=2.12
+ $X2=4.725 $Y2=2.12
r137 64 81 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.525 $Y=1.315
+ $X2=4.42 $Y2=1.315
r138 63 94 8.80565 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=5.915 $Y=1.315
+ $X2=6.24 $Y2=1.315
r139 63 64 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=5.915 $Y=1.315
+ $X2=4.525 $Y2=1.315
r140 59 61 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=4.56 $Y=2.34
+ $X2=4.56 $Y2=3.36
r141 57 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=2.205
+ $X2=4.56 $Y2=2.12
r142 57 59 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=4.56 $Y=2.205
+ $X2=4.56 $Y2=2.34
r143 53 81 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=1.23
+ $X2=4.42 $Y2=1.315
r144 53 55 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=4.42 $Y=1.23
+ $X2=4.42 $Y2=0.895
r145 52 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=2.12 $X2=3
+ $Y2=2.12
r146 51 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=2.12
+ $X2=4.56 $Y2=2.12
r147 51 52 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=4.395 $Y=2.12
+ $X2=3.165 $Y2=2.12
r148 50 79 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.965 $Y=1.315
+ $X2=2.86 $Y2=1.315
r149 49 81 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.315 $Y=1.315
+ $X2=4.42 $Y2=1.315
r150 49 50 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=4.315 $Y=1.315
+ $X2=2.965 $Y2=1.315
r151 45 47 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3 $Y=2.34 $X2=3
+ $Y2=3.36
r152 43 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=2.205 $X2=3
+ $Y2=2.12
r153 43 45 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3 $Y=2.205 $X2=3
+ $Y2=2.34
r154 39 79 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=1.23
+ $X2=2.86 $Y2=1.315
r155 39 41 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=2.86 $Y=1.23
+ $X2=2.86 $Y2=0.895
r156 37 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=2.12 $X2=3
+ $Y2=2.12
r157 37 38 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=2.835 $Y=2.12
+ $X2=1.605 $Y2=2.12
r158 35 79 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.755 $Y=1.315
+ $X2=2.86 $Y2=1.315
r159 35 36 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=2.755 $Y=1.315
+ $X2=1.405 $Y2=1.315
r160 31 33 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=1.44 $Y=2.34
+ $X2=1.44 $Y2=3.36
r161 29 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.44 $Y=2.205
+ $X2=1.605 $Y2=2.12
r162 29 31 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.44 $Y=2.205
+ $X2=1.44 $Y2=2.34
r163 25 36 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.3 $Y=1.23
+ $X2=1.405 $Y2=1.315
r164 25 27 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=1.3 $Y=1.23
+ $X2=1.3 $Y2=0.895
r165 8 71 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=5.98
+ $Y=2.215 $X2=6.12 $Y2=3.36
r166 8 69 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=5.98
+ $Y=2.215 $X2=6.12 $Y2=2.34
r167 7 61 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=4.42
+ $Y=2.215 $X2=4.56 $Y2=3.36
r168 7 59 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.42
+ $Y=2.215 $X2=4.56 $Y2=2.34
r169 6 47 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=2.86
+ $Y=2.215 $X2=3 $Y2=3.36
r170 6 45 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.86
+ $Y=2.215 $X2=3 $Y2=2.34
r171 5 33 300 $w=1.7e-07 $l=1.21298e-06 $layer=licon1_PDIFF $count=2 $X=1.3
+ $Y=2.215 $X2=1.44 $Y2=3.36
r172 5 31 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.3
+ $Y=2.215 $X2=1.44 $Y2=2.34
r173 4 89 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=5.98
+ $Y=0.705 $X2=6.12 $Y2=0.895
r174 3 55 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=4.28
+ $Y=0.705 $X2=4.42 $Y2=0.895
r175 2 41 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=2.72
+ $Y=0.705 $X2=2.86 $Y2=0.895
r176 1 27 91 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=2 $X=1.16
+ $Y=0.705 $X2=1.3 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_8%VGND 1 2 3 4 5 18 20 22 34 43 54 60 63 67 71
+ 77 80
r72 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.02 $Y=0.465
+ $X2=7.02 $Y2=0.465
r73 75 77 10.5793 $w=6.63e-07 $l=1.65e-07 $layer=LI1_cond $X=5.58 $Y=0.712
+ $X2=5.745 $Y2=0.712
r74 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.58 $Y=0.465
+ $X2=5.58 $Y2=0.465
r75 73 75 6.83473 $w=6.63e-07 $l=3.8e-07 $layer=LI1_cond $X=5.2 $Y=0.712
+ $X2=5.58 $Y2=0.712
r76 70 76 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=4.86 $Y=0.44
+ $X2=5.58 $Y2=0.44
r77 69 73 6.11529 $w=6.63e-07 $l=3.4e-07 $layer=LI1_cond $X=4.86 $Y=0.712
+ $X2=5.2 $Y2=0.712
r78 69 71 10.5793 $w=6.63e-07 $l=1.65e-07 $layer=LI1_cond $X=4.86 $Y=0.712
+ $X2=4.695 $Y2=0.712
r79 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.86 $Y=0.465
+ $X2=4.86 $Y2=0.465
r80 65 67 14.1765 $w=6.63e-07 $l=3.65e-07 $layer=LI1_cond $X=3.78 $Y=0.712
+ $X2=4.145 $Y2=0.712
r81 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.78 $Y=0.465
+ $X2=3.78 $Y2=0.465
r82 62 65 2.51806 $w=6.63e-07 $l=1.4e-07 $layer=LI1_cond $X=3.64 $Y=0.712
+ $X2=3.78 $Y2=0.712
r83 62 63 16.6946 $w=6.63e-07 $l=5.05e-07 $layer=LI1_cond $X=3.64 $Y=0.712
+ $X2=3.135 $Y2=0.712
r84 58 60 12.0182 $w=6.63e-07 $l=2.45e-07 $layer=LI1_cond $X=2.34 $Y=0.712
+ $X2=2.585 $Y2=0.712
r85 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.34 $Y=0.465
+ $X2=2.34 $Y2=0.465
r86 56 58 4.6764 $w=6.63e-07 $l=2.6e-07 $layer=LI1_cond $X=2.08 $Y=0.712
+ $X2=2.34 $Y2=0.712
r87 53 59 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.62 $Y=0.44
+ $X2=2.34 $Y2=0.44
r88 52 56 8.27363 $w=6.63e-07 $l=4.6e-07 $layer=LI1_cond $X=1.62 $Y=0.712
+ $X2=2.08 $Y2=0.712
r89 52 54 8.42098 $w=6.63e-07 $l=4.5e-08 $layer=LI1_cond $X=1.62 $Y=0.712
+ $X2=1.575 $Y2=0.712
r90 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.62 $Y=0.465
+ $X2=1.62 $Y2=0.465
r91 47 53 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.9 $Y=0.44
+ $X2=1.62 $Y2=0.44
r92 44 47 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.18 $Y=0.44
+ $X2=0.9 $Y2=0.44
r93 43 49 6.51124 $w=8.88e-07 $l=4.75e-07 $layer=LI1_cond $X=0.54 $Y=0.465
+ $X2=0.54 $Y2=0.94
r94 43 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.9 $Y=0.465
+ $X2=0.9 $Y2=0.465
r95 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.18 $Y=0.465
+ $X2=0.18 $Y2=0.465
r96 41 80 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=6.66 $Y=0.44
+ $X2=7.02 $Y2=0.44
r97 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.66 $Y=0.465
+ $X2=6.66 $Y2=0.465
r98 38 41 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.94 $Y=0.44
+ $X2=6.66 $Y2=0.44
r99 38 76 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=5.94 $Y=0.44
+ $X2=5.58 $Y2=0.44
r100 37 40 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=5.94 $Y=0.465
+ $X2=6.66 $Y2=0.465
r101 37 77 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.94 $Y=0.465
+ $X2=5.745 $Y2=0.465
r102 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.94 $Y=0.465
+ $X2=5.94 $Y2=0.465
r103 34 79 5.55669 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.735 $Y=0.465
+ $X2=6.92 $Y2=0.465
r104 34 40 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.735 $Y=0.465
+ $X2=6.66 $Y2=0.465
r105 33 70 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=4.5 $Y=0.44
+ $X2=4.86 $Y2=0.44
r106 33 66 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=4.5 $Y=0.44
+ $X2=3.78 $Y2=0.44
r107 32 71 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.5 $Y=0.465
+ $X2=4.695 $Y2=0.465
r108 32 67 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.5 $Y=0.465
+ $X2=4.145 $Y2=0.465
r109 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.5 $Y=0.465
+ $X2=4.5 $Y2=0.465
r110 28 59 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.06 $Y=0.44
+ $X2=2.34 $Y2=0.44
r111 27 63 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.06 $Y=0.465
+ $X2=3.135 $Y2=0.465
r112 27 60 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.06 $Y=0.465
+ $X2=2.585 $Y2=0.465
r113 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.06 $Y=0.465
+ $X2=3.06 $Y2=0.465
r114 22 66 0.069103 $w=3.7e-07 $l=1.8e-07 $layer=MET1_cond $X=3.6 $Y=0.44
+ $X2=3.78 $Y2=0.44
r115 22 28 0.207309 $w=3.7e-07 $l=5.4e-07 $layer=MET1_cond $X=3.6 $Y=0.44
+ $X2=3.06 $Y2=0.44
r116 18 79 2.55307 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=0.55
+ $X2=6.92 $Y2=0.465
r117 18 20 12.1474 $w=3.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.92 $Y=0.55
+ $X2=6.92 $Y2=0.94
r118 17 43 10.9281 $w=1.7e-07 $l=4.45e-07 $layer=LI1_cond $X=0.985 $Y=0.465
+ $X2=0.54 $Y2=0.465
r119 17 54 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.985 $Y=0.465
+ $X2=1.575 $Y2=0.465
r120 5 20 182 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_NDIFF $count=1 $X=6.76
+ $Y=0.705 $X2=6.91 $Y2=0.94
r121 4 73 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=5.06
+ $Y=0.705 $X2=5.2 $Y2=0.94
r122 3 62 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.5
+ $Y=0.705 $X2=3.64 $Y2=0.94
r123 2 56 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.94
+ $Y=0.705 $X2=2.08 $Y2=0.94
r124 1 49 91 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=2 $X=0.395
+ $Y=0.705 $X2=0.52 $Y2=0.94
.ends

