# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hvl__sdfrbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  20.16000 BY  4.070000 ;
  SYMMETRY X Y R90 ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.625000 2.330000 2.135000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.700000 0.685000 20.040000 3.755000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.435000 0.515000 17.835000 3.570000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAPARTIALMETALSIDEAREA  7.210000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685000 1.625000 11.245000 2.135000 ;
    END
    PORT
      LAYER li1 ;
        RECT 15.005000 1.425000 15.685000 2.120000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.235000 1.295000 5.635000 2.150000 ;
    END
    PORT
      LAYER met1 ;
        RECT  5.375000 1.920000  5.665000 1.965000 ;
        RECT  5.375000 1.965000 15.265000 2.105000 ;
        RECT  5.375000 2.105000  5.665000 2.150000 ;
        RECT 10.655000 1.920000 10.945000 1.965000 ;
        RECT 10.655000 2.105000 10.945000 2.150000 ;
        RECT 14.975000 1.920000 15.265000 1.965000 ;
        RECT 14.975000 2.105000 15.265000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.710000 1.975000 4.705000 2.155000 ;
        RECT 3.710000 2.155000 4.040000 2.480000 ;
        RECT 4.375000 1.295000 4.705000 1.975000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.655000 1.295000 0.985000 1.965000 ;
        RECT 0.815000 0.265000 1.685000 0.435000 ;
        RECT 0.815000 0.435000 0.985000 1.295000 ;
        RECT 1.515000 0.435000 1.685000 1.275000 ;
        RECT 1.515000 1.275000 4.195000 1.445000 ;
        RECT 3.485000 1.445000 4.195000 1.795000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.870000 1.850000 6.200000 2.520000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.365000 0.635000 1.115000 ;
    END
    PORT
      LAYER li1 ;
        RECT 10.770000 0.365000 11.805000 0.745000 ;
    END
    PORT
      LAYER li1 ;
        RECT 14.450000 0.365000 15.400000 0.895000 ;
    END
    PORT
      LAYER li1 ;
        RECT 16.725000 0.365000 17.255000 1.305000 ;
    END
    PORT
      LAYER li1 ;
        RECT 18.565000 0.365000 19.515000 1.475000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.275000 0.365000 6.225000 0.995000 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.870000 0.365000 7.720000 0.915000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 20.160000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 20.160000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 20.160000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 20.160000 4.155000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 20.160000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.090000 3.205000 0.985000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 11.955000 3.015000 12.545000 3.735000 ;
    END
    PORT
      LAYER li1 ;
        RECT 14.800000 2.675000 15.720000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 16.330000 2.185000 17.255000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 18.535000 2.175000 19.485000 3.755000 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.545000 3.365000 3.495000 3.735000 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.085000 3.365000 5.975000 3.755000 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.205000 2.205000 7.375000 3.705000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.925000 3.255000 10.875000 3.755000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 20.160000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  1.165000 0.615000  1.335000 2.315000 ;
      RECT  1.165000 2.315000  3.440000 2.485000 ;
      RECT  1.165000 2.485000  1.335000 3.205000 ;
      RECT  1.165000 3.205000  1.415000 3.705000 ;
      RECT  1.515000 2.665000  3.040000 2.835000 ;
      RECT  1.515000 2.835000  1.765000 2.995000 ;
      RECT  1.675000 3.235000  2.115000 3.735000 ;
      RECT  1.865000 0.265000  5.095000 0.435000 ;
      RECT  1.865000 0.435000  2.115000 0.995000 ;
      RECT  1.945000 3.015000  6.325000 3.185000 ;
      RECT  1.945000 3.185000  2.115000 3.235000 ;
      RECT  2.730000 1.625000  3.060000 2.315000 ;
      RECT  3.270000 2.485000  3.440000 2.665000 ;
      RECT  3.270000 2.665000  4.680000 2.835000 ;
      RECT  3.275000 0.615000  3.605000 0.925000 ;
      RECT  3.275000 0.925000  5.055000 1.095000 ;
      RECT  4.350000 2.325000  4.680000 2.665000 ;
      RECT  4.655000 3.185000  4.905000 3.735000 ;
      RECT  4.765000 0.435000  5.095000 0.755000 ;
      RECT  4.885000 1.095000  5.055000 3.015000 ;
      RECT  6.155000 3.185000  6.325000 3.635000 ;
      RECT  6.155000 3.635000  7.025000 3.805000 ;
      RECT  6.505000 0.495000  6.675000 1.505000 ;
      RECT  6.505000 1.505000  7.695000 1.675000 ;
      RECT  6.505000 1.675000  6.675000 3.455000 ;
      RECT  6.855000 1.855000  7.725000 2.025000 ;
      RECT  6.855000 2.025000  7.025000 3.635000 ;
      RECT  7.365000 1.345000  7.695000 1.505000 ;
      RECT  7.555000 2.025000  7.725000 3.255000 ;
      RECT  7.555000 3.255000  8.955000 3.425000 ;
      RECT  7.900000 0.265000  9.975000 0.435000 ;
      RECT  7.900000 0.435000  8.150000 0.995000 ;
      RECT  7.905000 0.995000  8.150000 2.225000 ;
      RECT  7.905000 2.225000  8.605000 3.015000 ;
      RECT  8.275000 3.425000  8.605000 3.755000 ;
      RECT  8.355000 3.015000  8.605000 3.075000 ;
      RECT  8.410000 0.615000  8.955000 0.995000 ;
      RECT  8.785000 0.995000  8.955000 3.255000 ;
      RECT  9.135000 0.615000  9.520000 0.995000 ;
      RECT  9.135000 0.995000  9.305000 2.905000 ;
      RECT  9.135000 2.905000 11.775000 3.075000 ;
      RECT  9.135000 3.075000  9.385000 3.755000 ;
      RECT  9.510000 2.005000  9.840000 2.315000 ;
      RECT  9.510000 2.315000 11.595000 2.485000 ;
      RECT  9.510000 2.485000  9.840000 2.675000 ;
      RECT  9.700000 0.435000  9.975000 0.925000 ;
      RECT  9.700000 0.925000 12.145000 1.095000 ;
      RECT  9.700000 1.095000  9.975000 1.755000 ;
      RECT 10.225000 1.275000 12.645000 1.445000 ;
      RECT 10.225000 1.445000 10.505000 1.945000 ;
      RECT 11.325000 2.665000 11.945000 2.835000 ;
      RECT 11.325000 2.835000 11.775000 2.905000 ;
      RECT 11.325000 3.075000 11.775000 3.735000 ;
      RECT 11.425000 1.875000 12.295000 2.045000 ;
      RECT 11.425000 2.045000 11.595000 2.315000 ;
      RECT 11.775000 2.225000 11.945000 2.665000 ;
      RECT 11.975000 0.265000 14.270000 0.435000 ;
      RECT 11.975000 0.435000 12.145000 0.925000 ;
      RECT 12.125000 2.045000 12.295000 2.175000 ;
      RECT 12.125000 2.175000 13.220000 2.345000 ;
      RECT 12.315000 0.615000 12.645000 1.275000 ;
      RECT 12.475000 1.445000 12.645000 1.825000 ;
      RECT 12.475000 1.825000 13.570000 1.995000 ;
      RECT 12.735000 2.525000 13.570000 2.695000 ;
      RECT 12.735000 2.695000 12.985000 3.755000 ;
      RECT 12.825000 0.435000 12.995000 1.475000 ;
      RECT 12.825000 1.475000 13.155000 1.645000 ;
      RECT 13.175000 0.615000 13.425000 1.125000 ;
      RECT 13.175000 1.125000 13.920000 1.295000 ;
      RECT 13.400000 1.995000 13.570000 2.525000 ;
      RECT 13.435000 2.875000 14.620000 3.045000 ;
      RECT 13.435000 3.045000 13.765000 3.755000 ;
      RECT 13.750000 1.295000 13.920000 2.875000 ;
      RECT 14.100000 0.435000 14.270000 2.555000 ;
      RECT 14.450000 1.075000 16.195000 1.245000 ;
      RECT 14.450000 1.245000 14.620000 2.875000 ;
      RECT 14.800000 2.300000 16.150000 2.495000 ;
      RECT 15.865000 1.245000 16.195000 1.655000 ;
      RECT 15.900000 2.495000 16.150000 3.175000 ;
      RECT 15.980000 1.835000 16.545000 2.005000 ;
      RECT 15.980000 2.005000 16.150000 2.300000 ;
      RECT 16.175000 0.515000 16.545000 0.895000 ;
      RECT 16.375000 0.895000 16.545000 1.835000 ;
      RECT 18.025000 0.685000 18.385000 1.655000 ;
      RECT 18.025000 1.655000 19.520000 1.985000 ;
      RECT 18.025000 1.985000 18.355000 2.985000 ;
    LAYER mcon ;
      RECT  0.095000  0.395000  0.265000 0.565000 ;
      RECT  0.095000  3.505000  0.265000 3.675000 ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.455000  0.395000  0.625000 0.565000 ;
      RECT  0.455000  3.505000  0.625000 3.675000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.815000  3.505000  0.985000 3.675000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.575000  3.505000  2.745000 3.675000 ;
      RECT  2.935000  3.505000  3.105000 3.675000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.295000  3.505000  3.465000 3.675000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.085000  3.505000  5.255000 3.675000 ;
      RECT  5.305000  0.395000  5.475000 0.565000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.950000  5.605000 2.120000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.445000  3.505000  5.615000 3.675000 ;
      RECT  5.665000  0.395000  5.835000 0.565000 ;
      RECT  5.805000  3.505000  5.975000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.025000  0.395000  6.195000 0.565000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  6.950000  0.395000  7.120000 0.565000 ;
      RECT  7.205000  3.505000  7.375000 3.675000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.470000  0.395000  7.640000 0.565000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.955000  3.505000 10.125000 3.675000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.315000  3.505000 10.485000 3.675000 ;
      RECT 10.675000  3.505000 10.845000 3.675000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.950000 10.885000 2.120000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.800000  0.395000 10.970000 0.565000 ;
      RECT 11.160000  0.395000 11.330000 0.565000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.520000  0.395000 11.690000 0.565000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 11.985000  3.505000 12.155000 3.675000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.345000  3.505000 12.515000 3.675000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.480000  0.395000 14.650000 0.565000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.815000  3.505000 14.985000 3.675000 ;
      RECT 14.840000  0.395000 15.010000 0.565000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  1.950000 15.205000 2.120000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.175000  3.505000 15.345000 3.675000 ;
      RECT 15.200000  0.395000 15.370000 0.565000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.535000  3.505000 15.705000 3.675000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.345000  3.505000 16.515000 3.675000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.705000  3.505000 16.875000 3.675000 ;
      RECT 16.725000  0.395000 16.895000 0.565000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 17.065000  3.505000 17.235000 3.675000 ;
      RECT 17.085000  0.395000 17.255000 0.565000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.985000 18.085000 4.155000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.985000 18.565000 4.155000 ;
      RECT 18.565000  3.505000 18.735000 3.675000 ;
      RECT 18.595000  0.395000 18.765000 0.565000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  3.985000 19.045000 4.155000 ;
      RECT 18.925000  3.505000 19.095000 3.675000 ;
      RECT 18.955000  0.395000 19.125000 0.565000 ;
      RECT 19.285000  3.505000 19.455000 3.675000 ;
      RECT 19.315000  0.395000 19.485000 0.565000 ;
      RECT 19.355000 -0.085000 19.525000 0.085000 ;
      RECT 19.355000  3.985000 19.525000 4.155000 ;
      RECT 19.835000 -0.085000 20.005000 0.085000 ;
      RECT 19.835000  3.985000 20.005000 4.155000 ;
  END
END sky130_fd_sc_hvl__sdfrbp_1
END LIBRARY
