* File: sky130_fd_sc_hvl__dfxbp_1.spice
* Created: Wed Sep  2 09:05:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__dfxbp_1.pex.spice"
.subckt sky130_fd_sc_hvl__dfxbp_1  VNB VPB CLK D VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1025 N_VGND_M1025_d N_CLK_M1025_g N_A_30_112#_M1025_s N_VNB_M1025_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1004 N_A_339_112#_M1004_d N_A_30_112#_M1004_g N_VGND_M1025_d N_VNB_M1025_b NHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1013 N_A_709_111#_M1013_d N_D_M1013_g N_VGND_M1013_s N_VNB_M1025_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1533 PD=0.7 PS=1.57 NRD=0 NRS=21.7056 M=1 R=0.84
+ SA=250000 SB=250006 A=0.21 P=1.84 MULT=1
MM1026 N_A_865_111#_M1026_d N_A_30_112#_M1026_g N_A_709_111#_M1013_d
+ N_VNB_M1025_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0
+ M=1 R=0.84 SA=250001 SB=250006 A=0.21 P=1.84 MULT=1
MM1018 A_1021_111# N_A_339_112#_M1018_g N_A_865_111#_M1026_d N_VNB_M1025_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1021 N_VGND_M1021_d N_A_1063_85#_M1021_g A_1021_111# N_VNB_M1025_b NHV L=0.5
+ W=0.42 AD=0.0879308 AS=0.0441 PD=0.807692 PS=0.63 NRD=25.7754 NRS=13.566 M=1
+ R=0.84 SA=250002 SB=250004 A=0.21 P=1.84 MULT=1
MM1023 N_A_1063_85#_M1023_d N_A_865_111#_M1023_g N_VGND_M1021_d N_VNB_M1025_b
+ NHV L=0.5 W=0.75 AD=0.157019 AS=0.157019 PD=1.44231 PS=1.44231 NRD=0 NRS=0 M=1
+ R=1.5 SA=250002 SB=250002 A=0.375 P=2.5 MULT=1
MM1024 N_A_1494_539#_M1024_d N_A_339_112#_M1024_g N_A_1063_85#_M1023_d
+ N_VNB_M1025_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.0879308 PD=0.7 PS=0.807692 NRD=0
+ NRS=25.7754 M=1 R=0.84 SA=250004 SB=250002 A=0.21 P=1.84 MULT=1
MM1007 A_1669_111# N_A_30_112#_M1007_g N_A_1494_539#_M1024_d N_VNB_M1025_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250005 SB=250002 A=0.21 P=1.84 MULT=1
MM1016 N_VGND_M1016_d N_A_1711_85#_M1016_g A_1669_111# N_VNB_M1025_b NHV L=0.5
+ W=0.42 AD=0.0879308 AS=0.0441 PD=0.807692 PS=0.63 NRD=25.7754 NRS=13.566 M=1
+ R=0.84 SA=250006 SB=250001 A=0.21 P=1.84 MULT=1
MM1009 N_A_1711_85#_M1009_d N_A_1494_539#_M1009_g N_VGND_M1016_d N_VNB_M1025_b
+ NHV L=0.5 W=0.75 AD=0.19875 AS=0.157019 PD=2.03 PS=1.44231 NRD=0 NRS=0 M=1
+ R=1.5 SA=250004 SB=250000 A=0.375 P=2.5 MULT=1
MM1010 N_VGND_M1010_d N_A_1711_85#_M1010_g N_Q_M1010_s N_VNB_M1025_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.19875 PD=2.07 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1014 N_VGND_M1014_d N_A_1711_85#_M1014_g N_A_2365_443#_M1014_s N_VNB_M1025_b
+ NHV L=0.5 W=0.42 AD=0.0933154 AS=0.1113 PD=0.822051 PS=1.37 NRD=31.2132 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1027 N_Q_N_M1027_d N_A_2365_443#_M1027_g N_VGND_M1014_d N_VNB_M1025_b NHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.166635 PD=2.03 PS=1.46795 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1012 N_VPWR_M1012_d N_CLK_M1012_g N_A_30_112#_M1012_s N_VPB_M1012_b PHV L=0.5
+ W=0.75 AD=0.105 AS=0.21375 PD=1.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1022 N_A_339_112#_M1022_d N_A_30_112#_M1022_g N_VPWR_M1012_d N_VPB_M1012_b PHV
+ L=0.5 W=0.75 AD=0.21375 AS=0.105 PD=2.07 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1006 N_A_709_111#_M1006_d N_D_M1006_g N_VPWR_M1006_s N_VPB_M1012_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250006 A=0.21 P=1.84 MULT=1
MM1019 N_A_865_111#_M1019_d N_A_339_112#_M1019_g N_A_709_111#_M1006_d
+ N_VPB_M1012_b PHV L=0.5 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0
+ M=1 R=0.84 SA=250001 SB=250006 A=0.21 P=1.84 MULT=1
MM1011 A_1021_539# N_A_30_112#_M1011_g N_A_865_111#_M1019_d N_VPB_M1012_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1015 N_VPWR_M1015_d N_A_1063_85#_M1015_g A_1021_539# N_VPB_M1012_b PHV L=0.5
+ W=0.42 AD=0.0920451 AS=0.0441 PD=0.81338 PS=0.63 NRD=45.458 NRS=22.729 M=1
+ R=0.84 SA=250002 SB=250004 A=0.21 P=1.84 MULT=1
MM1017 N_A_1063_85#_M1017_d N_A_865_111#_M1017_g N_VPWR_M1015_d N_VPB_M1012_b
+ PHV L=0.5 W=1 AD=0.14 AS=0.219155 PD=1.28 PS=1.93662 NRD=0 NRS=0 M=1 R=2
+ SA=250001 SB=250002 A=0.5 P=3 MULT=1
MM1000 N_A_1494_539#_M1000_d N_A_30_112#_M1000_g N_A_1063_85#_M1017_d
+ N_VPB_M1012_b PHV L=0.5 W=1 AD=0.219155 AS=0.14 PD=1.93662 PS=1.28 NRD=0 NRS=0
+ M=1 R=2 SA=250002 SB=250001 A=0.5 P=3 MULT=1
MM1002 A_1669_539# N_A_339_112#_M1002_g N_A_1494_539#_M1000_d N_VPB_M1012_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0920451 PD=0.63 PS=0.81338 NRD=22.729 NRS=43.1851
+ M=1 R=0.84 SA=250005 SB=250002 A=0.21 P=1.84 MULT=1
MM1008 N_VPWR_M1008_d N_A_1711_85#_M1008_g A_1669_539# N_VPB_M1012_b PHV L=0.5
+ W=0.42 AD=0.0920451 AS=0.0441 PD=0.81338 PS=0.63 NRD=43.1851 NRS=22.729 M=1
+ R=0.84 SA=250006 SB=250001 A=0.21 P=1.84 MULT=1
MM1003 N_A_1711_85#_M1003_d N_A_1494_539#_M1003_g N_VPWR_M1008_d N_VPB_M1012_b
+ PHV L=0.5 W=1 AD=0.265 AS=0.219155 PD=2.53 PS=1.93662 NRD=0 NRS=0 M=1 R=2
+ SA=250003 SB=250000 A=0.5 P=3 MULT=1
MM1001 N_VPWR_M1001_d N_A_1711_85#_M1001_g N_Q_M1001_s N_VPB_M1012_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.3975 PD=3.53 PS=3.53 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
MM1005 N_VPWR_M1005_d N_A_1711_85#_M1005_g N_A_2365_443#_M1005_s N_VPB_M1012_b
+ PHV L=0.5 W=0.75 AD=0.17 AS=0.19875 PD=1.26333 PS=2.03 NRD=29.2803 NRS=0 M=1
+ R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1020 N_Q_N_M1020_d N_A_2365_443#_M1020_g N_VPWR_M1005_d N_VPB_M1012_b PHV
+ L=0.5 W=1.5 AD=0.4275 AS=0.34 PD=3.57 PS=2.52667 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
DX28_noxref N_VNB_M1025_b N_VPB_M1012_b NWDIODE A=37.908 P=34.36
*
.include "sky130_fd_sc_hvl__dfxbp_1.pxi.spice"
*
.ends
*
*
