# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__schmittbuf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__schmittbuf_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.170000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.015000 1.855000 3.305000 2.150000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.860000 0.515000 5.195000 3.715000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 5.280000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 5.280000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 5.280000 4.155000 ;
      LAYER mcon ;
        RECT 0.155000 3.985000 0.325000 4.155000 ;
        RECT 0.635000 3.985000 0.805000 4.155000 ;
        RECT 1.115000 3.985000 1.285000 4.155000 ;
        RECT 1.595000 3.985000 1.765000 4.155000 ;
        RECT 2.075000 3.985000 2.245000 4.155000 ;
        RECT 2.555000 3.985000 2.725000 4.155000 ;
        RECT 3.035000 3.985000 3.205000 4.155000 ;
        RECT 3.515000 3.985000 3.685000 4.155000 ;
        RECT 3.995000 3.985000 4.165000 4.155000 ;
        RECT 4.475000 3.985000 4.645000 4.155000 ;
        RECT 4.955000 3.985000 5.125000 4.155000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 5.280000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 1.340000 1.975000 ;
        RECT -0.330000 1.975000 5.610000 4.485000 ;
        RECT  3.885000 1.885000 5.610000 1.975000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 5.280000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 1.805000 0.530000 1.975000 ;
      RECT 0.085000 1.975000 0.255000 3.485000 ;
      RECT 0.085000 3.485000 1.030000 3.655000 ;
      RECT 0.280000 1.090000 0.530000 1.805000 ;
      RECT 0.430000 2.165000 0.875000 2.335000 ;
      RECT 0.430000 2.335000 0.680000 3.085000 ;
      RECT 0.705000 0.570000 2.010000 0.795000 ;
      RECT 0.705000 0.795000 0.875000 2.165000 ;
      RECT 0.740000 3.405000 1.030000 3.485000 ;
      RECT 0.740000 3.655000 1.030000 3.735000 ;
      RECT 1.045000 1.655000 4.690000 1.685000 ;
      RECT 1.045000 1.685000 1.835000 1.985000 ;
      RECT 1.060000 0.975000 2.720000 1.145000 ;
      RECT 1.060000 1.145000 1.390000 1.410000 ;
      RECT 1.200000 2.295000 1.460000 3.235000 ;
      RECT 1.200000 3.235000 2.790000 3.405000 ;
      RECT 1.600000 1.315000 1.940000 1.505000 ;
      RECT 1.600000 1.505000 4.210000 1.645000 ;
      RECT 1.600000 1.645000 4.690000 1.655000 ;
      RECT 1.655000 1.985000 1.835000 2.330000 ;
      RECT 1.655000 2.330000 2.010000 3.065000 ;
      RECT 2.390000 1.145000 2.720000 1.335000 ;
      RECT 2.460000 2.320000 2.790000 3.235000 ;
      RECT 3.120000 0.375000 4.630000 1.285000 ;
      RECT 3.130000 3.405000 4.570000 3.735000 ;
      RECT 3.235000 2.320000 4.570000 3.405000 ;
      RECT 3.855000 1.685000 4.690000 2.055000 ;
    LAYER mcon ;
      RECT 3.210000 0.425000 3.380000 0.595000 ;
      RECT 3.225000 3.475000 3.395000 3.645000 ;
      RECT 3.570000 0.425000 3.740000 0.595000 ;
      RECT 3.585000 3.475000 3.755000 3.645000 ;
      RECT 3.945000 3.475000 4.115000 3.645000 ;
      RECT 3.980000 0.425000 4.150000 0.595000 ;
      RECT 4.305000 3.475000 4.475000 3.645000 ;
      RECT 4.410000 0.425000 4.580000 0.595000 ;
  END
END sky130_fd_sc_hvl__schmittbuf_1
END LIBRARY
