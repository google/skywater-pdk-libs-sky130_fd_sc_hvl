* NGSPICE file created from sky130_fd_sc_hvl__inv_4.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__inv_4 A VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB phv w=1.5e+06u l=500000u
+  ad=1.275e+12p pd=1.07e+07u as=8.4e+11p ps=7.12e+06u
M1001 Y A VGND VNB nhv w=750000u l=500000u
+  ad=4.2e+11p pd=4.12e+06u as=6.375e+11p ps=6.2e+06u
M1002 Y A VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A Y VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A Y VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A Y VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VGND VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends

