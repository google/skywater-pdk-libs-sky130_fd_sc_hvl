# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__o22ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__o22ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.805000 3.715000 2.120000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.250000 1.805000 2.755000 2.120000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.535000 0.550000 1.865000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.535000 1.595000 1.750000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.742500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.735000 0.615000 1.270000 1.355000 ;
        RECT 0.735000 1.355000 0.905000 1.930000 ;
        RECT 0.735000 1.930000 1.795000 2.100000 ;
        RECT 1.525000 2.100000 1.795000 2.175000 ;
        RECT 1.525000 2.175000 2.045000 3.260000 ;
        RECT 1.875000 3.260000 2.045000 3.755000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.840000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.840000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.840000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 4.170000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.840000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.985000 3.840000 4.155000 ;
      RECT 0.090000  2.280000 1.345000 3.755000 ;
      RECT 0.160000  0.265000 1.970000 0.435000 ;
      RECT 0.160000  0.435000 0.490000 1.355000 ;
      RECT 1.800000  0.435000 1.970000 1.455000 ;
      RECT 1.800000  1.455000 3.670000 1.625000 ;
      RECT 2.150000  0.365000 3.250000 1.275000 ;
      RECT 2.305000  2.300000 3.615000 3.755000 ;
      RECT 3.420000  0.525000 3.670000 1.455000 ;
    LAYER mcon ;
      RECT 0.095000  3.505000 0.265000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.455000  3.505000 0.625000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.815000  3.505000 0.985000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.175000  3.505000 1.345000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.200000  0.395000 2.370000 0.565000 ;
      RECT 2.335000  3.505000 2.505000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.560000  0.395000 2.730000 0.565000 ;
      RECT 2.695000  3.505000 2.865000 3.675000 ;
      RECT 2.920000  0.395000 3.090000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.055000  3.505000 3.225000 3.675000 ;
      RECT 3.415000  3.505000 3.585000 3.675000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
  END
END sky130_fd_sc_hvl__o22ai_1
END LIBRARY
