* File: sky130_fd_sc_hvl__lsbufhv2lv_1.pxi.spice
* Created: Fri Aug 28 09:36:50 2020
* 
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%VNB N_VNB_M1011_b VNB VNB N_VNB_c_24_p
+ N_VNB_c_5_p VNB VNB PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%VNB
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%VPB N_VPB_M1015_b N_VPB_X18_noxref_D1 VPB
+ N_VPB_c_85_p N_VPB_c_118_p N_VPB_c_71_n VPB
+ PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%VPB
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%LVPWR N_LVPWR_M1003_d N_LVPWR_M1001_d
+ N_LVPWR_M1003_b N_LVPWR_c_149_p N_LVPWR_c_128_n N_LVPWR_c_129_n LVPWR
+ N_LVPWR_c_126_n LVPWR PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%LVPWR
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A_30_1337# N_A_30_1337#_M1009_s
+ N_A_30_1337#_M1000_d N_A_30_1337#_c_214_n N_A_30_1337#_M1002_g
+ N_A_30_1337#_M1015_g N_A_30_1337#_c_196_n N_A_30_1337#_M1005_g
+ N_A_30_1337#_c_198_n N_A_30_1337#_c_199_n N_A_30_1337#_M1008_g
+ N_A_30_1337#_c_200_n N_A_30_1337#_M1012_g N_A_30_1337#_c_202_n
+ N_A_30_1337#_c_203_n N_A_30_1337#_M1014_g N_A_30_1337#_c_205_n
+ N_A_30_1337#_c_206_n N_A_30_1337#_c_207_n N_A_30_1337#_c_208_n
+ N_A_30_1337#_c_209_n N_A_30_1337#_c_210_n N_A_30_1337#_c_219_n
+ N_A_30_1337#_c_211_n N_A_30_1337#_c_212_n N_A_30_1337#_c_213_n
+ PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A_30_1337#
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A N_A_c_294_n N_A_M1000_g N_A_M1009_g
+ N_A_c_296_n N_A_c_297_n A A N_A_c_299_n PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A_30_207# N_A_30_207#_M1002_s
+ N_A_30_207#_M1015_d N_A_30_207#_M1004_g N_A_30_207#_c_322_n
+ N_A_30_207#_M1006_g N_A_30_207#_M1007_g N_A_30_207#_M1010_g
+ N_A_30_207#_c_326_n N_A_30_207#_c_327_n N_A_30_207#_c_328_n
+ N_A_30_207#_c_335_n N_A_30_207#_c_329_n N_A_30_207#_c_330_n
+ PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A_30_207#
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A_389_1337# N_A_389_1337#_M1005_d
+ N_A_389_1337#_M1008_d N_A_389_1337#_M1014_d N_A_389_1337#_M1013_d
+ N_A_389_1337#_M1001_g N_A_389_1337#_c_371_n N_A_389_1337#_c_372_n
+ N_A_389_1337#_c_373_n N_A_389_1337#_c_374_n N_A_389_1337#_c_375_n
+ N_A_389_1337#_c_376_n N_A_389_1337#_c_377_n N_A_389_1337#_c_393_n
+ N_A_389_1337#_c_378_n N_A_389_1337#_c_379_n N_A_389_1337#_c_380_n
+ PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A_389_1337#
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A_389_141# N_A_389_141#_M1004_s
+ N_A_389_141#_M1007_s N_A_389_141#_M1010_s N_A_389_141#_M1001_s
+ N_A_389_141#_c_445_n N_A_389_141#_c_446_n N_A_389_141#_c_447_n
+ N_A_389_141#_M1011_g N_A_389_141#_M1003_g N_A_389_141#_M1013_g
+ N_A_389_141#_c_450_n N_A_389_141#_c_451_n N_A_389_141#_c_452_n
+ N_A_389_141#_c_453_n N_A_389_141#_c_458_n N_A_389_141#_c_478_n
+ N_A_389_141#_c_454_n PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%A_389_141#
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%VPWR N_VPWR_M1015_s N_VPWR_M1000_s
+ N_VPWR_c_531_n N_VPWR_c_532_n VPWR VPWR N_VPWR_c_533_n N_VPWR_c_536_n VPWR
+ VPWR PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%VPWR
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%X N_X_M1011_s N_X_M1003_s X X X X X X
+ N_X_c_596_n PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%X
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%VGND N_VGND_M1002_d N_VGND_M1009_d
+ N_VGND_M1006_d N_VGND_M1007_d N_VGND_M1010_d N_VGND_M1008_s N_VGND_M1012_s
+ N_VGND_M1011_d VGND VGND N_VGND_c_611_n N_VGND_c_613_n N_VGND_c_615_n
+ N_VGND_c_617_n N_VGND_c_619_n N_VGND_c_621_n VGND VGND
+ PM_SKY130_FD_SC_HVL__LSBUFHV2LV_1%VGND
cc_1 N_VNB_M1011_b N_VPB_c_71_n 0.0458746f $X=-0.33 $Y=-0.265 $X2=7.92 $Y2=4.07
cc_2 N_VNB_M1011_b N_LVPWR_c_126_n 0.104679f $X=-0.33 $Y=-0.265 $X2=4.32
+ $Y2=4.068
cc_3 N_VNB_M1011_b N_A_30_1337#_M1002_g 0.0800155f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_4 N_VNB_M1011_b N_A_30_1337#_c_196_n 0.0441609f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_5 N_VNB_c_5_p N_A_30_1337#_c_196_n 0.00177683f $X=7.92 $Y=8.14 $X2=0 $Y2=0
cc_6 N_VNB_M1011_b N_A_30_1337#_c_198_n 0.0126934f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_7 N_VNB_M1011_b N_A_30_1337#_c_199_n 0.0347083f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_8 N_VNB_M1011_b N_A_30_1337#_c_200_n 0.0381344f $X=-0.33 $Y=-0.265 $X2=7.92
+ $Y2=4.07
cc_9 N_VNB_c_5_p N_A_30_1337#_c_200_n 0.00117942f $X=7.92 $Y=8.14 $X2=7.92
+ $Y2=4.07
cc_10 N_VNB_M1011_b N_A_30_1337#_c_202_n 0.0476552f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1011_b N_A_30_1337#_c_203_n 0.0442454f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_c_5_p N_A_30_1337#_c_203_n 0.00148776f $X=7.92 $Y=8.14 $X2=0 $Y2=0
cc_13 N_VNB_M1011_b N_A_30_1337#_c_205_n 0.0150462f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_M1011_b N_A_30_1337#_c_206_n 0.00795968f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_15 N_VNB_M1011_b N_A_30_1337#_c_207_n 0.00528668f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_16 N_VNB_M1011_b N_A_30_1337#_c_208_n 0.0013944f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_17 N_VNB_M1011_b N_A_30_1337#_c_209_n 0.0140388f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1011_b N_A_30_1337#_c_210_n 0.00634096f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_19 N_VNB_M1011_b N_A_30_1337#_c_211_n 0.0109898f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_20 N_VNB_M1011_b N_A_30_1337#_c_212_n 0.0496973f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_21 N_VNB_M1011_b N_A_30_1337#_c_213_n 0.0408601f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_22 N_VNB_M1011_b N_A_M1000_g 0.105199f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_23 N_VNB_M1011_b N_A_30_207#_M1004_g 0.0548441f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_24 N_VNB_c_24_p N_A_30_207#_M1004_g 0.00177683f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_25 N_VNB_M1011_b N_A_30_207#_c_322_n 0.0872215f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=3.955
cc_26 N_VNB_M1011_b N_A_30_207#_M1006_g 0.0532389f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_27 N_VNB_c_24_p N_A_30_207#_M1006_g 0.00133359f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_28 N_VNB_M1011_b N_A_30_207#_M1007_g 0.0731661f $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=4.07
cc_29 N_VNB_M1011_b N_A_30_207#_c_326_n 0.00528668f $X=-0.33 $Y=-0.265 $X2=7.92
+ $Y2=4.07
cc_30 N_VNB_M1011_b N_A_30_207#_c_327_n 6.51598e-19 $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=4.07
cc_31 N_VNB_M1011_b N_A_30_207#_c_328_n 0.0140388f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_32 N_VNB_M1011_b N_A_30_207#_c_329_n 0.00352805f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_33 N_VNB_M1011_b N_A_30_207#_c_330_n 0.0063605f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_M1011_b N_A_389_1337#_c_371_n 0.0191968f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_35 N_VNB_M1011_b N_A_389_1337#_c_372_n 0.0402584f $X=-0.33 $Y=-0.265 $X2=7.92
+ $Y2=4.07
cc_36 N_VNB_M1011_b N_A_389_1337#_c_373_n 0.00924932f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_37 N_VNB_M1011_b N_A_389_1337#_c_374_n 0.00489685f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_38 N_VNB_M1011_b N_A_389_1337#_c_375_n 0.0803719f $X=-0.33 $Y=-0.265 $X2=4.32
+ $Y2=4.068
cc_39 N_VNB_M1011_b N_A_389_1337#_c_376_n 0.0640209f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_M1011_b N_A_389_1337#_c_377_n 0.0735354f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_41 N_VNB_M1011_b N_A_389_1337#_c_378_n 0.0853837f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_42 N_VNB_M1011_b N_A_389_1337#_c_379_n 0.0144603f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_M1011_b N_A_389_1337#_c_380_n 0.018029f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_44 N_VNB_M1011_b N_A_389_141#_c_445_n 0.221183f $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=4.07
cc_45 N_VNB_M1011_b N_A_389_141#_c_446_n 0.0285954f $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=4.07
cc_46 N_VNB_M1011_b N_A_389_141#_c_447_n 0.037708f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_47 N_VNB_M1011_b N_A_389_141#_M1011_g 0.029045f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_c_24_p N_A_389_141#_M1011_g 5.48702e-19 $X=7.92 $Y=0 $X2=0 $Y2=0
cc_49 N_VNB_M1011_b N_A_389_141#_c_450_n 0.0448303f $X=-0.33 $Y=-0.265 $X2=7.92
+ $Y2=4.07
cc_50 N_VNB_M1011_b N_A_389_141#_c_451_n 0.0477688f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_51 N_VNB_M1011_b N_A_389_141#_c_452_n 0.0167391f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_52 N_VNB_M1011_b N_A_389_141#_c_453_n 0.00864539f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_53 N_VNB_M1011_b N_A_389_141#_c_454_n 0.0424485f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_54 N_VNB_M1011_b VPWR 0.0472087f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_55 N_VNB_M1011_b VPWR 0.127845f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_56 N_VNB_M1011_b N_X_c_596_n 0.0304474f $X=-0.33 $Y=-0.265 $X2=7.92 $Y2=4.07
cc_57 N_VNB_M1011_b N_VGND_c_611_n 0.0469969f $X=-0.33 $Y=-0.265 $X2=7.92
+ $Y2=4.07
cc_58 N_VNB_c_24_p N_VGND_c_611_n 0.00159492f $X=7.92 $Y=0 $X2=7.92 $Y2=4.07
cc_59 N_VNB_M1011_b N_VGND_c_613_n 0.0405793f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_60 N_VNB_c_5_p N_VGND_c_613_n 0.00159492f $X=7.92 $Y=8.14 $X2=0 $Y2=0
cc_61 N_VNB_M1011_b N_VGND_c_615_n 0.0472241f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_62 N_VNB_c_5_p N_VGND_c_615_n 0.00159492f $X=7.92 $Y=8.14 $X2=0 $Y2=0
cc_63 N_VNB_M1011_b N_VGND_c_617_n 0.0918106f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_64 N_VNB_c_24_p N_VGND_c_617_n 0.00159492f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_65 N_VNB_M1011_b N_VGND_c_619_n 0.0936208f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_66 N_VNB_c_24_p N_VGND_c_619_n 0.00159492f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_67 N_VNB_M1011_b N_VGND_c_621_n 0.334411f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_68 N_VNB_c_24_p N_VGND_c_621_n 0.873341f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_69 N_VNB_M1011_b VGND 0.361606f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_70 N_VNB_c_5_p VGND 0.873432f $X=7.92 $Y=8.14 $X2=0 $Y2=0
cc_71 N_VPB_c_71_n N_LVPWR_M1003_b 0.00876039f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_72 N_VPB_c_71_n N_LVPWR_c_128_n 0.0459925f $X=7.92 $Y=4.07 $X2=0.24 $Y2=0
cc_73 N_VPB_c_71_n N_LVPWR_c_129_n 0.0121537f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_74 N_VPB_M1015_b N_LVPWR_c_126_n 0.0260448f $X=-0.33 $Y=1.885 $X2=0.24
+ $Y2=8.14
cc_75 N_VPB_X18_noxref_D1 N_LVPWR_c_126_n 0.0692382f $X=7 $Y=1.885 $X2=0.24
+ $Y2=8.14
cc_76 N_VPB_M1015_b N_A_30_1337#_c_214_n 0.05835f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_77 N_VPB_M1015_b N_A_30_1337#_M1002_g 0.0435401f $X=-0.33 $Y=1.885 $X2=-0.33
+ $Y2=-0.265
cc_78 N_VPB_M1015_b N_A_30_1337#_c_208_n 8.1289e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_79 N_VPB_M1015_b N_A_30_1337#_c_209_n 0.00462706f $X=-0.33 $Y=1.885 $X2=0.24
+ $Y2=0
cc_80 N_VPB_M1015_b N_A_30_1337#_c_210_n 0.0108734f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_81 N_VPB_M1015_b N_A_30_1337#_c_219_n 0.0470269f $X=-0.33 $Y=1.885 $X2=4.32
+ $Y2=0.058
cc_82 N_VPB_M1015_b N_A_30_1337#_c_211_n 0.0161651f $X=-0.33 $Y=1.885 $X2=4.08
+ $Y2=8.14
cc_83 N_VPB_M1015_b N_A_30_1337#_c_212_n 0.0483344f $X=-0.33 $Y=1.885 $X2=4.32
+ $Y2=8.14
cc_84 N_VPB_c_85_p N_A_30_1337#_c_212_n 0.00283754f $X=0.72 $Y=4.07 $X2=4.32
+ $Y2=8.14
cc_85 N_VPB_c_71_n N_A_30_1337#_c_212_n 0.0230371f $X=7.92 $Y=4.07 $X2=4.32
+ $Y2=8.14
cc_86 N_VPB_M1015_b N_A_30_1337#_c_213_n 0.0127287f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_87 N_VPB_M1015_b N_A_c_294_n 0.0218752f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_88 N_VPB_M1015_b N_A_M1000_g 0.0427957f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_89 N_VPB_M1015_b N_A_c_296_n 0.0151278f $X=-0.33 $Y=1.885 $X2=-0.33
+ $Y2=-0.265
cc_90 N_VPB_M1015_b N_A_c_297_n 0.0308178f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_91 N_VPB_M1015_b A 0.0061586f $X=-0.33 $Y=1.885 $X2=0 $Y2=8.025
cc_92 N_VPB_M1015_b N_A_c_299_n 0.0455794f $X=-0.33 $Y=1.885 $X2=0.24 $Y2=0
cc_93 N_VPB_M1015_b N_A_30_207#_c_322_n 0.0148597f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_94 N_VPB_c_71_n N_A_30_207#_M1007_g 0.011079f $X=7.92 $Y=4.07 $X2=0.24 $Y2=0
cc_95 N_VPB_M1015_b N_A_30_207#_c_327_n 6.9836e-19 $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_96 N_VPB_M1015_b N_A_30_207#_c_328_n 0.00363373f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_97 N_VPB_M1015_b N_A_30_207#_c_335_n 0.00729926f $X=-0.33 $Y=1.885 $X2=0.24
+ $Y2=8.14
cc_98 N_VPB_M1015_b N_A_30_207#_c_329_n 0.00135355f $X=-0.33 $Y=1.885 $X2=7.92
+ $Y2=8.14
cc_99 N_VPB_M1015_b N_A_30_207#_c_330_n 0.00992608f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_100 N_VPB_c_71_n N_A_389_1337#_M1001_g 0.00401315f $X=7.92 $Y=4.07 $X2=0
+ $Y2=0
cc_101 N_VPB_c_71_n N_A_389_1337#_c_378_n 0.0244033f $X=7.92 $Y=4.07 $X2=4.08
+ $Y2=0
cc_102 N_VPB_c_71_n N_A_389_141#_c_445_n 0.0145164f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_103 N_VPB_c_71_n N_A_389_141#_c_451_n 0.0266466f $X=7.92 $Y=4.07 $X2=7.92
+ $Y2=8.14
cc_104 N_VPB_c_71_n N_A_389_141#_c_452_n 0.0331169f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_105 N_VPB_c_71_n N_A_389_141#_c_458_n 0.00397161f $X=7.92 $Y=4.07 $X2=4.08
+ $Y2=8.14
cc_106 N_VPB_M1015_b N_VPWR_c_531_n 0.0557649f $X=-0.33 $Y=1.885 $X2=-0.33
+ $Y2=-0.265
cc_107 N_VPB_M1015_b N_VPWR_c_532_n 0.0629033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_108 N_VPB_M1015_b N_VPWR_c_533_n 0.0169807f $X=-0.33 $Y=1.885 $X2=7.92 $Y2=0
cc_109 N_VPB_c_85_p N_VPWR_c_533_n 0.022423f $X=0.72 $Y=4.07 $X2=7.92 $Y2=0
cc_110 N_VPB_c_71_n N_VPWR_c_533_n 0.00163118f $X=7.92 $Y=4.07 $X2=7.92 $Y2=0
cc_111 N_VPB_M1015_b N_VPWR_c_536_n 0.0167014f $X=-0.33 $Y=1.885 $X2=0.24
+ $Y2=8.14
cc_112 N_VPB_c_85_p N_VPWR_c_536_n 0.0224257f $X=0.72 $Y=4.07 $X2=0.24 $Y2=8.14
cc_113 N_VPB_c_71_n N_VPWR_c_536_n 0.00162748f $X=7.92 $Y=4.07 $X2=0.24 $Y2=8.14
cc_114 N_VPB_M1015_b VPWR 0.0368664f $X=-0.33 $Y=1.885 $X2=7.92 $Y2=8.14
cc_115 N_VPB_X18_noxref_D1 VPWR 0.0422008f $X=7 $Y=1.885 $X2=7.92 $Y2=8.14
cc_116 N_VPB_c_85_p VPWR 0.00454266f $X=0.72 $Y=4.07 $X2=7.92 $Y2=8.14
cc_117 N_VPB_c_118_p VPWR 0.00678484f $X=7.92 $Y=4.07 $X2=7.92 $Y2=8.14
cc_118 N_VPB_c_71_n VPWR 0.84712f $X=7.92 $Y=4.07 $X2=7.92 $Y2=8.14
cc_119 N_VPB_M1015_b VPWR 0.0523976f $X=-0.33 $Y=1.885 $X2=4.08 $Y2=0
cc_120 N_VPB_X18_noxref_D1 VPWR 0.0764274f $X=7 $Y=1.885 $X2=4.08 $Y2=0
cc_121 N_VPB_c_85_p VPWR 0.00454266f $X=0.72 $Y=4.07 $X2=4.08 $Y2=0
cc_122 N_VPB_c_118_p VPWR 0.00678484f $X=7.92 $Y=4.07 $X2=4.08 $Y2=0
cc_123 N_VPB_c_71_n VPWR 0.849059f $X=7.92 $Y=4.07 $X2=4.08 $Y2=0
cc_124 N_VPB_c_71_n N_VGND_c_617_n 0.00710099f $X=7.92 $Y=4.07 $X2=0 $Y2=0
cc_125 N_LVPWR_c_126_n N_A_30_1337#_c_214_n 0.00980342f $X=4.605 $Y=3.19 $X2=0
+ $Y2=0
cc_126 N_LVPWR_c_126_n N_A_30_1337#_c_210_n 0.0715684f $X=4.605 $Y=3.19 $X2=0
+ $Y2=0
cc_127 N_LVPWR_c_126_n N_A_30_1337#_c_219_n 0.00467827f $X=4.605 $Y=3.19
+ $X2=4.32 $Y2=0.058
cc_128 N_LVPWR_c_126_n N_A_30_1337#_c_212_n 0.0202991f $X=4.605 $Y=3.19 $X2=4.32
+ $Y2=8.14
cc_129 N_LVPWR_c_126_n N_A_30_207#_M1007_g 0.0185311f $X=4.605 $Y=3.19 $X2=0.24
+ $Y2=0
cc_130 N_LVPWR_c_126_n N_A_30_207#_c_335_n 0.0014457f $X=4.605 $Y=3.19 $X2=0.24
+ $Y2=8.14
cc_131 N_LVPWR_c_128_n N_A_389_1337#_M1013_d 0.00148638f $X=4.265 $Y=4.085 $X2=0
+ $Y2=0
cc_132 N_LVPWR_c_126_n N_A_389_1337#_M1013_d 0.00259992f $X=4.605 $Y=3.19 $X2=0
+ $Y2=0
cc_133 N_LVPWR_M1003_b N_A_389_1337#_M1001_g 0.0272031f $X=3.53 $Y=1.925 $X2=0
+ $Y2=0
cc_134 N_LVPWR_c_128_n N_A_389_1337#_M1001_g 0.00592637f $X=4.265 $Y=4.085 $X2=0
+ $Y2=0
cc_135 N_LVPWR_c_129_n N_A_389_1337#_M1001_g 0.00695404f $X=4.265 $Y=4.42 $X2=0
+ $Y2=0
cc_136 N_LVPWR_M1003_b N_A_389_1337#_c_372_n 0.00221896f $X=3.53 $Y=1.925
+ $X2=7.92 $Y2=0
cc_137 N_LVPWR_M1003_b N_A_389_1337#_c_374_n 0.00160726f $X=3.53 $Y=1.925 $X2=0
+ $Y2=0
cc_138 N_LVPWR_c_129_n N_A_389_1337#_c_376_n 0.0213021f $X=4.265 $Y=4.42 $X2=0
+ $Y2=0
cc_139 N_LVPWR_M1003_b N_A_389_1337#_c_377_n 0.0155782f $X=3.53 $Y=1.925
+ $X2=7.92 $Y2=8.14
cc_140 N_LVPWR_c_129_n N_A_389_1337#_c_377_n 0.00617974f $X=4.265 $Y=4.42
+ $X2=7.92 $Y2=8.14
cc_141 N_LVPWR_M1003_b N_A_389_1337#_c_393_n 0.0073482f $X=3.53 $Y=1.925 $X2=0
+ $Y2=0
cc_142 N_LVPWR_c_149_p N_A_389_1337#_c_393_n 0.00152476f $X=4.265 $Y=2.25 $X2=0
+ $Y2=0
cc_143 N_LVPWR_M1003_b N_A_389_1337#_c_378_n 0.0365288f $X=3.53 $Y=1.925
+ $X2=4.08 $Y2=0
cc_144 N_LVPWR_c_149_p N_A_389_1337#_c_378_n 0.00299067f $X=4.265 $Y=2.25
+ $X2=4.08 $Y2=0
cc_145 N_LVPWR_c_128_n N_A_389_1337#_c_378_n 0.0764335f $X=4.265 $Y=4.085
+ $X2=4.08 $Y2=0
cc_146 N_LVPWR_c_129_n N_A_389_1337#_c_378_n 0.041929f $X=4.265 $Y=4.42 $X2=4.08
+ $Y2=0
cc_147 N_LVPWR_c_126_n N_A_389_1337#_c_378_n 0.0273372f $X=4.605 $Y=3.19
+ $X2=4.08 $Y2=0
cc_148 N_LVPWR_M1003_b N_A_389_1337#_c_380_n 0.00943291f $X=3.53 $Y=1.925 $X2=0
+ $Y2=0
cc_149 N_LVPWR_c_128_n N_A_389_1337#_c_380_n 0.00991797f $X=4.265 $Y=4.085 $X2=0
+ $Y2=0
cc_150 N_LVPWR_c_126_n N_A_389_1337#_c_380_n 0.0161079f $X=4.605 $Y=3.19 $X2=0
+ $Y2=0
cc_151 N_LVPWR_c_128_n N_A_389_141#_c_445_n 0.016492f $X=4.265 $Y=4.085 $X2=0
+ $Y2=0
cc_152 N_LVPWR_c_129_n N_A_389_141#_c_445_n 0.0010372f $X=4.265 $Y=4.42 $X2=0
+ $Y2=0
cc_153 N_LVPWR_c_126_n N_A_389_141#_c_445_n 0.0215479f $X=4.605 $Y=3.19 $X2=0
+ $Y2=0
cc_154 N_LVPWR_M1003_b N_A_389_141#_c_446_n 0.0103185f $X=3.53 $Y=1.925 $X2=0
+ $Y2=0
cc_155 N_LVPWR_M1003_b N_A_389_141#_M1003_g 0.018503f $X=3.53 $Y=1.925 $X2=7.92
+ $Y2=0
cc_156 N_LVPWR_c_149_p N_A_389_141#_M1003_g 4.70317e-19 $X=4.265 $Y=2.25
+ $X2=7.92 $Y2=0
cc_157 N_LVPWR_c_128_n N_A_389_141#_M1003_g 0.0116728f $X=4.265 $Y=4.085
+ $X2=7.92 $Y2=0
cc_158 N_LVPWR_c_126_n N_A_389_141#_M1003_g 0.00809621f $X=4.605 $Y=3.19
+ $X2=7.92 $Y2=0
cc_159 N_LVPWR_M1003_b N_A_389_141#_M1013_g 0.022397f $X=3.53 $Y=1.925 $X2=0
+ $Y2=0
cc_160 N_LVPWR_c_149_p N_A_389_141#_M1013_g 5.94561e-19 $X=4.265 $Y=2.25 $X2=0
+ $Y2=0
cc_161 N_LVPWR_c_128_n N_A_389_141#_M1013_g 0.0176706f $X=4.265 $Y=4.085 $X2=0
+ $Y2=0
cc_162 N_LVPWR_c_126_n N_A_389_141#_M1013_g 0.00740956f $X=4.605 $Y=3.19 $X2=0
+ $Y2=0
cc_163 N_LVPWR_M1003_b N_A_389_141#_c_450_n 0.00702821f $X=3.53 $Y=1.925 $X2=0
+ $Y2=0
cc_164 N_LVPWR_c_149_p N_A_389_141#_c_450_n 0.00309844f $X=4.265 $Y=2.25 $X2=0
+ $Y2=0
cc_165 N_LVPWR_c_126_n N_A_389_141#_c_451_n 0.0407972f $X=4.605 $Y=3.19 $X2=7.92
+ $Y2=8.14
cc_166 N_LVPWR_M1003_b N_A_389_141#_c_452_n 0.00461606f $X=3.53 $Y=1.925 $X2=0
+ $Y2=0
cc_167 N_LVPWR_M1003_b N_A_389_141#_c_458_n 0.00246153f $X=3.53 $Y=1.925
+ $X2=4.08 $Y2=8.14
cc_168 N_LVPWR_c_128_n N_A_389_141#_c_458_n 0.0133262f $X=4.265 $Y=4.085
+ $X2=4.08 $Y2=8.14
cc_169 N_LVPWR_c_129_n N_A_389_141#_c_458_n 0.0115197f $X=4.265 $Y=4.42 $X2=4.08
+ $Y2=8.14
cc_170 N_LVPWR_M1003_b N_A_389_141#_c_478_n 0.00198099f $X=3.53 $Y=1.925
+ $X2=4.32 $Y2=8.082
cc_171 N_LVPWR_c_129_n N_A_389_141#_c_478_n 0.00508153f $X=4.265 $Y=4.42
+ $X2=4.32 $Y2=8.082
cc_172 N_LVPWR_c_126_n N_VPWR_c_531_n 0.0466946f $X=4.605 $Y=3.19 $X2=-0.33
+ $Y2=-0.265
cc_173 N_LVPWR_c_126_n N_VPWR_c_533_n 0.00197188f $X=4.605 $Y=3.19 $X2=7.92
+ $Y2=0
cc_174 N_LVPWR_M1003_b VPWR 0.00424322f $X=3.53 $Y=1.925 $X2=7.92 $Y2=8.14
cc_175 N_LVPWR_c_128_n VPWR 0.0761117f $X=4.265 $Y=4.085 $X2=7.92 $Y2=8.14
cc_176 N_LVPWR_c_126_n VPWR 0.838276f $X=4.605 $Y=3.19 $X2=7.92 $Y2=8.14
cc_177 N_LVPWR_M1003_b VPWR 0.0327385f $X=3.53 $Y=1.925 $X2=4.08 $Y2=0
cc_178 N_LVPWR_c_128_n VPWR 0.0031715f $X=4.265 $Y=4.085 $X2=4.08 $Y2=0
cc_179 N_LVPWR_c_129_n VPWR 0.0423398f $X=4.265 $Y=4.42 $X2=4.08 $Y2=0
cc_180 N_LVPWR_c_126_n N_X_M1003_s 5.28909e-19 $X=4.605 $Y=3.19 $X2=0 $Y2=0
cc_181 N_LVPWR_M1003_b N_X_c_596_n 0.00665255f $X=3.53 $Y=1.925 $X2=0 $Y2=0
cc_182 N_LVPWR_c_149_p N_X_c_596_n 0.00357017f $X=4.265 $Y=2.25 $X2=0 $Y2=0
cc_183 N_LVPWR_c_128_n N_X_c_596_n 0.0202758f $X=4.265 $Y=4.085 $X2=0 $Y2=0
cc_184 N_LVPWR_c_126_n N_X_c_596_n 0.0514471f $X=4.605 $Y=3.19 $X2=0 $Y2=0
cc_185 N_LVPWR_c_128_n N_VGND_c_617_n 0.0102587f $X=4.265 $Y=4.085 $X2=0 $Y2=0
cc_186 N_LVPWR_c_126_n N_VGND_c_617_n 0.0704096f $X=4.605 $Y=3.19 $X2=0 $Y2=0
cc_187 N_LVPWR_c_149_p N_VGND_c_619_n 0.010688f $X=4.265 $Y=2.25 $X2=0 $Y2=0
cc_188 N_A_30_1337#_c_207_n N_A_M1000_g 0.00571833f $X=0.295 $Y=6.895 $X2=0
+ $Y2=0
cc_189 N_A_30_1337#_c_208_n N_A_M1000_g 0.0724091f $X=0.95 $Y=6.397 $X2=0 $Y2=0
cc_190 N_A_30_1337#_c_211_n N_A_M1000_g 0.0136055f $X=1.075 $Y=5.715 $X2=0 $Y2=0
cc_191 N_A_30_1337#_c_213_n N_A_M1000_g 0.0233088f $X=1.61 $Y=6.07 $X2=0 $Y2=0
cc_192 N_A_30_1337#_c_212_n N_A_c_296_n 0.00918492f $X=1.35 $Y=5.55 $X2=-0.33
+ $Y2=-0.265
cc_193 N_A_30_1337#_c_211_n A 0.0156547f $X=1.075 $Y=5.715 $X2=0 $Y2=8.025
cc_194 N_A_30_1337#_c_212_n A 0.0271564f $X=1.35 $Y=5.55 $X2=0 $Y2=8.025
cc_195 N_A_30_1337#_c_211_n N_A_c_299_n 0.00712362f $X=1.075 $Y=5.715 $X2=0.24
+ $Y2=0
cc_196 N_A_30_1337#_c_212_n N_A_c_299_n 0.00237131f $X=1.35 $Y=5.55 $X2=0.24
+ $Y2=0
cc_197 N_A_30_1337#_M1002_g N_A_30_207#_M1004_g 0.0218679f $X=0.685 $Y=1.245
+ $X2=-0.33 $Y2=-0.265
cc_198 N_A_30_1337#_c_210_n N_A_30_207#_c_322_n 0.00187442f $X=1.47 $Y=2.96
+ $X2=0 $Y2=0
cc_199 N_A_30_1337#_c_210_n N_A_30_207#_M1007_g 8.76986e-19 $X=1.47 $Y=2.96
+ $X2=0.24 $Y2=0
cc_200 N_A_30_1337#_c_212_n N_A_30_207#_M1007_g 0.00160599f $X=1.35 $Y=5.55
+ $X2=0.24 $Y2=0
cc_201 N_A_30_1337#_M1002_g N_A_30_207#_c_326_n 0.00571833f $X=0.685 $Y=1.245
+ $X2=7.92 $Y2=0
cc_202 N_A_30_1337#_M1002_g N_A_30_207#_c_327_n 0.0728299f $X=0.685 $Y=1.245
+ $X2=0 $Y2=0
cc_203 N_A_30_1337#_M1002_g N_A_30_207#_c_335_n 0.0104872f $X=0.685 $Y=1.245
+ $X2=0.24 $Y2=8.14
cc_204 N_A_30_1337#_c_210_n N_A_30_207#_c_335_n 0.01246f $X=1.47 $Y=2.96
+ $X2=0.24 $Y2=8.14
cc_205 N_A_30_1337#_c_219_n N_A_30_207#_c_335_n 0.0056527f $X=1.135 $Y=2.96
+ $X2=0.24 $Y2=8.14
cc_206 N_A_30_1337#_c_210_n N_A_30_207#_c_329_n 0.00982452f $X=1.47 $Y=2.96
+ $X2=7.92 $Y2=8.14
cc_207 N_A_30_1337#_c_196_n N_A_389_1337#_c_371_n 0.0269434f $X=1.695 $Y=6.61
+ $X2=0 $Y2=0
cc_208 N_A_30_1337#_c_198_n N_A_389_1337#_c_371_n 0.0109819f $X=2.225 $Y=6.535
+ $X2=0 $Y2=0
cc_209 N_A_30_1337#_c_199_n N_A_389_1337#_c_371_n 0.027654f $X=2.475 $Y=6.46
+ $X2=0 $Y2=0
cc_210 N_A_30_1337#_c_200_n N_A_389_1337#_c_371_n 0.0197273f $X=2.475 $Y=6.61
+ $X2=0 $Y2=0
cc_211 N_A_30_1337#_c_205_n N_A_389_1337#_c_371_n 0.00413022f $X=1.695 $Y=6.535
+ $X2=0 $Y2=0
cc_212 N_A_30_1337#_c_206_n N_A_389_1337#_c_371_n 0.00310572f $X=2.475 $Y=6.535
+ $X2=0 $Y2=0
cc_213 N_A_30_1337#_c_212_n N_A_389_1337#_c_371_n 0.0952854f $X=1.35 $Y=5.55
+ $X2=0 $Y2=0
cc_214 N_A_30_1337#_c_213_n N_A_389_1337#_c_371_n 0.00499425f $X=1.61 $Y=6.07
+ $X2=0 $Y2=0
cc_215 N_A_30_1337#_c_199_n N_A_389_1337#_c_372_n 0.0195038f $X=2.475 $Y=6.46
+ $X2=7.92 $Y2=0
cc_216 N_A_30_1337#_c_212_n N_A_389_1337#_c_373_n 0.0218587f $X=1.35 $Y=5.55
+ $X2=0 $Y2=0
cc_217 N_A_30_1337#_c_199_n N_A_389_1337#_c_374_n 0.00244389f $X=2.475 $Y=6.46
+ $X2=0 $Y2=0
cc_218 N_A_30_1337#_c_202_n N_A_389_1337#_c_375_n 0.00715826f $X=3.005 $Y=6.535
+ $X2=0.24 $Y2=8.14
cc_219 N_A_30_1337#_c_203_n N_A_389_1337#_c_375_n 0.0234318f $X=3.255 $Y=6.61
+ $X2=0.24 $Y2=8.14
cc_220 N_A_30_1337#_c_199_n N_A_389_1337#_c_379_n 9.97257e-19 $X=2.475 $Y=6.46
+ $X2=4.32 $Y2=0
cc_221 N_A_30_1337#_c_202_n N_A_389_1337#_c_379_n 0.00572917f $X=3.005 $Y=6.535
+ $X2=4.32 $Y2=0
cc_222 N_A_30_1337#_c_210_n N_A_389_141#_c_451_n 0.0211293f $X=1.47 $Y=2.96
+ $X2=7.92 $Y2=8.14
cc_223 N_A_30_1337#_c_219_n N_A_389_141#_c_451_n 0.00185275f $X=1.135 $Y=2.96
+ $X2=7.92 $Y2=8.14
cc_224 N_A_30_1337#_c_212_n N_A_389_141#_c_451_n 0.0876228f $X=1.35 $Y=5.55
+ $X2=7.92 $Y2=8.14
cc_225 N_A_30_1337#_c_212_n N_A_389_141#_c_453_n 0.0258593f $X=1.35 $Y=5.55
+ $X2=4.08 $Y2=0
cc_226 N_A_30_1337#_c_214_n N_VPWR_c_531_n 0.019601f $X=0.685 $Y=2.515 $X2=-0.33
+ $Y2=-0.265
cc_227 N_A_30_1337#_M1002_g N_VPWR_c_531_n 0.00669099f $X=0.685 $Y=1.245
+ $X2=-0.33 $Y2=-0.265
cc_228 N_A_30_1337#_c_210_n N_VPWR_c_531_n 0.0198736f $X=1.47 $Y=2.96 $X2=-0.33
+ $Y2=-0.265
cc_229 N_A_30_1337#_c_208_n N_VPWR_c_532_n 0.00144394f $X=0.95 $Y=6.397 $X2=0
+ $Y2=0
cc_230 N_A_30_1337#_c_209_n N_VPWR_c_532_n 0.0128286f $X=0.42 $Y=6.397 $X2=0
+ $Y2=0
cc_231 N_A_30_1337#_c_214_n N_VPWR_c_533_n 0.00481379f $X=0.685 $Y=2.515
+ $X2=7.92 $Y2=0
cc_232 N_A_30_1337#_c_210_n N_VPWR_c_533_n 0.00270294f $X=1.47 $Y=2.96 $X2=7.92
+ $Y2=0
cc_233 N_A_30_1337#_c_214_n VPWR 0.0030611f $X=0.685 $Y=2.515 $X2=7.92 $Y2=8.14
cc_234 N_A_30_1337#_c_210_n VPWR 0.0080616f $X=1.47 $Y=2.96 $X2=7.92 $Y2=8.14
cc_235 N_A_30_1337#_c_212_n VPWR 0.0354957f $X=1.35 $Y=5.55 $X2=7.92 $Y2=8.14
cc_236 N_A_30_1337#_c_212_n VPWR 0.0502411f $X=1.35 $Y=5.55 $X2=4.08 $Y2=0
cc_237 N_A_30_1337#_M1002_g N_VGND_c_611_n 0.0210102f $X=0.685 $Y=1.245 $X2=0
+ $Y2=0
cc_238 N_A_30_1337#_c_196_n N_VGND_c_613_n 0.0347688f $X=1.695 $Y=6.61 $X2=0
+ $Y2=0
cc_239 N_A_30_1337#_c_208_n N_VGND_c_613_n 0.00372166f $X=0.95 $Y=6.397 $X2=0
+ $Y2=0
cc_240 N_A_30_1337#_c_211_n N_VGND_c_613_n 0.0442967f $X=1.075 $Y=5.715 $X2=0
+ $Y2=0
cc_241 N_A_30_1337#_c_196_n N_VGND_c_615_n 8.23467e-19 $X=1.695 $Y=6.61 $X2=7.92
+ $Y2=0
cc_242 N_A_30_1337#_c_199_n N_VGND_c_615_n 0.0363562f $X=2.475 $Y=6.46 $X2=7.92
+ $Y2=0
cc_243 N_A_30_1337#_c_200_n N_VGND_c_615_n 0.0417041f $X=2.475 $Y=6.61 $X2=7.92
+ $Y2=0
cc_244 N_A_30_1337#_c_202_n N_VGND_c_615_n 0.0209666f $X=3.005 $Y=6.535 $X2=7.92
+ $Y2=0
cc_245 N_A_30_1337#_c_203_n N_VGND_c_615_n 0.0378199f $X=3.255 $Y=6.61 $X2=7.92
+ $Y2=0
cc_246 N_A_30_1337#_c_206_n N_VGND_c_615_n 0.00557872f $X=2.475 $Y=6.535
+ $X2=7.92 $Y2=0
cc_247 N_A_30_1337#_M1002_g N_VGND_c_621_n 0.0136209f $X=0.685 $Y=1.245 $X2=0
+ $Y2=0
cc_248 N_A_30_1337#_c_196_n VGND 0.026803f $X=1.695 $Y=6.61 $X2=0 $Y2=0
cc_249 N_A_30_1337#_c_200_n VGND 0.0175283f $X=2.475 $Y=6.61 $X2=0 $Y2=0
cc_250 N_A_30_1337#_c_203_n VGND 0.022837f $X=3.255 $Y=6.61 $X2=0 $Y2=0
cc_251 N_A_30_1337#_c_207_n VGND 0.0108023f $X=0.295 $Y=6.895 $X2=0 $Y2=0
cc_252 N_A_c_294_n N_VPWR_c_532_n 0.0135528f $X=0.685 $Y=5.625 $X2=0 $Y2=0
cc_253 N_A_M1000_g N_VPWR_c_532_n 0.00667092f $X=0.685 $Y=5.715 $X2=0 $Y2=0
cc_254 N_A_c_297_n N_VPWR_c_532_n 0.0094178f $X=0.935 $Y=5.035 $X2=0 $Y2=0
cc_255 A N_VPWR_c_532_n 0.0274931f $X=1.115 $Y=4.91 $X2=0 $Y2=0
cc_256 N_A_c_294_n N_VPWR_c_536_n 0.00347108f $X=0.685 $Y=5.625 $X2=0.24
+ $Y2=8.14
cc_257 N_A_c_297_n N_VPWR_c_536_n 0.00232677f $X=0.935 $Y=5.035 $X2=0.24
+ $Y2=8.14
cc_258 A N_VPWR_c_536_n 0.00576436f $X=1.115 $Y=4.91 $X2=0.24 $Y2=8.14
cc_259 N_A_c_297_n VPWR 0.019692f $X=0.935 $Y=5.035 $X2=4.08 $Y2=0
cc_260 A VPWR 0.0311181f $X=1.115 $Y=4.91 $X2=4.08 $Y2=0
cc_261 N_A_M1000_g N_VGND_c_613_n 0.0303358f $X=0.685 $Y=5.715 $X2=0 $Y2=0
cc_262 N_A_M1000_g VGND 0.0147494f $X=0.685 $Y=5.715 $X2=0 $Y2=0
cc_263 N_A_30_207#_c_322_n N_A_389_141#_c_445_n 0.0204856f $X=2.475 $Y=1.65
+ $X2=0 $Y2=0
cc_264 N_A_30_207#_M1006_g N_A_389_141#_c_447_n 0.0204856f $X=2.475 $Y=1.08
+ $X2=0.24 $Y2=0
cc_265 N_A_30_207#_M1004_g N_A_389_141#_c_451_n 0.0312302f $X=1.695 $Y=1.08
+ $X2=7.92 $Y2=8.14
cc_266 N_A_30_207#_c_322_n N_A_389_141#_c_451_n 0.0314645f $X=2.475 $Y=1.65
+ $X2=7.92 $Y2=8.14
cc_267 N_A_30_207#_M1006_g N_A_389_141#_c_451_n 0.0247916f $X=2.475 $Y=1.08
+ $X2=7.92 $Y2=8.14
cc_268 N_A_30_207#_M1007_g N_A_389_141#_c_451_n 0.0560519f $X=2.475 $Y=2.5
+ $X2=7.92 $Y2=8.14
cc_269 N_A_30_207#_c_329_n N_A_389_141#_c_451_n 0.0264057f $X=1.597 $Y=1.73
+ $X2=7.92 $Y2=8.14
cc_270 N_A_30_207#_c_330_n N_A_389_141#_c_451_n 0.0261027f $X=1.61 $Y=1.73
+ $X2=7.92 $Y2=8.14
cc_271 N_A_30_207#_M1007_g N_A_389_141#_c_452_n 0.014357f $X=2.475 $Y=2.5 $X2=0
+ $Y2=0
cc_272 N_A_30_207#_c_327_n N_VPWR_c_531_n 0.00135625f $X=0.95 $Y=1.73 $X2=-0.33
+ $Y2=-0.265
cc_273 N_A_30_207#_c_328_n N_VPWR_c_531_n 0.0121965f $X=0.42 $Y=1.73 $X2=-0.33
+ $Y2=-0.265
cc_274 N_A_30_207#_M1007_g VPWR 0.00700858f $X=2.475 $Y=2.5 $X2=7.92 $Y2=8.14
cc_275 N_A_30_207#_M1004_g N_VGND_c_611_n 0.034756f $X=1.695 $Y=1.08 $X2=0 $Y2=0
cc_276 N_A_30_207#_c_327_n N_VGND_c_611_n 0.0452382f $X=0.95 $Y=1.73 $X2=0 $Y2=0
cc_277 N_A_30_207#_M1004_g N_VGND_c_617_n 8.52469e-19 $X=1.695 $Y=1.08 $X2=0
+ $Y2=0
cc_278 N_A_30_207#_c_322_n N_VGND_c_617_n 0.0166231f $X=2.475 $Y=1.65 $X2=0
+ $Y2=0
cc_279 N_A_30_207#_M1006_g N_VGND_c_617_n 0.0475723f $X=2.475 $Y=1.08 $X2=0
+ $Y2=0
cc_280 N_A_30_207#_M1007_g N_VGND_c_617_n 0.0727695f $X=2.475 $Y=2.5 $X2=0 $Y2=0
cc_281 N_A_30_207#_M1004_g N_VGND_c_621_n 0.026803f $X=1.695 $Y=1.08 $X2=0 $Y2=0
cc_282 N_A_30_207#_M1006_g N_VGND_c_621_n 0.0199218f $X=2.475 $Y=1.08 $X2=0
+ $Y2=0
cc_283 N_A_30_207#_c_326_n N_VGND_c_621_n 0.0108023f $X=0.295 $Y=1.245 $X2=0
+ $Y2=0
cc_284 N_A_389_1337#_M1001_g N_A_389_141#_c_445_n 0.00684085f $X=4.05 $Y=4.835
+ $X2=0 $Y2=0
cc_285 N_A_389_1337#_c_372_n N_A_389_141#_c_445_n 0.0025108f $X=3.29 $Y=5.32
+ $X2=0 $Y2=0
cc_286 N_A_389_1337#_c_393_n N_A_389_141#_M1013_g 0.00246524f $X=4.695 $Y=2.25
+ $X2=0 $Y2=0
cc_287 N_A_389_1337#_c_378_n N_A_389_141#_M1013_g 0.00354403f $X=5.045 $Y=5.595
+ $X2=0 $Y2=0
cc_288 N_A_389_1337#_c_372_n N_A_389_141#_c_452_n 0.0207526f $X=3.29 $Y=5.32
+ $X2=0 $Y2=0
cc_289 N_A_389_1337#_c_373_n N_A_389_141#_c_453_n 0.00637574f $X=2.25 $Y=5.32
+ $X2=4.08 $Y2=0
cc_290 N_A_389_1337#_M1001_g N_A_389_141#_c_458_n 6.48264e-19 $X=4.05 $Y=4.835
+ $X2=4.08 $Y2=8.14
cc_291 N_A_389_1337#_M1001_g N_A_389_141#_c_478_n 0.00154299f $X=4.05 $Y=4.835
+ $X2=4.32 $Y2=8.082
cc_292 N_A_389_1337#_c_372_n N_A_389_141#_c_478_n 0.0187941f $X=3.29 $Y=5.32
+ $X2=4.32 $Y2=8.082
cc_293 N_A_389_1337#_c_376_n N_A_389_141#_c_478_n 0.0117776f $X=4.92 $Y=5.72
+ $X2=4.32 $Y2=8.082
cc_294 N_A_389_1337#_c_377_n N_A_389_141#_c_478_n 0.00593478f $X=4.22 $Y=5.72
+ $X2=4.32 $Y2=8.082
cc_295 N_A_389_1337#_c_379_n N_A_389_141#_c_478_n 0.00846878f $X=3.55 $Y=5.72
+ $X2=4.32 $Y2=8.082
cc_296 N_A_389_1337#_c_372_n N_A_389_141#_c_454_n 0.00485191f $X=3.29 $Y=5.32
+ $X2=0 $Y2=0
cc_297 N_A_389_1337#_c_378_n VPWR 0.033301f $X=5.045 $Y=5.595 $X2=7.92 $Y2=8.14
cc_298 N_A_389_1337#_M1001_g VPWR 0.00830624f $X=4.05 $Y=4.835 $X2=4.08 $Y2=0
cc_299 N_A_389_1337#_c_372_n VPWR 0.0326833f $X=3.29 $Y=5.32 $X2=4.08 $Y2=0
cc_300 N_A_389_1337#_c_373_n VPWR 0.00868385f $X=2.25 $Y=5.32 $X2=4.08 $Y2=0
cc_301 N_A_389_1337#_c_378_n VPWR 0.0490299f $X=5.045 $Y=5.595 $X2=4.08 $Y2=0
cc_302 N_A_389_1337#_c_371_n N_VGND_c_613_n 0.0260785f $X=2.085 $Y=5.78 $X2=0
+ $Y2=0
cc_303 N_A_389_1337#_c_371_n N_VGND_c_615_n 0.0968722f $X=2.085 $Y=5.78 $X2=7.92
+ $Y2=0
cc_304 N_A_389_1337#_c_372_n N_VGND_c_615_n 0.0501196f $X=3.29 $Y=5.32 $X2=7.92
+ $Y2=0
cc_305 N_A_389_1337#_c_375_n N_VGND_c_615_n 0.074602f $X=3.645 $Y=6.83 $X2=7.92
+ $Y2=0
cc_306 N_A_389_1337#_c_377_n N_VGND_c_615_n 9.46477e-19 $X=4.22 $Y=5.72 $X2=7.92
+ $Y2=0
cc_307 N_A_389_1337#_c_379_n N_VGND_c_615_n 0.0212281f $X=3.55 $Y=5.72 $X2=7.92
+ $Y2=0
cc_308 N_A_389_1337#_c_393_n N_VGND_c_619_n 0.00587594f $X=4.695 $Y=2.25 $X2=0
+ $Y2=0
cc_309 N_A_389_1337#_c_371_n VGND 0.014218f $X=2.085 $Y=5.78 $X2=0 $Y2=0
cc_310 N_A_389_1337#_c_375_n VGND 0.0143529f $X=3.645 $Y=6.83 $X2=0 $Y2=0
cc_311 N_A_389_141#_c_445_n VPWR 0.0184873f $X=3.335 $Y=4.265 $X2=7.92 $Y2=8.14
cc_312 N_A_389_141#_c_451_n VPWR 0.0320303f $X=2.085 $Y=0.85 $X2=7.92 $Y2=8.14
cc_313 N_A_389_141#_M1001_s VPWR 6.02657e-19 $X=3.71 $Y=4.275 $X2=4.08 $Y2=0
cc_314 N_A_389_141#_c_445_n VPWR 0.00321729f $X=3.335 $Y=4.265 $X2=4.08 $Y2=0
cc_315 N_A_389_141#_c_452_n VPWR 0.0755659f $X=3.71 $Y=4.425 $X2=4.08 $Y2=0
cc_316 N_A_389_141#_c_453_n VPWR 0.0218642f $X=2.25 $Y=4.425 $X2=4.08 $Y2=0
cc_317 N_A_389_141#_c_458_n VPWR 0.0119352f $X=3.835 $Y=4.595 $X2=4.08 $Y2=0
cc_318 N_A_389_141#_c_478_n VPWR 0.0211576f $X=3.835 $Y=5.25 $X2=4.08 $Y2=0
cc_319 N_A_389_141#_c_454_n VPWR 0.00330503f $X=3.17 $Y=4.43 $X2=4.08 $Y2=0
cc_320 N_A_389_141#_c_445_n N_X_c_596_n 0.0427695f $X=3.335 $Y=4.265 $X2=0 $Y2=0
cc_321 N_A_389_141#_c_446_n N_X_c_596_n 0.048541f $X=3.975 $Y=1.8 $X2=0 $Y2=0
cc_322 N_A_389_141#_c_447_n N_X_c_596_n 0.00617995f $X=3.5 $Y=1.8 $X2=0 $Y2=0
cc_323 N_A_389_141#_M1011_g N_X_c_596_n 0.00765192f $X=4.05 $Y=1.125 $X2=0 $Y2=0
cc_324 N_A_389_141#_M1003_g N_X_c_596_n 0.00503276f $X=4.05 $Y=2.665 $X2=0 $Y2=0
cc_325 N_A_389_141#_c_451_n N_VGND_c_611_n 0.0260785f $X=2.085 $Y=0.85 $X2=0
+ $Y2=0
cc_326 N_A_389_141#_c_447_n N_VGND_c_617_n 0.0386285f $X=3.5 $Y=1.8 $X2=0 $Y2=0
cc_327 N_A_389_141#_c_451_n N_VGND_c_617_n 0.142032f $X=2.085 $Y=0.85 $X2=0
+ $Y2=0
cc_328 N_A_389_141#_c_452_n N_VGND_c_617_n 0.0153592f $X=3.71 $Y=4.425 $X2=0
+ $Y2=0
cc_329 N_A_389_141#_c_454_n N_VGND_c_617_n 0.00233733f $X=3.17 $Y=4.43 $X2=0
+ $Y2=0
cc_330 N_A_389_141#_M1011_g N_VGND_c_619_n 0.00744837f $X=4.05 $Y=1.125 $X2=0
+ $Y2=0
cc_331 N_A_389_141#_c_450_n N_VGND_c_619_n 0.0169724f $X=4.48 $Y=1.8 $X2=0 $Y2=0
cc_332 N_A_389_141#_M1011_g N_VGND_c_621_n 0.00523016f $X=4.05 $Y=1.125 $X2=0
+ $Y2=0
cc_333 N_A_389_141#_c_451_n N_VGND_c_621_n 0.014218f $X=2.085 $Y=0.85 $X2=0
+ $Y2=0
cc_334 VPWR N_X_c_596_n 0.00225327f $X=4.32 $Y=3.63 $X2=0 $Y2=0
cc_335 VPWR N_VGND_c_617_n 0.0518341f $X=4.32 $Y=3.63 $X2=0 $Y2=0
cc_336 N_X_c_596_n N_VGND_c_617_n 0.131929f $X=3.835 $Y=0.9 $X2=0 $Y2=0
cc_337 N_X_c_596_n N_VGND_c_619_n 0.00339639f $X=3.835 $Y=0.9 $X2=0 $Y2=0
cc_338 N_X_c_596_n N_VGND_c_621_n 0.0199684f $X=3.835 $Y=0.9 $X2=0 $Y2=0
