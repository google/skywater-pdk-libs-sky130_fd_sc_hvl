* File: sky130_fd_sc_hvl__decap_4.pex.spice
* Created: Fri Aug 28 09:33:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__DECAP_4%VNB 5 7 11 25
r10 7 25 6.64328e-05 $w=1.92e-06 $l=1e-09 $layer=MET1_cond $X=0.96 $Y=0.057
+ $X2=0.96 $Y2=0.058
r11 7 11 0.00378667 $w=1.92e-06 $l=5.7e-08 $layer=MET1_cond $X=0.96 $Y=0.057
+ $X2=0.96 $Y2=0
r12 5 11 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r13 5 11 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__DECAP_4%VPB 4 6 14 21
r12 10 21 0.00378667 $w=1.92e-06 $l=5.7e-08 $layer=MET1_cond $X=0.96 $Y=4.07
+ $X2=0.96 $Y2=4.013
r13 10 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=4.07
+ $X2=1.68 $Y2=4.07
r14 9 14 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=1.68 $Y2=4.07
r15 9 10 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r16 6 21 6.64328e-05 $w=1.92e-06 $l=1e-09 $layer=MET1_cond $X=0.96 $Y=4.012
+ $X2=0.96 $Y2=4.013
r17 4 14 91 $w=1.7e-07 $l=1.72198e-06 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=1.68 $Y2=4.07
r18 4 9 91 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__DECAP_4%VGND 1 9 14 15 17 21 26
r26 32 33 5.39275 $w=6.9e-07 $l=3.05e-07 $layer=LI1_cond $X=0.335 $Y=0.807
+ $X2=0.64 $Y2=0.807
r27 29 32 0.618841 $w=6.9e-07 $l=3.5e-08 $layer=LI1_cond $X=0.3 $Y=0.807
+ $X2=0.335 $Y2=0.807
r28 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.3 $Y=0.48 $X2=0.3
+ $Y2=0.48
r29 23 26 0.275706 $w=8.83e-07 $l=2e-08 $layer=LI1_cond $X=1.595 $Y=0.807
+ $X2=1.615 $Y2=0.807
r30 23 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.595 $Y=0.48
+ $X2=1.595 $Y2=0.48
r31 21 33 2.89971 $w=8.85e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=0.807
+ $X2=0.64 $Y2=0.807
r32 21 23 10.8904 $w=8.83e-07 $l=7.9e-07 $layer=LI1_cond $X=0.805 $Y=0.807
+ $X2=1.595 $Y2=0.807
r33 17 30 0.00265731 $w=1.92e-06 $l=4e-08 $layer=MET1_cond $X=0.96 $Y=0.44
+ $X2=0.96 $Y2=0.48
r34 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.865 $X2=0.64 $Y2=1.865
r35 12 33 5.06645 $w=3.3e-07 $l=4.43e-07 $layer=LI1_cond $X=0.64 $Y=1.25
+ $X2=0.64 $Y2=0.807
r36 12 14 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.64 $Y=1.25
+ $X2=0.64 $Y2=1.865
r37 10 15 124.152 $w=3.3e-07 $l=7.1e-07 $layer=POLY_cond $X=0.64 $Y=2.575
+ $X2=0.64 $Y2=1.865
r38 9 10 57.2398 $w=1e-06 $l=6.3e-07 $layer=POLY_cond $X=0.975 $Y=3.205
+ $X2=0.975 $Y2=2.575
r39 1 32 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.595 $X2=0.335 $Y2=0.76
r40 1 26 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=1.475
+ $Y=0.595 $X2=1.615 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HVL__DECAP_4%VPWR 1 7 9 12 13 15 29 31
r24 28 31 2.62243 $w=1.068e-06 $l=2.3e-07 $layer=LI1_cond $X=1.385 $Y=3.22
+ $X2=1.615 $Y2=3.22
r25 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.385 $Y=3.645
+ $X2=1.385 $Y2=3.645
r26 26 28 2.33738 $w=1.068e-06 $l=2.05e-07 $layer=LI1_cond $X=1.18 $Y=3.22
+ $X2=1.385 $Y2=3.22
r27 24 26 6.84112 $w=1.068e-06 $l=6e-07 $layer=LI1_cond $X=0.58 $Y=3.22 $X2=1.18
+ $Y2=3.22
r28 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.58 $Y=3.645
+ $X2=0.58 $Y2=3.645
r29 20 24 2.79346 $w=1.068e-06 $l=2.45e-07 $layer=LI1_cond $X=0.335 $Y=3.22
+ $X2=0.58 $Y2=3.22
r30 15 29 0.16316 $w=3.7e-07 $l=4.25e-07 $layer=MET1_cond $X=0.96 $Y=3.63
+ $X2=1.385 $Y2=3.63
r31 15 25 0.145884 $w=3.7e-07 $l=3.8e-07 $layer=MET1_cond $X=0.96 $Y=3.63
+ $X2=0.58 $Y2=3.63
r32 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.865 $X2=1.18 $Y2=1.865
r33 10 26 7.77329 $w=3.3e-07 $l=5.35e-07 $layer=LI1_cond $X=1.18 $Y=2.685
+ $X2=1.18 $Y2=3.22
r34 10 12 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=1.18 $Y=2.685
+ $X2=1.18 $Y2=1.865
r35 7 13 47.1522 $w=4.6e-07 $l=3.9e-07 $layer=POLY_cond $X=1.245 $Y=1.475
+ $X2=1.245 $Y2=1.865
r36 7 9 38.5285 $w=1e-06 $l=5.15393e-07 $layer=POLY_cond $X=1.245 $Y=1.475
+ $X2=1.224 $Y2=0.97
r37 1 31 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.475
+ $Y=2.705 $X2=1.615 $Y2=3.56
r38 1 31 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.475
+ $Y=2.705 $X2=1.615 $Y2=2.85
r39 1 20 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.475
+ $Y=2.705 $X2=0.335 $Y2=3.56
r40 1 20 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.475
+ $Y=2.705 $X2=0.335 $Y2=2.85
.ends

