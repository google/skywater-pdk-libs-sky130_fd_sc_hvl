# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__inv_16
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__inv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  18.00000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  1.400000 1.565000  2.290000 1.895000 ;
        RECT  2.960000 1.565000  3.850000 1.895000 ;
        RECT  4.520000 1.565000  5.410000 1.895000 ;
        RECT  6.080000 1.565000  6.970000 1.895000 ;
        RECT  7.640000 1.565000  8.530000 1.895000 ;
        RECT  9.200000 1.565000 10.090000 1.895000 ;
        RECT 10.760000 1.565000 11.650000 1.895000 ;
      LAYER mcon ;
        RECT  1.595000 1.580000  1.765000 1.750000 ;
        RECT  1.955000 1.580000  2.125000 1.750000 ;
        RECT  3.145000 1.580000  3.315000 1.750000 ;
        RECT  3.505000 1.580000  3.675000 1.750000 ;
        RECT  4.705000 1.580000  4.875000 1.750000 ;
        RECT  5.065000 1.580000  5.235000 1.750000 ;
        RECT  6.265000 1.580000  6.435000 1.750000 ;
        RECT  6.625000 1.580000  6.795000 1.750000 ;
        RECT  7.825000 1.580000  7.995000 1.750000 ;
        RECT  8.185000 1.580000  8.355000 1.750000 ;
        RECT  9.385000 1.580000  9.555000 1.750000 ;
        RECT  9.745000 1.580000  9.915000 1.750000 ;
        RECT 10.945000 1.580000 11.115000 1.750000 ;
        RECT 11.305000 1.580000 11.475000 1.750000 ;
      LAYER met1 ;
        RECT  1.535000 1.550000  2.185000 1.580000 ;
        RECT  1.535000 1.580000 11.535000 1.750000 ;
        RECT  1.535000 1.750000  2.185000 1.780000 ;
        RECT  3.085000 1.550000  3.735000 1.580000 ;
        RECT  3.085000 1.750000  3.735000 1.780000 ;
        RECT  4.645000 1.550000  5.295000 1.580000 ;
        RECT  4.645000 1.750000  5.295000 1.780000 ;
        RECT  6.205000 1.550000  6.855000 1.580000 ;
        RECT  6.205000 1.750000  6.855000 1.780000 ;
        RECT  7.765000 1.550000  8.415000 1.580000 ;
        RECT  7.765000 1.750000  8.415000 1.780000 ;
        RECT  9.325000 1.550000  9.975000 1.580000 ;
        RECT  9.325000 1.750000  9.975000 1.780000 ;
        RECT 10.885000 1.550000 11.535000 1.580000 ;
        RECT 10.885000 1.750000 11.535000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  5.040000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.900000 0.795000  1.230000 3.755000 ;
        RECT  2.460000 0.795000  2.790000 3.755000 ;
        RECT  4.020000 0.795000  4.350000 3.755000 ;
        RECT  5.580000 0.795000  5.910000 3.755000 ;
        RECT  7.140000 0.795000  7.470000 3.755000 ;
        RECT  8.700000 0.795000  9.030000 3.755000 ;
        RECT 10.260000 0.795000 10.590000 3.755000 ;
        RECT 11.820000 0.795000 12.150000 3.755000 ;
      LAYER mcon ;
        RECT  0.985000 2.320000  1.155000 2.490000 ;
        RECT  2.545000 2.320000  2.715000 2.490000 ;
        RECT  4.105000 2.320000  4.275000 2.490000 ;
        RECT  5.665000 2.320000  5.835000 2.490000 ;
        RECT  7.225000 2.320000  7.395000 2.490000 ;
        RECT  8.785000 2.320000  8.955000 2.490000 ;
        RECT 10.345000 2.320000 10.515000 2.490000 ;
        RECT 11.905000 2.320000 12.075000 2.490000 ;
      LAYER met1 ;
        RECT  0.925000 2.290000  1.215000 2.320000 ;
        RECT  0.925000 2.320000 12.135000 2.490000 ;
        RECT  0.925000 2.490000  1.215000 2.520000 ;
        RECT  2.485000 2.290000  2.775000 2.320000 ;
        RECT  2.485000 2.490000  2.775000 2.520000 ;
        RECT  4.045000 2.290000  4.335000 2.320000 ;
        RECT  4.045000 2.490000  4.335000 2.520000 ;
        RECT  5.605000 2.290000  5.895000 2.320000 ;
        RECT  5.605000 2.490000  5.895000 2.520000 ;
        RECT  7.165000 2.290000  7.455000 2.320000 ;
        RECT  7.165000 2.490000  7.455000 2.520000 ;
        RECT  8.725000 2.290000  9.015000 2.320000 ;
        RECT  8.725000 2.490000  9.015000 2.520000 ;
        RECT 10.285000 2.290000 10.575000 2.320000 ;
        RECT 10.285000 2.490000 10.575000 2.520000 ;
        RECT 11.845000 2.290000 12.135000 2.320000 ;
        RECT 11.845000 2.490000 12.135000 2.520000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.095000 0.375000  0.630000 1.475000 ;
        RECT  1.400000 0.375000  2.290000 1.395000 ;
        RECT  2.960000 0.375000  3.850000 1.395000 ;
        RECT  4.520000 0.375000  5.410000 1.395000 ;
        RECT  6.080000 0.375000  6.970000 1.395000 ;
        RECT  7.640000 0.375000  8.530000 1.395000 ;
        RECT  9.200000 0.375000 10.090000 1.395000 ;
        RECT 10.760000 0.375000 11.650000 1.395000 ;
        RECT 12.320000 0.375000 12.935000 1.395000 ;
      LAYER mcon ;
        RECT  0.095000 0.425000  0.265000 0.595000 ;
        RECT  0.455000 0.425000  0.625000 0.595000 ;
        RECT  1.400000 0.425000  1.570000 0.595000 ;
        RECT  1.760000 0.425000  1.930000 0.595000 ;
        RECT  2.120000 0.425000  2.290000 0.595000 ;
        RECT  2.960000 0.425000  3.130000 0.595000 ;
        RECT  3.320000 0.425000  3.490000 0.595000 ;
        RECT  3.680000 0.425000  3.850000 0.595000 ;
        RECT  4.520000 0.425000  4.690000 0.595000 ;
        RECT  4.880000 0.425000  5.050000 0.595000 ;
        RECT  5.240000 0.425000  5.410000 0.595000 ;
        RECT  6.080000 0.425000  6.250000 0.595000 ;
        RECT  6.440000 0.425000  6.610000 0.595000 ;
        RECT  6.800000 0.425000  6.970000 0.595000 ;
        RECT  7.640000 0.425000  7.810000 0.595000 ;
        RECT  8.000000 0.425000  8.170000 0.595000 ;
        RECT  8.360000 0.425000  8.530000 0.595000 ;
        RECT  9.200000 0.425000  9.370000 0.595000 ;
        RECT  9.560000 0.425000  9.730000 0.595000 ;
        RECT  9.920000 0.425000 10.090000 0.595000 ;
        RECT 10.760000 0.425000 10.930000 0.595000 ;
        RECT 11.120000 0.425000 11.290000 0.595000 ;
        RECT 11.480000 0.425000 11.650000 0.595000 ;
        RECT 12.365000 0.425000 12.535000 0.595000 ;
        RECT 12.725000 0.425000 12.895000 0.595000 ;
      LAYER met1 ;
        RECT 0.000000 0.255000 13.440000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 13.440000 0.085000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.115000 13.440000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 13.440000 4.155000 ;
      LAYER mcon ;
        RECT  0.155000 3.985000  0.325000 4.155000 ;
        RECT  0.635000 3.985000  0.805000 4.155000 ;
        RECT  1.115000 3.985000  1.285000 4.155000 ;
        RECT  1.595000 3.985000  1.765000 4.155000 ;
        RECT  2.075000 3.985000  2.245000 4.155000 ;
        RECT  2.555000 3.985000  2.725000 4.155000 ;
        RECT  3.035000 3.985000  3.205000 4.155000 ;
        RECT  3.515000 3.985000  3.685000 4.155000 ;
        RECT  3.995000 3.985000  4.165000 4.155000 ;
        RECT  4.475000 3.985000  4.645000 4.155000 ;
        RECT  4.955000 3.985000  5.125000 4.155000 ;
        RECT  5.435000 3.985000  5.605000 4.155000 ;
        RECT  5.915000 3.985000  6.085000 4.155000 ;
        RECT  6.395000 3.985000  6.565000 4.155000 ;
        RECT  6.875000 3.985000  7.045000 4.155000 ;
        RECT  7.355000 3.985000  7.525000 4.155000 ;
        RECT  7.835000 3.985000  8.005000 4.155000 ;
        RECT  8.315000 3.985000  8.485000 4.155000 ;
        RECT  8.795000 3.985000  8.965000 4.155000 ;
        RECT  9.275000 3.985000  9.445000 4.155000 ;
        RECT  9.755000 3.985000  9.925000 4.155000 ;
        RECT 10.235000 3.985000 10.405000 4.155000 ;
        RECT 10.715000 3.985000 10.885000 4.155000 ;
        RECT 11.195000 3.985000 11.365000 4.155000 ;
        RECT 11.675000 3.985000 11.845000 4.155000 ;
        RECT 12.155000 3.985000 12.325000 4.155000 ;
        RECT 12.635000 3.985000 12.805000 4.155000 ;
        RECT 13.115000 3.985000 13.285000 4.155000 ;
      LAYER met1 ;
        RECT 0.000000 3.955000 13.440000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.125000 2.175000  0.655000 3.755000 ;
        RECT  1.400000 2.175000  2.290000 3.755000 ;
        RECT  2.960000 2.175000  3.850000 3.755000 ;
        RECT  4.520000 2.175000  5.410000 3.755000 ;
        RECT  6.080000 2.175000  6.970000 3.755000 ;
        RECT  7.640000 2.175000  8.530000 3.755000 ;
        RECT  9.200000 2.175000 10.090000 3.755000 ;
        RECT 10.760000 2.175000 11.650000 3.755000 ;
        RECT 12.320000 2.175000 12.935000 3.675000 ;
      LAYER mcon ;
        RECT  0.125000 3.475000  0.295000 3.645000 ;
        RECT  0.485000 3.475000  0.655000 3.645000 ;
        RECT  1.400000 3.475000  1.570000 3.645000 ;
        RECT  1.760000 3.475000  1.930000 3.645000 ;
        RECT  2.120000 3.475000  2.290000 3.645000 ;
        RECT  2.960000 3.475000  3.130000 3.645000 ;
        RECT  3.320000 3.475000  3.490000 3.645000 ;
        RECT  3.680000 3.475000  3.850000 3.645000 ;
        RECT  4.520000 3.475000  4.690000 3.645000 ;
        RECT  4.880000 3.475000  5.050000 3.645000 ;
        RECT  5.240000 3.475000  5.410000 3.645000 ;
        RECT  6.080000 3.475000  6.250000 3.645000 ;
        RECT  6.440000 3.475000  6.610000 3.645000 ;
        RECT  6.800000 3.475000  6.970000 3.645000 ;
        RECT  7.640000 3.475000  7.810000 3.645000 ;
        RECT  8.000000 3.475000  8.170000 3.645000 ;
        RECT  8.360000 3.475000  8.530000 3.645000 ;
        RECT  9.200000 3.475000  9.370000 3.645000 ;
        RECT  9.560000 3.475000  9.730000 3.645000 ;
        RECT  9.920000 3.475000 10.090000 3.645000 ;
        RECT 10.760000 3.475000 10.930000 3.645000 ;
        RECT 11.120000 3.475000 11.290000 3.645000 ;
        RECT 11.480000 3.475000 11.650000 3.645000 ;
        RECT 12.365000 3.475000 12.535000 3.645000 ;
        RECT 12.725000 3.475000 12.895000 3.645000 ;
      LAYER met1 ;
        RECT 0.000000 3.445000 13.440000 3.815000 ;
    END
  END VPWR
END sky130_fd_sc_hvl__inv_16
