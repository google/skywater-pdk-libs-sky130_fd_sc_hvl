* File: sky130_fd_sc_hvl__sdfrtp_1.spice
* Created: Fri Aug 28 09:39:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__sdfrtp_1.pex.spice"
.subckt sky130_fd_sc_hvl__sdfrtp_1  VNB VPB SCD SCE D RESET_B CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* D	D
* SCE	SCE
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1002 noxref_24 N_SCD_M1002_g N_noxref_23_M1002_s N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250000 SB=250004 A=0.21 P=1.84 MULT=1
MM1016 N_A_65_649#_M1016_d N_SCE_M1016_g noxref_24 N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250001 SB=250003 A=0.21 P=1.84 MULT=1
MM1038 noxref_25 N_A_116_451#_M1038_g N_A_65_649#_M1016_d N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1004 N_noxref_23_M1004_d N_D_M1004_g noxref_25 N_VNB_M1002_b NHV L=0.5 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250002
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1024 N_VGND_M1024_d N_RESET_B_M1024_g N_noxref_23_M1004_d N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250003 SB=250001 A=0.21 P=1.84 MULT=1
MM1012 N_A_116_451#_M1012_d N_SCE_M1012_g N_VGND_M1024_d N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250004
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1022 N_A_1312_126#_M1022_d N_A_1212_100#_M1022_g N_A_65_649#_M1022_s
+ N_VNB_M1002_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1001 A_1468_126# N_A_1212_471#_M1001_g N_A_1312_126#_M1022_d N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1010 A_1610_126# N_A_1510_100#_M1010_g A_1468_126# N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=13.566 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1013 N_VGND_M1013_d N_RESET_B_M1013_g A_1610_126# N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1032 N_VGND_M1032_d N_A_1212_100#_M1032_g N_A_1212_471#_M1032_s N_VNB_M1002_b
+ NHV L=0.5 W=0.42 AD=0.0973538 AS=0.1113 PD=0.832821 PS=1.37 NRD=25.7754 NRS=0
+ M=1 R=0.84 SA=250000 SB=250005 A=0.21 P=1.84 MULT=1
MM1007 N_A_1510_100#_M1007_d N_A_1312_126#_M1007_g N_VGND_M1032_d N_VNB_M1002_b
+ NHV L=0.5 W=0.75 AD=0.105 AS=0.173846 PD=1.03 PS=1.48718 NRD=0 NRS=5.3124 M=1
+ R=1.5 SA=250001 SB=250003 A=0.375 P=2.5 MULT=1
MM1030 N_A_2360_115#_M1030_d N_A_1212_471#_M1030_g N_A_1510_100#_M1007_d
+ N_VNB_M1002_b NHV L=0.5 W=0.75 AD=0.166635 AS=0.105 PD=1.46795 PS=1.03 NRD=0
+ NRS=0 M=1 R=1.5 SA=250001 SB=250002 A=0.375 P=2.5 MULT=1
MM1000 A_2539_181# N_A_1212_100#_M1000_g N_A_2360_115#_M1030_d N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.11235 AS=0.0933154 PD=0.955 PS=0.822051 NRD=57.6726
+ NRS=31.2132 M=1 R=0.84 SA=250003 SB=250003 A=0.21 P=1.84 MULT=1
MM1021 N_VGND_M1021_d N_A_2616_417#_M1021_g A_2539_181# N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.0609 AS=0.11235 PD=0.71 PS=0.955 NRD=0 NRS=57.6726 M=1 R=0.84
+ SA=250004 SB=250002 A=0.21 P=1.84 MULT=1
MM1025 A_2904_181# N_RESET_B_M1025_g N_VGND_M1021_d N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0609 PD=0.63 PS=0.71 NRD=13.566 NRS=2.7132 M=1 R=0.84
+ SA=250004 SB=250001 A=0.21 P=1.84 MULT=1
MM1031 N_A_2616_417#_M1031_d N_A_2360_115#_M1031_g A_2904_181# N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250005 SB=250000 A=0.21 P=1.84 MULT=1
MM1033 N_VGND_M1033_d N_CLK_M1033_g N_A_1212_100#_M1033_s N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1005 N_VGND_M1005_d N_A_2360_115#_M1005_g N_A_3417_443#_M1005_s N_VNB_M1002_b
+ NHV L=0.5 W=0.42 AD=0.0879308 AS=0.1197 PD=0.807692 PS=1.41 NRD=25.7754 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1034 N_Q_M1034_d N_A_3417_443#_M1034_g N_VGND_M1005_d N_VNB_M1002_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.157019 PD=2.03 PS=1.44231 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1008 A_222_649# N_A_116_451#_M1008_g N_A_65_649#_M1008_s N_VPB_M1008_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250000 SB=250004 A=0.21 P=1.84 MULT=1
MM1011 N_VPWR_M1011_d N_SCD_M1011_g A_222_649# N_VPB_M1008_b PHV L=0.5 W=0.42
+ AD=0.063 AS=0.0441 PD=0.72 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84 SA=250001
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1035 A_524_649# N_SCE_M1035_g N_VPWR_M1011_d N_VPB_M1008_b PHV L=0.5 W=0.42
+ AD=0.0441 AS=0.063 PD=0.63 PS=0.72 NRD=22.729 NRS=9.0916 M=1 R=0.84 SA=250002
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1037 N_A_65_649#_M1037_d N_D_M1037_g A_524_649# N_VPB_M1008_b PHV L=0.5 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84 SA=250002
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1019 N_VPWR_M1019_d N_RESET_B_M1019_g N_A_65_649#_M1037_d N_VPB_M1008_b PHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=0.99 PS=0.7 NRD=2.2729 NRS=0 M=1 R=0.84
+ SA=250003 SB=250001 A=0.21 P=1.84 MULT=1
MM1014 N_A_116_451#_M1014_d N_SCE_M1014_g N_VPWR_M1019_d N_VPB_M1008_b PHV L=0.5
+ W=0.42 AD=0.1197 AS=0.1197 PD=1.41 PS=0.99 NRD=0 NRS=129.594 M=1 R=0.84
+ SA=250004 SB=250000 A=0.21 P=1.84 MULT=1
MM1026 N_A_1312_126#_M1026_d N_A_1212_471#_M1026_g N_A_65_649#_M1026_s
+ N_VPB_M1008_b PHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1003 A_1468_641# N_A_1212_100#_M1003_g N_A_1312_126#_M1026_d N_VPB_M1008_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250001 SB=250002 A=0.21 P=1.84 MULT=1
MM1015 N_VPWR_M1015_d N_A_1510_100#_M1015_g A_1468_641# N_VPB_M1008_b PHV L=0.5
+ W=0.42 AD=0.0756 AS=0.0441 PD=0.78 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1027 N_A_1312_126#_M1027_d N_RESET_B_M1027_g N_VPWR_M1015_d N_VPB_M1008_b PHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0756 PD=1.41 PS=0.78 NRD=0 NRS=36.3664 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1020 N_VPWR_M1020_d N_A_1212_100#_M1020_g N_A_1212_471#_M1020_s N_VPB_M1008_b
+ PHV L=0.5 W=0.75 AD=0.148929 AS=0.19875 PD=1.17857 PS=2.03 NRD=36.5574 NRS=0
+ M=1 R=1.5 SA=250000 SB=250004 A=0.375 P=2.5 MULT=1
MM1009 N_A_1510_100#_M1009_d N_A_1312_126#_M1009_g N_VPWR_M1020_d N_VPB_M1008_b
+ PHV L=0.5 W=1 AD=0.14 AS=0.198571 PD=1.28 PS=1.57143 NRD=0 NRS=0 M=1 R=2
+ SA=250001 SB=250003 A=0.5 P=3 MULT=1
MM1036 N_A_2360_115#_M1036_d N_A_1212_100#_M1036_g N_A_1510_100#_M1009_d
+ N_VPB_M1008_b PHV L=0.5 W=1 AD=0.275493 AS=0.14 PD=2.0493 PS=1.28 NRD=15.2609
+ NRS=0 M=1 R=2 SA=250001 SB=250002 A=0.5 P=3 MULT=1
MM1023 A_2574_543# N_A_1212_471#_M1023_g N_A_2360_115#_M1036_d N_VPB_M1008_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.115707 PD=0.63 PS=0.860704 NRD=22.729 NRS=43.1851
+ M=1 R=0.84 SA=250003 SB=250003 A=0.21 P=1.84 MULT=1
MM1039 N_VPWR_M1039_d N_A_2616_417#_M1039_g A_2574_543# N_VPB_M1008_b PHV L=0.5
+ W=0.42 AD=0.156925 AS=0.0441 PD=1.305 PS=0.63 NRD=144.893 NRS=22.729 M=1
+ R=0.84 SA=250003 SB=250003 A=0.21 P=1.84 MULT=1
MM1006 N_A_2616_417#_M1006_d N_RESET_B_M1006_g N_VPWR_M1039_d N_VPB_M1008_b PHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.156925 PD=0.7 PS=1.305 NRD=0 NRS=144.893 M=1
+ R=0.84 SA=250004 SB=250002 A=0.21 P=1.84 MULT=1
MM1028 N_VPWR_M1028_d N_A_2360_115#_M1028_g N_A_2616_417#_M1006_d N_VPB_M1008_b
+ PHV L=0.5 W=0.42 AD=0.107638 AS=0.0588 PD=0.890256 PS=0.7 NRD=95.4809 NRS=0
+ M=1 R=0.84 SA=250005 SB=250001 A=0.21 P=1.84 MULT=1
MM1018 N_A_1212_100#_M1018_d N_CLK_M1018_g N_VPWR_M1028_d N_VPB_M1008_b PHV
+ L=0.5 W=0.75 AD=0.21375 AS=0.192212 PD=2.07 PS=1.58974 NRD=0 NRS=0 M=1 R=1.5
+ SA=250003 SB=250000 A=0.375 P=2.5 MULT=1
MM1029 N_VPWR_M1029_d N_A_2360_115#_M1029_g N_A_3417_443#_M1029_s N_VPB_M1008_b
+ PHV L=0.5 W=0.75 AD=0.17 AS=0.21375 PD=1.26333 PS=2.07 NRD=29.2803 NRS=0 M=1
+ R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1017 N_Q_M1017_d N_A_3417_443#_M1017_g N_VPWR_M1029_d N_VPB_M1008_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.34 PD=3.57 PS=2.52667 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
DX40_noxref N_VNB_M1002_b N_VPB_M1008_b NWDIODE A=51.636 P=44.92
*
.include "sky130_fd_sc_hvl__sdfrtp_1.pxi.spice"
*
.ends
*
*
