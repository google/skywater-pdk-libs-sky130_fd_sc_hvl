* File: sky130_fd_sc_hvl__o21ai_1.pxi.spice
* Created: Wed Sep  2 09:08:59 2020
* 
x_PM_SKY130_FD_SC_HVL__O21AI_1%VNB N_VNB_M1003_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__O21AI_1%VNB
x_PM_SKY130_FD_SC_HVL__O21AI_1%VPB N_VPB_M1000_b VPB N_VPB_c_27_p VPB
+ PM_SKY130_FD_SC_HVL__O21AI_1%VPB
x_PM_SKY130_FD_SC_HVL__O21AI_1%A1 N_A1_M1003_g N_A1_M1000_g A1 A1 N_A1_c_52_n
+ PM_SKY130_FD_SC_HVL__O21AI_1%A1
x_PM_SKY130_FD_SC_HVL__O21AI_1%A2 A2 A2 N_A2_M1004_g N_A2_M1001_g
+ PM_SKY130_FD_SC_HVL__O21AI_1%A2
x_PM_SKY130_FD_SC_HVL__O21AI_1%B1 N_B1_M1002_g N_B1_M1005_g B1 B1 N_B1_c_107_n
+ PM_SKY130_FD_SC_HVL__O21AI_1%B1
x_PM_SKY130_FD_SC_HVL__O21AI_1%VPWR N_VPWR_M1000_s N_VPWR_M1005_d VPWR
+ N_VPWR_c_133_n N_VPWR_c_136_n N_VPWR_c_139_n PM_SKY130_FD_SC_HVL__O21AI_1%VPWR
x_PM_SKY130_FD_SC_HVL__O21AI_1%Y N_Y_M1002_d N_Y_M1001_d N_Y_c_159_n N_Y_c_160_n
+ N_Y_c_161_n Y Y Y Y N_Y_c_163_n Y PM_SKY130_FD_SC_HVL__O21AI_1%Y
x_PM_SKY130_FD_SC_HVL__O21AI_1%A_30_107# N_A_30_107#_M1003_s N_A_30_107#_M1004_d
+ N_A_30_107#_c_195_n N_A_30_107#_c_201_n N_A_30_107#_c_197_n
+ N_A_30_107#_c_198_n PM_SKY130_FD_SC_HVL__O21AI_1%A_30_107#
x_PM_SKY130_FD_SC_HVL__O21AI_1%VGND N_VGND_M1003_d VGND N_VGND_c_225_n
+ PM_SKY130_FD_SC_HVL__O21AI_1%VGND
cc_1 N_VNB_M1003_b N_A1_M1003_g 0.0496344f $X=-0.33 $Y=-0.265 $X2=0.685 $Y2=0.91
cc_2 N_VNB_c_2_p N_A1_M1003_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.685 $Y2=0.91
cc_3 N_VNB_M1003_b N_A1_c_52_n 0.0909093f $X=-0.33 $Y=-0.265 $X2=0.69 $Y2=1.67
cc_4 N_VNB_M1003_b A2 0.0122868f $X=-0.33 $Y=-0.265 $X2=0.685 $Y2=0.91
cc_5 N_VNB_M1003_b N_A2_M1004_g 0.0828476f $X=-0.33 $Y=-0.265 $X2=0.775
+ $Y2=2.965
cc_6 N_VNB_c_2_p N_A2_M1004_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.775 $Y2=2.965
cc_7 N_VNB_M1003_b N_B1_M1002_g 0.0540153f $X=-0.33 $Y=-0.265 $X2=0.685 $Y2=0.91
cc_8 N_VNB_c_2_p N_B1_M1002_g 0.0023273f $X=0.24 $Y=0 $X2=0.685 $Y2=0.91
cc_9 N_VNB_M1003_b B1 0.0210764f $X=-0.33 $Y=-0.265 $X2=0.635 $Y2=1.58
cc_10 N_VNB_M1003_b N_B1_c_107_n 0.0621325f $X=-0.33 $Y=-0.265 $X2=0.69 $Y2=1.75
cc_11 N_VNB_M1003_b N_Y_c_159_n 0.00831213f $X=-0.33 $Y=-0.265 $X2=0.155
+ $Y2=1.58
cc_12 N_VNB_M1003_b N_Y_c_160_n 0.00176215f $X=-0.33 $Y=-0.265 $X2=0.635
+ $Y2=1.58
cc_13 N_VNB_M1003_b N_Y_c_161_n 0.044488f $X=-0.33 $Y=-0.265 $X2=0.685 $Y2=1.75
cc_14 N_VNB_c_2_p N_Y_c_161_n 8.20017e-19 $X=0.24 $Y=0 $X2=0.685 $Y2=1.75
cc_15 N_VNB_M1003_b N_Y_c_163_n 0.00211554f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_16 N_VNB_M1003_b N_A_30_107#_c_195_n 0.031352f $X=-0.33 $Y=-0.265 $X2=0.155
+ $Y2=1.58
cc_17 N_VNB_c_2_p N_A_30_107#_c_195_n 8.20017e-19 $X=0.24 $Y=0 $X2=0.155
+ $Y2=1.58
cc_18 N_VNB_M1003_b N_A_30_107#_c_197_n 0.010957f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_19 N_VNB_M1003_b N_A_30_107#_c_198_n 0.01098f $X=-0.33 $Y=-0.265 $X2=0.69
+ $Y2=1.67
cc_20 N_VNB_c_2_p N_A_30_107#_c_198_n 8.71357e-19 $X=0.24 $Y=0 $X2=0.69 $Y2=1.67
cc_21 N_VNB_M1003_b VGND 0.0957605f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_22 N_VNB_c_2_p VGND 0.359489f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_23 N_VNB_M1003_b N_VGND_c_225_n 0.0439761f $X=-0.33 $Y=-0.265 $X2=0.775
+ $Y2=2.965
cc_24 N_VNB_c_2_p N_VGND_c_225_n 0.00252795f $X=0.24 $Y=0 $X2=0.775 $Y2=2.965
cc_25 N_VPB_M1000_b N_A1_M1000_g 0.0405731f $X=-0.33 $Y=1.885 $X2=0.775
+ $Y2=2.965
cc_26 VPB N_A1_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.775 $Y2=2.965
cc_27 N_VPB_c_27_p N_A1_M1000_g 0.0137101f $X=3.12 $Y=4.07 $X2=0.775 $Y2=2.965
cc_28 N_VPB_M1000_b N_A1_c_52_n 0.0389273f $X=-0.33 $Y=1.885 $X2=0.69 $Y2=1.67
cc_29 N_VPB_M1000_b N_A2_M1004_g 0.05108f $X=-0.33 $Y=1.885 $X2=0.775 $Y2=2.965
cc_30 VPB N_A2_M1004_g 0.00970178f $X=0 $Y=3.955 $X2=0.775 $Y2=2.965
cc_31 N_VPB_c_27_p N_A2_M1004_g 0.0176589f $X=3.12 $Y=4.07 $X2=0.775 $Y2=2.965
cc_32 N_VPB_M1000_b N_B1_M1005_g 0.0410229f $X=-0.33 $Y=1.885 $X2=0.775
+ $Y2=2.965
cc_33 VPB N_B1_M1005_g 0.00970178f $X=0 $Y=3.955 $X2=0.775 $Y2=2.965
cc_34 N_VPB_c_27_p N_B1_M1005_g 0.0158814f $X=3.12 $Y=4.07 $X2=0.775 $Y2=2.965
cc_35 N_VPB_M1000_b B1 0.0214441f $X=-0.33 $Y=1.885 $X2=0.635 $Y2=1.58
cc_36 N_VPB_M1000_b N_B1_c_107_n 0.0269326f $X=-0.33 $Y=1.885 $X2=0.69 $Y2=1.75
cc_37 N_VPB_M1000_b N_VPWR_c_133_n 0.0720466f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_38 VPB N_VPWR_c_133_n 0.00377264f $X=0 $Y=3.955 $X2=0.635 $Y2=1.58
cc_39 N_VPB_c_27_p N_VPWR_c_133_n 0.0481158f $X=3.12 $Y=4.07 $X2=0.635 $Y2=1.58
cc_40 N_VPB_M1000_b N_VPWR_c_136_n 0.0771136f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_136_n 0.00341542f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_42 N_VPB_c_27_p N_VPWR_c_136_n 0.0489311f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_43 N_VPB_M1000_b N_VPWR_c_139_n 0.0483213f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_139_n 0.356745f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_45 N_VPB_c_27_p N_VPWR_c_139_n 0.0155472f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_46 N_VPB_M1000_b Y 0.00493291f $X=-0.33 $Y=1.885 $X2=0.69 $Y2=1.67
cc_47 VPB Y 0.00178441f $X=0 $Y=3.955 $X2=0.69 $Y2=1.67
cc_48 N_VPB_c_27_p Y 0.0242307f $X=3.12 $Y=4.07 $X2=0.69 $Y2=1.67
cc_49 N_VPB_M1000_b N_Y_c_163_n 5.46551e-19 $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_50 A1 A2 0.0192186f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_51 N_A1_c_52_n A2 0.00243451f $X=0.69 $Y=1.67 $X2=0 $Y2=0
cc_52 N_A1_M1003_g N_A2_M1004_g 0.0305346f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_53 A1 N_A2_M1004_g 5.64228e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_54 N_A1_c_52_n N_A2_M1004_g 0.16649f $X=0.69 $Y=1.67 $X2=0 $Y2=0
cc_55 N_A1_M1000_g N_VPWR_c_133_n 0.098289f $X=0.775 $Y=2.965 $X2=0.24 $Y2=0
cc_56 A1 N_VPWR_c_133_n 0.035216f $X=0.635 $Y=1.58 $X2=0.24 $Y2=0
cc_57 N_A1_c_52_n N_VPWR_c_133_n 0.0115742f $X=0.69 $Y=1.67 $X2=0.24 $Y2=0
cc_58 N_A1_M1000_g N_VPWR_c_139_n 0.00233065f $X=0.775 $Y=2.965 $X2=0 $Y2=0
cc_59 N_A1_M1000_g Y 0.00194962f $X=0.775 $Y=2.965 $X2=0 $Y2=0
cc_60 N_A1_c_52_n Y 4.52574e-19 $X=0.69 $Y=1.67 $X2=0 $Y2=0
cc_61 N_A1_M1003_g N_A_30_107#_c_195_n 0.0179396f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_62 N_A1_M1003_g N_A_30_107#_c_201_n 0.0274902f $X=0.685 $Y=0.91 $X2=0.24
+ $Y2=0
cc_63 A1 N_A_30_107#_c_201_n 0.0221274f $X=0.635 $Y=1.58 $X2=0.24 $Y2=0
cc_64 N_A1_c_52_n N_A_30_107#_c_201_n 0.00283794f $X=0.69 $Y=1.67 $X2=0.24 $Y2=0
cc_65 N_A1_M1003_g N_A_30_107#_c_197_n 0.00390282f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_66 A1 N_A_30_107#_c_197_n 0.0265402f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_67 N_A1_c_52_n N_A_30_107#_c_197_n 0.00856016f $X=0.69 $Y=1.67 $X2=0 $Y2=0
cc_68 N_A1_M1003_g VGND 0.0059694f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_69 N_A1_M1003_g N_VGND_c_225_n 0.0323077f $X=0.685 $Y=0.91 $X2=0 $Y2=0
cc_70 N_A2_M1004_g N_B1_M1002_g 0.0669296f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_71 A2 N_B1_c_107_n 9.3531e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_72 N_A2_M1004_g N_VPWR_c_133_n 0.0059943f $X=1.485 $Y=0.91 $X2=0.24 $Y2=0
cc_73 N_A2_M1004_g N_VPWR_c_136_n 5.02847e-19 $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_74 N_A2_M1004_g N_VPWR_c_139_n 0.0221283f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_75 A2 N_Y_c_160_n 0.010701f $X=1.595 $Y=1.58 $X2=0.24 $Y2=0
cc_76 N_A2_M1004_g N_Y_c_160_n 0.00175919f $X=1.485 $Y=0.91 $X2=0.24 $Y2=0
cc_77 A2 Y 0.0176514f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_78 N_A2_M1004_g Y 0.0707834f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_79 A2 N_Y_c_163_n 0.0108283f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_80 N_A2_M1004_g N_Y_c_163_n 0.00395465f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_81 A2 N_A_30_107#_c_201_n 0.0384286f $X=1.595 $Y=1.58 $X2=0.24 $Y2=0
cc_82 N_A2_M1004_g N_A_30_107#_c_201_n 0.0260301f $X=1.485 $Y=0.91 $X2=0.24
+ $Y2=0
cc_83 N_A2_M1004_g N_A_30_107#_c_198_n 0.0167032f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_84 N_A2_M1004_g VGND 0.005327f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_85 N_A2_M1004_g N_VGND_c_225_n 0.0320804f $X=1.485 $Y=0.91 $X2=0 $Y2=0
cc_86 N_B1_M1005_g N_VPWR_c_136_n 0.0680107f $X=2.265 $Y=2.965 $X2=0 $Y2=0
cc_87 B1 N_VPWR_c_136_n 0.0668027f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_88 N_B1_c_107_n N_VPWR_c_136_n 9.69005e-19 $X=2.49 $Y=1.89 $X2=0 $Y2=0
cc_89 N_B1_M1005_g N_VPWR_c_139_n 0.010749f $X=2.265 $Y=2.965 $X2=0 $Y2=0
cc_90 B1 N_Y_c_159_n 0.037472f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_91 N_B1_c_107_n N_Y_c_159_n 0.0378807f $X=2.49 $Y=1.89 $X2=0 $Y2=0
cc_92 N_B1_c_107_n N_Y_c_160_n 0.00854995f $X=2.49 $Y=1.89 $X2=0.24 $Y2=0
cc_93 N_B1_M1002_g N_Y_c_161_n 0.0318362f $X=2.265 $Y=0.91 $X2=0 $Y2=0
cc_94 N_B1_c_107_n N_Y_c_161_n 0.00710882f $X=2.49 $Y=1.89 $X2=0 $Y2=0
cc_95 N_B1_M1005_g Y 0.0405921f $X=2.265 $Y=2.965 $X2=0 $Y2=0
cc_96 B1 Y 4.60971e-19 $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_97 N_B1_c_107_n Y 0.00564292f $X=2.49 $Y=1.89 $X2=0 $Y2=0
cc_98 B1 N_Y_c_163_n 0.0231453f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_99 N_B1_c_107_n N_Y_c_163_n 0.0145461f $X=2.49 $Y=1.89 $X2=0 $Y2=0
cc_100 N_B1_M1002_g N_A_30_107#_c_201_n 0.00496761f $X=2.265 $Y=0.91 $X2=0.24
+ $Y2=0
cc_101 N_B1_M1002_g N_A_30_107#_c_198_n 0.0169926f $X=2.265 $Y=0.91 $X2=0 $Y2=0
cc_102 N_B1_M1002_g VGND 0.0301625f $X=2.265 $Y=0.91 $X2=0 $Y2=0
cc_103 N_B1_M1002_g N_VGND_c_225_n 8.39127e-19 $X=2.265 $Y=0.91 $X2=0 $Y2=0
cc_104 N_VPWR_c_139_n A_205_443# 0.00809061f $X=3.055 $Y=3.59 $X2=0 $Y2=3.985
cc_105 N_VPWR_c_136_n N_Y_c_159_n 0.00249128f $X=2.655 $Y=2.385 $X2=0.24
+ $Y2=4.07
cc_106 N_VPWR_c_133_n Y 0.0249574f $X=0.385 $Y=2.34 $X2=3.12 $Y2=4.07
cc_107 N_VPWR_c_136_n Y 0.108311f $X=2.655 $Y=2.385 $X2=3.12 $Y2=4.07
cc_108 N_VPWR_c_139_n Y 0.0558588f $X=3.055 $Y=3.59 $X2=3.12 $Y2=4.07
cc_109 N_Y_c_160_n N_A_30_107#_c_201_n 0.00377899f $X=2.145 $Y=1.54 $X2=0.24
+ $Y2=0
cc_110 N_Y_c_161_n N_A_30_107#_c_201_n 0.00614935f $X=2.655 $Y=0.66 $X2=0.24
+ $Y2=0
cc_111 Y N_A_30_107#_c_201_n 0.00584864f $X=1.595 $Y=1.95 $X2=0.24 $Y2=0
cc_112 N_Y_c_161_n N_A_30_107#_c_198_n 0.0187895f $X=2.655 $Y=0.66 $X2=0 $Y2=0
cc_113 N_Y_c_161_n VGND 0.0354771f $X=2.655 $Y=0.66 $X2=0 $Y2=0
cc_114 N_A_30_107#_c_201_n N_VGND_M1003_d 0.00525032f $X=1.71 $Y=1.19 $X2=0
+ $Y2=0
cc_115 N_A_30_107#_c_195_n VGND 0.0332558f $X=0.295 $Y=0.66 $X2=0 $Y2=0
cc_116 N_A_30_107#_c_201_n VGND 0.0141109f $X=1.71 $Y=1.19 $X2=0 $Y2=0
cc_117 N_A_30_107#_c_198_n VGND 0.0324443f $X=1.875 $Y=0.66 $X2=0 $Y2=0
cc_118 N_A_30_107#_c_195_n N_VGND_c_225_n 0.0307506f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_119 N_A_30_107#_c_201_n N_VGND_c_225_n 0.0540633f $X=1.71 $Y=1.19 $X2=0 $Y2=0
cc_120 N_A_30_107#_c_198_n N_VGND_c_225_n 0.0307506f $X=1.875 $Y=0.66 $X2=0
+ $Y2=0
