* File: sky130_fd_sc_hvl__a22o_1.spice
* Created: Fri Aug 28 09:32:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__a22o_1.pex.spice"
.subckt sky130_fd_sc_hvl__a22o_1  VNB VPB B2 B1 A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_83_81#_M1008_g N_X_M1008_s N_VNB_M1008_b NHV L=0.5
+ W=0.75 AD=0.4425 AS=0.19875 PD=1.93 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250004 A=0.375 P=2.5 MULT=1
MM1002 A_519_107# N_B2_M1002_g N_VGND_M1008_d N_VNB_M1008_b NHV L=0.5 W=0.75
+ AD=0.07875 AS=0.4425 PD=0.96 PS=1.93 NRD=7.5924 NRS=0 M=1 R=1.5 SA=250002
+ SB=250002 A=0.375 P=2.5 MULT=1
MM1001 N_A_83_81#_M1001_d N_B1_M1001_g A_519_107# N_VNB_M1008_b NHV L=0.5 W=0.75
+ AD=0.114375 AS=0.07875 PD=1.055 PS=0.96 NRD=3.7962 NRS=7.5924 M=1 R=1.5
+ SA=250002 SB=250002 A=0.375 P=2.5 MULT=1
MM1006 A_822_107# N_A1_M1006_g N_A_83_81#_M1001_d N_VNB_M1008_b NHV L=0.5 W=0.75
+ AD=0.07875 AS=0.114375 PD=0.96 PS=1.055 NRD=7.5924 NRS=0 M=1 R=1.5 SA=250003
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g A_822_107# N_VNB_M1008_b NHV L=0.5 W=0.75
+ AD=0.21375 AS=0.07875 PD=2.07 PS=0.96 NRD=0 NRS=7.5924 M=1 R=1.5 SA=250004
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_A_83_81#_M1009_g N_X_M1009_s N_VPB_M1009_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.4275 PD=3.57 PS=3.57 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
MM1000 N_A_83_81#_M1000_d N_B2_M1000_g N_A_316_443#_M1000_s N_VPB_M1009_b PHV
+ L=0.5 W=1.5 AD=0.21 AS=0.6675 PD=1.78 PS=3.89 NRD=0 NRS=20.3606 M=1 R=3
+ SA=250000 SB=250002 A=0.75 P=4 MULT=1
MM1004 N_A_316_443#_M1004_d N_B1_M1004_g N_A_83_81#_M1000_d N_VPB_M1009_b PHV
+ L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001
+ SB=250002 A=0.75 P=4 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_316_443#_M1004_d N_VPB_M1009_b PHV L=0.5
+ W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002 SB=250001
+ A=0.75 P=4 MULT=1
MM1005 N_A_316_443#_M1005_d N_A2_M1005_g N_VPWR_M1003_d N_VPB_M1009_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250003
+ SB=250000 A=0.75 P=4 MULT=1
DX10_noxref N_VNB_M1008_b N_VPB_M1009_b NWDIODE A=15.444 P=17.08
*
.include "sky130_fd_sc_hvl__a22o_1.pxi.spice"
*
.ends
*
*
