* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__nand2_1 A B VGND VNB VPB VPWR Y
M1000 a_233_111# B VGND VNB nhv w=750000u l=500000u
+  ad=1.575e+11p pd=1.92e+06u as=2.1375e+11p ps=2.07e+06u
M1001 Y A a_233_111# VNB nhv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
M1002 VPWR A Y VPB phv w=1.5e+06u l=500000u
+  ad=8.55e+11p pd=7.14e+06u as=4.2e+11p ps=3.56e+06u
M1003 Y B VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
