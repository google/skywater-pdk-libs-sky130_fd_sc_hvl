* NGSPICE file created from sky130_fd_sc_hvl__nand2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hvl__nand2_1 A B VGND VNB VPB VPWR Y
M1000 a_233_111# B VGND VNB nhv w=750000u l=500000u
+  ad=1.575e+11p pd=1.92e+06u as=2.1375e+11p ps=2.07e+06u
M1001 Y A a_233_111# VNB nhv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=0p ps=0u
M1002 VPWR A Y VPB phv w=1.5e+06u l=500000u
+  ad=8.55e+11p pd=7.14e+06u as=4.2e+11p ps=3.56e+06u
M1003 Y B VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends

