* File: sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3.pex.spice
* Created: Fri Aug 28 09:37:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%VNB 9 11 12 23 35 42 49
c227 9 0 3.71401e-19 $X=-0.33 $Y=-0.265
r228 29 49 6.4 $w=2.3e-07 $l=9.975e-06 $layer=MET1_cond $X=0.24 $Y=8.14
+ $X2=10.215 $Y2=8.14
r229 17 42 6.4 $w=2.3e-07 $l=9.975e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=10.215
+ $Y2=0
r230 12 35 7.85324 $w=2.3e-07 $l=1.224e-05 $layer=MET1_cond $X=12.48 $Y=8.14
+ $X2=24.72 $Y2=8.14
r231 12 49 1.45323 $w=2.3e-07 $l=2.265e-06 $layer=MET1_cond $X=12.48 $Y=8.14
+ $X2=10.215 $Y2=8.14
r232 11 23 7.85324 $w=2.3e-07 $l=1.224e-05 $layer=MET1_cond $X=12.48 $Y=0
+ $X2=24.72 $Y2=0
r233 11 42 1.45323 $w=2.3e-07 $l=2.265e-06 $layer=MET1_cond $X=12.48 $Y=0
+ $X2=10.215 $Y2=0
r234 9 35 0.357692 $w=1.7e-07 $l=4.42e-06 $layer=mcon $count=26 $X=24.72 $Y=8.14
+ $X2=24.72 $Y2=8.14
r235 9 29 0.357692 $w=1.7e-07 $l=4.42e-06 $layer=mcon $count=26 $X=0.24 $Y=8.14
+ $X2=0.24 $Y2=8.14
r236 9 23 0.357692 $w=1.7e-07 $l=4.42e-06 $layer=mcon $count=26 $X=24.72 $Y=0
+ $X2=24.72 $Y2=0
r237 9 17 0.357692 $w=1.7e-07 $l=4.42e-06 $layer=mcon $count=26 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%VPB 7 11 13 15 22 29 37
c168 13 0 2.86262e-19 $X=0 $Y=3.955
c169 7 0 5.88701e-20 $X=-0.33 $Y=1.885
r170 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.6 $Y=4.07 $X2=0.6
+ $Y2=4.07
r171 27 29 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.445 $Y=4.07
+ $X2=0.6 $Y2=4.07
r172 23 37 0.32401 $w=2.3e-07 $l=5.05e-07 $layer=MET1_cond $X=9.71 $Y=4.07
+ $X2=10.215 $Y2=4.07
r173 23 30 5.84502 $w=2.3e-07 $l=9.11e-06 $layer=MET1_cond $X=9.71 $Y=4.07
+ $X2=0.6 $Y2=4.07
r174 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.71 $Y=4.07
+ $X2=9.71 $Y2=4.07
r175 18 30 0.230978 $w=2.3e-07 $l=3.6e-07 $layer=MET1_cond $X=0.24 $Y=4.07
+ $X2=0.6 $Y2=4.07
r176 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r177 15 27 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.36 $Y=4.07
+ $X2=0.445 $Y2=4.07
r178 15 17 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.36 $Y=4.07
+ $X2=0.24 $Y2=4.07
r179 13 37 1.45323 $w=2.3e-07 $l=2.265e-06 $layer=MET1_cond $X=12.48 $Y=4.07
+ $X2=10.215 $Y2=4.07
r180 9 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.445 $Y=4.155
+ $X2=0.445 $Y2=4.07
r181 9 11 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=0.445 $Y=4.155
+ $X2=0.445 $Y2=4.875
r182 7 22 91 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=9.135 $Y=3.985 $X2=9.71 $Y2=4.07
r183 7 17 182 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=1 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
r184 7 11 182 $w=1.7e-07 $l=1.09002e-06 $layer=licon1_NTAP_notbjt $count=1 $X=0
+ $Y=3.985 $X2=0.445 $Y2=4.875
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%LVPWR 1 2 3 4 5 6 7 8 28
+ 32 34 40 44 45 46 47 50 54 56 58 60 63 67 69 73 77 78 80 83 87 92
c193 78 0 1.46493e-19 $X=18.88 $Y=3.62
c194 77 0 1.39769e-19 $X=18.85 $Y=4.52
r195 89 90 7.36913 $w=7.45e-07 $l=4.5e-07 $layer=LI1_cond $X=20.042 $Y=4.07
+ $X2=20.042 $Y2=4.52
r196 88 89 7.36913 $w=7.45e-07 $l=4.5e-07 $layer=LI1_cond $X=20.042 $Y=3.62
+ $X2=20.042 $Y2=4.07
r197 86 88 7.61477 $w=7.45e-07 $l=4.65e-07 $layer=LI1_cond $X=20.042 $Y=3.155
+ $X2=20.042 $Y2=3.62
r198 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.245 $Y=3.155
+ $X2=20.245 $Y2=3.155
r199 83 87 3.8701 $w=2.85e-07 $l=7.765e-06 $layer=MET1_cond $X=12.48 $Y=3.162
+ $X2=20.245 $Y2=3.162
r200 83 92 1.12888 $w=2.85e-07 $l=2.265e-06 $layer=MET1_cond $X=12.48 $Y=3.162
+ $X2=10.215 $Y2=3.162
r201 80 82 2.5376 $w=6.25e-07 $l=1.3e-07 $layer=LI1_cond $X=20.042 $Y=5.64
+ $X2=20.042 $Y2=5.77
r202 73 75 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=21.235 $Y=4.94
+ $X2=21.235 $Y2=5.64
r203 71 73 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=21.235 $Y=4.605
+ $X2=21.235 $Y2=4.94
r204 70 90 9.73363 $w=1.7e-07 $l=3.78e-07 $layer=LI1_cond $X=20.42 $Y=4.52
+ $X2=20.042 $Y2=4.52
r205 69 71 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=21.07 $Y=4.52
+ $X2=21.235 $Y2=4.605
r206 69 70 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=21.07 $Y=4.52
+ $X2=20.42 $Y2=4.52
r207 65 86 7.98612 $w=7.45e-07 $l=2.81521e-07 $layer=LI1_cond $X=19.82 $Y=3.02
+ $X2=20.042 $Y2=3.155
r208 65 67 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=19.82 $Y=3.02
+ $X2=19.82 $Y2=2.84
r209 61 80 3.82348 $w=7.55e-07 $l=2.12e-07 $layer=LI1_cond $X=20.042 $Y=5.428
+ $X2=20.042 $Y2=5.64
r210 61 63 7.73094 $w=7.53e-07 $l=4.88e-07 $layer=LI1_cond $X=20.042 $Y=5.428
+ $X2=20.042 $Y2=4.94
r211 60 90 1.37351 $w=7.55e-07 $l=8.5e-08 $layer=LI1_cond $X=20.042 $Y=4.605
+ $X2=20.042 $Y2=4.52
r212 60 63 5.3071 $w=7.53e-07 $l=3.35e-07 $layer=LI1_cond $X=20.042 $Y=4.605
+ $X2=20.042 $Y2=4.94
r213 59 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.965 $Y=3.62
+ $X2=18.88 $Y2=3.62
r214 58 88 9.73363 $w=1.7e-07 $l=3.77e-07 $layer=LI1_cond $X=19.665 $Y=3.62
+ $X2=20.042 $Y2=3.62
r215 58 59 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=19.665 $Y=3.62
+ $X2=18.965 $Y2=3.62
r216 57 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.935 $Y=4.52
+ $X2=18.85 $Y2=4.52
r217 56 90 9.73363 $w=1.7e-07 $l=3.77e-07 $layer=LI1_cond $X=19.665 $Y=4.52
+ $X2=20.042 $Y2=4.52
r218 56 57 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=19.665 $Y=4.52
+ $X2=18.935 $Y2=4.52
r219 52 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.88 $Y=3.535
+ $X2=18.88 $Y2=3.62
r220 52 54 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=18.88 $Y=3.535
+ $X2=18.88 $Y2=2.84
r221 48 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.85 $Y=4.605
+ $X2=18.85 $Y2=4.52
r222 48 50 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=18.85 $Y=4.605
+ $X2=18.85 $Y2=4.94
r223 46 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.795 $Y=3.62
+ $X2=18.88 $Y2=3.62
r224 46 47 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=18.795 $Y=3.62
+ $X2=18.065 $Y2=3.62
r225 44 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.765 $Y=4.52
+ $X2=18.85 $Y2=4.52
r226 44 45 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=18.765 $Y=4.52
+ $X2=18.035 $Y2=4.52
r227 40 43 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=17.94 $Y=2.5
+ $X2=17.94 $Y2=3.2
r228 38 47 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=17.94 $Y=3.535
+ $X2=18.065 $Y2=3.62
r229 38 43 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=17.94 $Y=3.535
+ $X2=17.94 $Y2=3.2
r230 34 89 5.52765 $w=3.3e-07 $l=3.77e-07 $layer=LI1_cond $X=19.665 $Y=4.07
+ $X2=20.042 $Y2=4.07
r231 34 36 44.5262 $w=3.28e-07 $l=1.275e-06 $layer=LI1_cond $X=19.665 $Y=4.07
+ $X2=18.39 $Y2=4.07
r232 30 45 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=17.91 $Y=4.605
+ $X2=18.035 $Y2=4.52
r233 30 32 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=17.91 $Y=4.605
+ $X2=17.91 $Y2=4.94
r234 28 36 91 $w=1.7e-07 $l=6.36082e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=17.795 $Y=3.985 $X2=18.39 $Y2=4.07
r235 8 75 400 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=21.085
+ $Y=4.795 $X2=21.235 $Y2=5.64
r236 8 73 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=21.085
+ $Y=4.795 $X2=21.235 $Y2=4.94
r237 7 82 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=20.2
+ $Y=4.795 $X2=20.335 $Y2=5.77
r238 7 63 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=20.2
+ $Y=4.795 $X2=20.335 $Y2=4.94
r239 6 67 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=19.63
+ $Y=2.225 $X2=19.78 $Y2=2.84
r240 5 80 400 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=19.6
+ $Y=4.795 $X2=19.75 $Y2=5.64
r241 5 63 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=19.6
+ $Y=4.795 $X2=19.75 $Y2=4.94
r242 4 54 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=18.73
+ $Y=2.225 $X2=18.88 $Y2=2.84
r243 3 50 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=18.7
+ $Y=4.795 $X2=18.85 $Y2=4.94
r244 2 43 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=17.835
+ $Y=2.225 $X2=17.98 $Y2=3.2
r245 2 40 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=17.835
+ $Y=2.225 $X2=17.98 $Y2=2.5
r246 1 32 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=17.805
+ $Y=4.795 $X2=17.95 $Y2=4.94
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%VGND 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 60 64 67 70 71 73 75 81 86 87 89 95 101 107 113 119
+ 125 129 131 133 135 137 139 141 145 149 151 153 155 157 161 163 167 169 171
+ 173 175 176 178 179 181 182 184 185 187 188 190 191 193 194 195 196 197 198
+ 199 200 201 213 222 269 280 283 291 307
c251 13 0 7.44113e-20 $X=17.8 $Y=6.645
r252 282 283 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=21.265 $Y=7.63
+ $X2=21.265 $Y2=7.63
r253 279 280 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=19.825 $Y=0.51
+ $X2=19.825 $Y2=0.51
r254 277 283 1.28992 $w=3.7e-07 $l=3.36e-06 $layer=MET1_cond $X=17.905 $Y=7.7
+ $X2=21.265 $Y2=7.7
r255 276 277 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=17.905 $Y=7.63
+ $X2=17.905 $Y2=7.63
r256 274 280 0.737098 $w=3.7e-07 $l=1.92e-06 $layer=MET1_cond $X=17.905 $Y=0.44
+ $X2=19.825 $Y2=0.44
r257 273 274 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=17.905 $Y=0.51
+ $X2=17.905 $Y2=0.51
r258 270 291 1.99439 $w=3.7e-07 $l=5.195e-06 $layer=MET1_cond $X=5.02 $Y=0.44
+ $X2=10.215 $Y2=0.44
r259 269 270 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.02 $Y=0.37
+ $X2=5.02 $Y2=0.37
r260 266 269 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=4.84 $Y=0.37
+ $X2=5.02 $Y2=0.37
r261 265 270 0.579697 $w=3.7e-07 $l=1.51e-06 $layer=MET1_cond $X=3.51 $Y=0.44
+ $X2=5.02 $Y2=0.44
r262 264 265 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.51 $Y=0.37
+ $X2=3.51 $Y2=0.37
r263 261 262 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.95 $Y=0.37
+ $X2=1.95 $Y2=0.37
r264 258 259 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=7.685
+ $X2=1.2 $Y2=7.685
r265 256 277 1.25345 $w=3.7e-07 $l=3.265e-06 $layer=MET1_cond $X=14.64 $Y=7.7
+ $X2=17.905 $Y2=7.7
r266 255 256 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.64 $Y=7.685
+ $X2=14.64 $Y2=7.685
r267 253 256 0.370469 $w=3.7e-07 $l=9.65e-07 $layer=MET1_cond $X=13.675 $Y=7.7
+ $X2=14.64 $Y2=7.7
r268 252 255 48.3525 $w=2.28e-07 $l=9.65e-07 $layer=LI1_cond $X=13.675 $Y=7.685
+ $X2=14.64 $Y2=7.685
r269 252 253 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.675 $Y=7.685
+ $X2=13.675 $Y2=7.685
r270 250 253 0.182355 $w=3.7e-07 $l=4.75e-07 $layer=MET1_cond $X=13.2 $Y=7.7
+ $X2=13.675 $Y2=7.7
r271 249 250 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=7.685
+ $X2=13.2 $Y2=7.685
r272 246 249 48.102 $w=2.28e-07 $l=9.6e-07 $layer=LI1_cond $X=12.24 $Y=7.685
+ $X2=13.2 $Y2=7.685
r273 246 247 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=7.685
+ $X2=12.24 $Y2=7.685
r274 244 247 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=7.7
+ $X2=12.24 $Y2=7.7
r275 244 307 0.489479 $w=3.7e-07 $l=1.275e-06 $layer=MET1_cond $X=11.76 $Y=7.7
+ $X2=10.485 $Y2=7.7
r276 243 244 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.76 $Y=7.685
+ $X2=11.76 $Y2=7.685
r277 241 307 0.247619 $w=3.7e-07 $l=6.45e-07 $layer=MET1_cond $X=9.84 $Y=7.7
+ $X2=10.485 $Y2=7.7
r278 240 243 96.2039 $w=2.28e-07 $l=1.92e-06 $layer=LI1_cond $X=9.84 $Y=7.685
+ $X2=11.76 $Y2=7.685
r279 240 241 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=7.685
+ $X2=9.84 $Y2=7.685
r280 238 241 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=7.7
+ $X2=9.84 $Y2=7.7
r281 237 238 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=7.685
+ $X2=9.36 $Y2=7.685
r282 235 238 0.737098 $w=3.7e-07 $l=1.92e-06 $layer=MET1_cond $X=7.44 $Y=7.7
+ $X2=9.36 $Y2=7.7
r283 234 237 96.2039 $w=2.28e-07 $l=1.92e-06 $layer=LI1_cond $X=7.44 $Y=7.685
+ $X2=9.36 $Y2=7.685
r284 234 235 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=7.685
+ $X2=7.44 $Y2=7.685
r285 232 235 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=7.7
+ $X2=7.44 $Y2=7.7
r286 231 232 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=7.685
+ $X2=6.96 $Y2=7.685
r287 229 232 0.737098 $w=3.7e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=7.7
+ $X2=6.96 $Y2=7.7
r288 228 231 96.2039 $w=2.28e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=7.685
+ $X2=6.96 $Y2=7.685
r289 228 229 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=7.685
+ $X2=5.04 $Y2=7.685
r290 225 265 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=3.15 $Y=0.44
+ $X2=3.51 $Y2=0.44
r291 224 225 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.15 $Y=0.37
+ $X2=3.15 $Y2=0.37
r292 222 264 3.40825 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=3.395 $Y=0.37
+ $X2=3.51 $Y2=0.37
r293 222 224 12.276 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.395 $Y=0.37
+ $X2=3.15 $Y2=0.37
r294 221 229 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=7.7
+ $X2=5.04 $Y2=7.7
r295 220 221 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=7.685
+ $X2=4.56 $Y2=7.685
r296 218 221 0.737098 $w=3.7e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=7.7
+ $X2=4.56 $Y2=7.7
r297 217 220 96.2039 $w=2.28e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=7.685
+ $X2=4.56 $Y2=7.685
r298 217 218 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=7.685
+ $X2=2.64 $Y2=7.685
r299 214 225 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=2.31 $Y=0.44
+ $X2=3.15 $Y2=0.44
r300 214 262 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=2.31 $Y=0.44
+ $X2=1.95 $Y2=0.44
r301 213 214 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.31 $Y=0.37
+ $X2=2.31 $Y2=0.37
r302 211 261 3.40825 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=2.065 $Y=0.37
+ $X2=1.95 $Y2=0.37
r303 211 213 12.276 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.065 $Y=0.37
+ $X2=2.31 $Y2=0.37
r304 210 218 0.184275 $w=3.7e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=7.7
+ $X2=2.64 $Y2=7.7
r305 210 259 0.368549 $w=3.7e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=7.7
+ $X2=1.2 $Y2=7.7
r306 209 210 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=7.685
+ $X2=2.16 $Y2=7.685
r307 207 258 3.33465 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=1.28 $Y=7.685
+ $X2=1.17 $Y2=7.685
r308 207 209 44.0935 $w=2.28e-07 $l=8.8e-07 $layer=LI1_cond $X=1.28 $Y=7.685
+ $X2=2.16 $Y2=7.685
r309 201 250 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=12.48 $Y=7.7
+ $X2=13.2 $Y2=7.7
r310 201 247 0.0921373 $w=3.7e-07 $l=2.4e-07 $layer=MET1_cond $X=12.48 $Y=7.7
+ $X2=12.24 $Y2=7.7
r311 200 274 2.08269 $w=3.7e-07 $l=5.425e-06 $layer=MET1_cond $X=12.48 $Y=0.44
+ $X2=17.905 $Y2=0.44
r312 200 291 0.869546 $w=3.7e-07 $l=2.265e-06 $layer=MET1_cond $X=12.48 $Y=0.44
+ $X2=10.215 $Y2=0.44
r313 195 255 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=14.665 $Y=7.685
+ $X2=14.64 $Y2=7.685
r314 193 249 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=13.335 $Y=7.685
+ $X2=13.2 $Y2=7.685
r315 193 194 4.97762 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=13.335 $Y=7.685
+ $X2=13.445 $Y2=7.685
r316 192 252 6.01275 $w=2.28e-07 $l=1.2e-07 $layer=LI1_cond $X=13.555 $Y=7.685
+ $X2=13.675 $Y2=7.685
r317 192 194 4.97762 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=13.555 $Y=7.685
+ $X2=13.445 $Y2=7.685
r318 190 243 3.50744 $w=2.28e-07 $l=7e-08 $layer=LI1_cond $X=11.83 $Y=7.685
+ $X2=11.76 $Y2=7.685
r319 190 191 4.97762 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=11.83 $Y=7.685
+ $X2=11.94 $Y2=7.685
r320 189 246 9.52018 $w=2.28e-07 $l=1.9e-07 $layer=LI1_cond $X=12.05 $Y=7.685
+ $X2=12.24 $Y2=7.685
r321 189 191 4.97762 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=12.05 $Y=7.685
+ $X2=11.94 $Y2=7.685
r322 187 237 5.51168 $w=2.28e-07 $l=1.1e-07 $layer=LI1_cond $X=9.47 $Y=7.685
+ $X2=9.36 $Y2=7.685
r323 187 188 4.97762 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=9.47 $Y=7.685
+ $X2=9.58 $Y2=7.685
r324 186 240 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=9.69 $Y=7.685
+ $X2=9.84 $Y2=7.685
r325 186 188 4.97762 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=9.69 $Y=7.685
+ $X2=9.58 $Y2=7.685
r326 184 231 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=7.11 $Y=7.685
+ $X2=6.96 $Y2=7.685
r327 184 185 4.97762 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=7.11 $Y=7.685
+ $X2=7.22 $Y2=7.685
r328 183 234 5.51168 $w=2.28e-07 $l=1.1e-07 $layer=LI1_cond $X=7.33 $Y=7.685
+ $X2=7.44 $Y2=7.685
r329 183 185 4.97762 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=7.33 $Y=7.685
+ $X2=7.22 $Y2=7.685
r330 181 220 9.52018 $w=2.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.75 $Y=7.685
+ $X2=4.56 $Y2=7.685
r331 181 182 4.97762 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.75 $Y=7.685
+ $X2=4.86 $Y2=7.685
r332 180 228 3.50744 $w=2.28e-07 $l=7e-08 $layer=LI1_cond $X=4.97 $Y=7.685
+ $X2=5.04 $Y2=7.685
r333 180 182 4.97762 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.97 $Y=7.685
+ $X2=4.86 $Y2=7.685
r334 178 209 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=7.685
+ $X2=2.16 $Y2=7.685
r335 178 179 4.97762 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=2.36 $Y=7.685
+ $X2=2.47 $Y2=7.685
r336 177 217 3.00637 $w=2.28e-07 $l=6e-08 $layer=LI1_cond $X=2.58 $Y=7.685
+ $X2=2.64 $Y2=7.685
r337 177 179 4.97762 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=2.58 $Y=7.685
+ $X2=2.47 $Y2=7.685
r338 171 282 3.27362 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=21.25 $Y=7.515
+ $X2=21.25 $Y2=7.63
r339 171 173 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=21.25 $Y=7.515
+ $X2=21.25 $Y2=6.79
r340 170 199 5.53409 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=20.435 $Y=7.63
+ $X2=20.31 $Y2=7.63
r341 169 282 3.55828 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=21.125 $Y=7.63
+ $X2=21.25 $Y2=7.63
r342 169 170 34.5733 $w=2.28e-07 $l=6.9e-07 $layer=LI1_cond $X=21.125 $Y=7.63
+ $X2=20.435 $Y2=7.63
r343 165 199 1.04409 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=20.31 $Y=7.515
+ $X2=20.31 $Y2=7.63
r344 165 167 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=20.31 $Y=7.515
+ $X2=20.31 $Y2=6.79
r345 164 198 6.89714 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=19.95 $Y=7.63
+ $X2=19.785 $Y2=7.63
r346 163 199 5.53409 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=20.185 $Y=7.63
+ $X2=20.31 $Y2=7.63
r347 163 164 11.775 $w=2.28e-07 $l=2.35e-07 $layer=LI1_cond $X=20.185 $Y=7.63
+ $X2=19.95 $Y2=7.63
r348 159 198 0.0811015 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=19.785 $Y=7.515
+ $X2=19.785 $Y2=7.63
r349 159 161 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=19.785 $Y=7.515
+ $X2=19.785 $Y2=6.79
r350 155 279 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=19.785 $Y=0.625
+ $X2=19.785 $Y2=0.51
r351 155 157 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=19.785 $Y=0.625
+ $X2=19.785 $Y2=0.98
r352 154 197 6.89714 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=19.04 $Y=0.51
+ $X2=18.875 $Y2=0.51
r353 153 279 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=19.62 $Y=0.51
+ $X2=19.785 $Y2=0.51
r354 153 154 29.0616 $w=2.28e-07 $l=5.8e-07 $layer=LI1_cond $X=19.62 $Y=0.51
+ $X2=19.04 $Y2=0.51
r355 152 196 6.89714 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=19.02 $Y=7.63
+ $X2=18.855 $Y2=7.63
r356 151 198 6.89714 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=19.62 $Y=7.63
+ $X2=19.785 $Y2=7.63
r357 151 152 30.0637 $w=2.28e-07 $l=6e-07 $layer=LI1_cond $X=19.62 $Y=7.63
+ $X2=19.02 $Y2=7.63
r358 147 197 0.0811015 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=18.875 $Y=0.625
+ $X2=18.875 $Y2=0.51
r359 147 149 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=18.875 $Y=0.625
+ $X2=18.875 $Y2=0.98
r360 143 196 0.0811015 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=18.855 $Y=7.515
+ $X2=18.855 $Y2=7.63
r361 143 145 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=18.855 $Y=7.515
+ $X2=18.855 $Y2=7.16
r362 142 276 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=18.11 $Y=7.63
+ $X2=17.945 $Y2=7.63
r363 141 196 6.89714 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=18.69 $Y=7.63
+ $X2=18.855 $Y2=7.63
r364 141 142 29.0616 $w=2.28e-07 $l=5.8e-07 $layer=LI1_cond $X=18.69 $Y=7.63
+ $X2=18.11 $Y2=7.63
r365 140 273 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=18.11 $Y=0.51
+ $X2=17.945 $Y2=0.51
r366 139 197 6.89714 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=18.71 $Y=0.51
+ $X2=18.875 $Y2=0.51
r367 139 140 30.0637 $w=2.28e-07 $l=6e-07 $layer=LI1_cond $X=18.71 $Y=0.51
+ $X2=18.11 $Y2=0.51
r368 135 276 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=17.945 $Y=7.515
+ $X2=17.945 $Y2=7.63
r369 135 137 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=17.945 $Y=7.515
+ $X2=17.945 $Y2=7.16
r370 131 273 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=17.945 $Y=0.625
+ $X2=17.945 $Y2=0.51
r371 131 133 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=17.945 $Y=0.625
+ $X2=17.945 $Y2=0.9
r372 127 195 6.82087 $w=2.3e-07 $l=1.60857e-07 $layer=LI1_cond $X=14.775 $Y=7.57
+ $X2=14.665 $Y2=7.685
r373 127 129 63.3844 $w=2.18e-07 $l=1.21e-06 $layer=LI1_cond $X=14.775 $Y=7.57
+ $X2=14.775 $Y2=6.36
r374 123 194 1.50311 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=13.445 $Y=7.57
+ $X2=13.445 $Y2=7.685
r375 123 125 63.3844 $w=2.18e-07 $l=1.21e-06 $layer=LI1_cond $X=13.445 $Y=7.57
+ $X2=13.445 $Y2=6.36
r376 119 122 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=11.94 $Y=6.36
+ $X2=11.94 $Y2=7.04
r377 117 191 1.50311 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=11.94 $Y=7.57
+ $X2=11.94 $Y2=7.685
r378 117 122 27.7634 $w=2.18e-07 $l=5.3e-07 $layer=LI1_cond $X=11.94 $Y=7.57
+ $X2=11.94 $Y2=7.04
r379 113 116 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=9.58 $Y=6.36
+ $X2=9.58 $Y2=7.04
r380 111 188 1.50311 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=9.58 $Y=7.57
+ $X2=9.58 $Y2=7.685
r381 111 116 27.7634 $w=2.18e-07 $l=5.3e-07 $layer=LI1_cond $X=9.58 $Y=7.57
+ $X2=9.58 $Y2=7.04
r382 107 110 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=7.22 $Y=6.36
+ $X2=7.22 $Y2=7.04
r383 105 185 1.50311 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=7.22 $Y=7.57
+ $X2=7.22 $Y2=7.685
r384 105 110 27.7634 $w=2.18e-07 $l=5.3e-07 $layer=LI1_cond $X=7.22 $Y=7.57
+ $X2=7.22 $Y2=7.04
r385 101 104 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=4.86 $Y=6.36
+ $X2=4.86 $Y2=7.04
r386 99 182 1.50311 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=4.86 $Y=7.57
+ $X2=4.86 $Y2=7.685
r387 99 104 27.7634 $w=2.18e-07 $l=5.3e-07 $layer=LI1_cond $X=4.86 $Y=7.57
+ $X2=4.86 $Y2=7.04
r388 95 97 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.84 $Y=0.81
+ $X2=4.84 $Y2=1.49
r389 93 266 0.716491 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=4.84 $Y=0.485
+ $X2=4.84 $Y2=0.37
r390 93 95 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.84 $Y=0.485
+ $X2=4.84 $Y2=0.81
r391 89 91 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.51 $Y=0.81
+ $X2=3.51 $Y2=1.49
r392 87 264 3.40825 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=3.51 $Y=0.485
+ $X2=3.51 $Y2=0.37
r393 87 89 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.51 $Y=0.485
+ $X2=3.51 $Y2=0.81
r394 86 179 1.50311 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=2.47 $Y=7.57
+ $X2=2.47 $Y2=7.685
r395 86 176 19.1201 $w=2.18e-07 $l=3.65e-07 $layer=LI1_cond $X=2.47 $Y=7.57
+ $X2=2.47 $Y2=7.205
r396 81 84 34.8294 $w=2.23e-07 $l=6.8e-07 $layer=LI1_cond $X=2.472 $Y=6.36
+ $X2=2.472 $Y2=7.04
r397 79 176 5.73661 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=2.472 $Y=7.093
+ $X2=2.472 $Y2=7.205
r398 79 84 2.71464 $w=2.23e-07 $l=5.3e-08 $layer=LI1_cond $X=2.472 $Y=7.093
+ $X2=2.472 $Y2=7.04
r399 75 77 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.95 $Y=0.81
+ $X2=1.95 $Y2=1.49
r400 73 261 3.40825 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=1.95 $Y=0.485
+ $X2=1.95 $Y2=0.37
r401 73 75 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.95 $Y=0.485
+ $X2=1.95 $Y2=0.81
r402 71 205 16.2827 $w=6.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=7.015
+ $X2=1.465 $Y2=6.85
r403 70 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.625
+ $Y=7.015 $X2=1.625 $Y2=7.015
r404 68 175 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=1.28 $Y=7.015
+ $X2=1.17 $Y2=7.015
r405 68 70 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.28 $Y=7.015
+ $X2=1.625 $Y2=7.015
r406 67 258 3.48622 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=1.17 $Y=7.57
+ $X2=1.17 $Y2=7.685
r407 66 175 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.17 $Y=7.18
+ $X2=1.17 $Y2=7.015
r408 66 67 20.4297 $w=2.18e-07 $l=3.9e-07 $layer=LI1_cond $X=1.17 $Y=7.18
+ $X2=1.17 $Y2=7.57
r409 62 175 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.17 $Y=6.85
+ $X2=1.17 $Y2=7.015
r410 62 64 25.668 $w=2.18e-07 $l=4.9e-07 $layer=LI1_cond $X=1.17 $Y=6.85
+ $X2=1.17 $Y2=6.36
r411 60 205 45.4775 $w=5e-07 $l=4.25e-07 $layer=POLY_cond $X=1.56 $Y=6.425
+ $X2=1.56 $Y2=6.85
r412 19 173 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=21.07
+ $Y=6.645 $X2=21.21 $Y2=6.79
r413 18 167 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=20.205
+ $Y=6.645 $X2=20.35 $Y2=6.79
r414 17 157 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=19.645
+ $Y=0.755 $X2=19.785 $Y2=0.98
r415 16 161 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=19.615
+ $Y=6.645 $X2=19.785 $Y2=6.79
r416 15 149 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=18.735
+ $Y=0.755 $X2=18.875 $Y2=0.98
r417 14 145 182 $w=1.7e-07 $l=6.02557e-07 $layer=licon1_NDIFF $count=1 $X=18.665
+ $Y=6.645 $X2=18.855 $Y2=7.16
r418 13 137 182 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_NDIFF $count=1 $X=17.8
+ $Y=6.645 $X2=17.945 $Y2=7.16
r419 12 133 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=17.8
+ $Y=0.755 $X2=17.945 $Y2=0.9
r420 11 129 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.635
+ $Y=6.215 $X2=14.775 $Y2=6.36
r421 10 125 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=13.305
+ $Y=6.215 $X2=13.445 $Y2=6.36
r422 9 122 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1
+ $X=11.8 $Y=6.215 $X2=11.94 $Y2=7.04
r423 9 119 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1
+ $X=11.8 $Y=6.215 $X2=11.94 $Y2=6.36
r424 8 116 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1
+ $X=9.44 $Y=6.215 $X2=9.58 $Y2=7.04
r425 8 113 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1
+ $X=9.44 $Y=6.215 $X2=9.58 $Y2=6.36
r426 7 110 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1
+ $X=7.08 $Y=6.215 $X2=7.22 $Y2=7.04
r427 7 107 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1
+ $X=7.08 $Y=6.215 $X2=7.22 $Y2=6.36
r428 6 104 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1
+ $X=4.72 $Y=6.215 $X2=4.86 $Y2=7.04
r429 6 101 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1
+ $X=4.72 $Y=6.215 $X2=4.86 $Y2=6.36
r430 5 97 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1 $X=4.7
+ $Y=0.665 $X2=4.84 $Y2=1.49
r431 5 95 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.7
+ $Y=0.665 $X2=4.84 $Y2=0.81
r432 4 91 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1 $X=3.37
+ $Y=0.665 $X2=3.51 $Y2=1.49
r433 4 89 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.37
+ $Y=0.665 $X2=3.51 $Y2=0.81
r434 3 84 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1
+ $X=2.375 $Y=6.215 $X2=2.5 $Y2=7.04
r435 3 81 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1
+ $X=2.375 $Y=6.215 $X2=2.5 $Y2=6.36
r436 2 77 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1 $X=1.81
+ $Y=0.665 $X2=1.95 $Y2=1.49
r437 2 75 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.81
+ $Y=0.665 $X2=1.95 $Y2=0.81
r438 1 64 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=6.215 $X2=1.17 $Y2=6.36
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_262_107# 1 2 3 4 15 19
+ 21 25 29 31 35 39 41 42 43 46 50 56 60 64 70 74 75
r126 70 72 53.4314 $w=2.18e-07 $l=1.02e-06 $layer=LI1_cond $X=5.62 $Y=2.57
+ $X2=5.62 $Y2=3.59
r127 68 75 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=5.62 $Y=2.14
+ $X2=5.62 $Y2=2.03
r128 68 70 22.525 $w=2.18e-07 $l=4.3e-07 $layer=LI1_cond $X=5.62 $Y=2.14
+ $X2=5.62 $Y2=2.57
r129 64 67 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=5.62 $Y=0.81
+ $X2=5.62 $Y2=1.49
r130 62 75 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=5.62 $Y=1.92
+ $X2=5.62 $Y2=2.03
r131 62 67 22.525 $w=2.18e-07 $l=4.3e-07 $layer=LI1_cond $X=5.62 $Y=1.92
+ $X2=5.62 $Y2=1.49
r132 61 74 2.39845 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.17 $Y=2.03
+ $X2=4.06 $Y2=2.03
r133 60 75 1.34256 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=5.51 $Y=2.03
+ $X2=5.62 $Y2=2.03
r134 60 61 70.1943 $w=2.18e-07 $l=1.34e-06 $layer=LI1_cond $X=5.51 $Y=2.03
+ $X2=4.17 $Y2=2.03
r135 56 58 53.4314 $w=2.18e-07 $l=1.02e-06 $layer=LI1_cond $X=4.06 $Y=2.57
+ $X2=4.06 $Y2=3.59
r136 54 74 3.75657 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=2.195
+ $X2=4.06 $Y2=2.03
r137 54 56 19.6439 $w=2.18e-07 $l=3.75e-07 $layer=LI1_cond $X=4.06 $Y=2.195
+ $X2=4.06 $Y2=2.57
r138 50 53 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=4.06 $Y=0.81
+ $X2=4.06 $Y2=1.49
r139 48 74 3.75657 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=1.865
+ $X2=4.06 $Y2=2.03
r140 48 53 19.6439 $w=2.18e-07 $l=3.75e-07 $layer=LI1_cond $X=4.06 $Y=1.865
+ $X2=4.06 $Y2=1.49
r141 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.515
+ $Y=2.03 $X2=3.515 $Y2=2.03
r142 43 74 2.39845 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=3.95 $Y=2.03
+ $X2=4.06 $Y2=2.03
r143 43 45 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=3.95 $Y=2.03
+ $X2=3.515 $Y2=2.03
r144 33 46 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=3.12 $Y=2.03
+ $X2=3.515 $Y2=2.03
r145 33 39 185.12 $w=5e-07 $l=1.73e-06 $layer=POLY_cond $X=3.12 $Y=2.195
+ $X2=3.12 $Y2=3.925
r146 33 35 74.9041 $w=5e-07 $l=7e-07 $layer=POLY_cond $X=3.12 $Y=1.865 $X2=3.12
+ $Y2=1.165
r147 32 42 60.25 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=2.59 $Y=2.03 $X2=2.34
+ $Y2=2.03
r148 31 33 52.6045 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=2.87 $Y=2.03
+ $X2=3.12 $Y2=2.03
r149 31 32 92.8416 $w=2e-07 $l=2.8e-07 $layer=POLY_cond $X=2.87 $Y=2.03 $X2=2.59
+ $Y2=2.03
r150 27 42 9.64 $w=5e-07 $l=1e-07 $layer=POLY_cond $X=2.34 $Y=2.13 $X2=2.34
+ $Y2=2.03
r151 27 29 192.076 $w=5e-07 $l=1.795e-06 $layer=POLY_cond $X=2.34 $Y=2.13
+ $X2=2.34 $Y2=3.925
r152 23 42 9.64 $w=5e-07 $l=1e-07 $layer=POLY_cond $X=2.34 $Y=1.93 $X2=2.34
+ $Y2=2.03
r153 23 25 81.8595 $w=5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.34 $Y=1.93
+ $X2=2.34 $Y2=1.165
r154 22 41 18.8672 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=1.81 $Y=2.03 $X2=1.56
+ $Y2=2.03
r155 21 42 60.25 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=2.09 $Y=2.03 $X2=2.34
+ $Y2=2.03
r156 21 22 92.8416 $w=2e-07 $l=2.8e-07 $layer=POLY_cond $X=2.09 $Y=2.03 $X2=1.81
+ $Y2=2.03
r157 17 41 9.03033 $w=5e-07 $l=1e-07 $layer=POLY_cond $X=1.56 $Y=2.13 $X2=1.56
+ $Y2=2.03
r158 17 19 192.076 $w=5e-07 $l=1.795e-06 $layer=POLY_cond $X=1.56 $Y=2.13
+ $X2=1.56 $Y2=3.925
r159 13 41 9.03033 $w=5e-07 $l=1e-07 $layer=POLY_cond $X=1.56 $Y=1.93 $X2=1.56
+ $Y2=2.03
r160 13 15 81.8595 $w=5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.56 $Y=1.93
+ $X2=1.56 $Y2=1.165
r161 4 72 300 $w=1.7e-07 $l=1.23301e-06 $layer=licon1_PDIFF $count=2 $X=5.48
+ $Y=2.425 $X2=5.62 $Y2=3.59
r162 4 70 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=5.48
+ $Y=2.425 $X2=5.62 $Y2=2.57
r163 3 58 300 $w=1.7e-07 $l=1.22591e-06 $layer=licon1_PDIFF $count=2 $X=3.935
+ $Y=2.425 $X2=4.06 $Y2=3.59
r164 3 56 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=3.935
+ $Y=2.425 $X2=4.06 $Y2=2.57
r165 2 67 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1 $X=5.48
+ $Y=0.665 $X2=5.62 $Y2=1.49
r166 2 64 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.48
+ $Y=0.665 $X2=5.62 $Y2=0.81
r167 1 53 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1
+ $X=3.935 $Y=0.665 $X2=4.06 $Y2=1.49
r168 1 50 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1
+ $X=3.935 $Y=0.665 $X2=4.06 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_840_107# 1 2 3 4 15 19
+ 21 25 29 31 34 35 36 39 41 42 44 49 54 57 61 62 65 69 73 76 77 81
r157 78 80 22.525 $w=2.18e-07 $l=4.3e-07 $layer=LI1_cond $X=7.97 $Y=5.865
+ $X2=8.4 $Y2=5.865
r158 76 77 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.87
+ $Y=5.07 $X2=7.87 $Y2=5.07
r159 71 73 20.1678 $w=2.18e-07 $l=3.85e-07 $layer=LI1_cond $X=12.665 $Y=5.975
+ $X2=12.665 $Y2=6.36
r160 70 81 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=10.87 $Y=5.865
+ $X2=10.76 $Y2=5.865
r161 69 71 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=12.555 $Y=5.865
+ $X2=12.665 $Y2=5.975
r162 69 70 88.2667 $w=2.18e-07 $l=1.685e-06 $layer=LI1_cond $X=12.555 $Y=5.865
+ $X2=10.87 $Y2=5.865
r163 65 67 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=10.76 $Y=6.36
+ $X2=10.76 $Y2=7.04
r164 63 81 1.34256 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=10.76 $Y=5.975
+ $X2=10.76 $Y2=5.865
r165 63 65 20.1678 $w=2.18e-07 $l=3.85e-07 $layer=LI1_cond $X=10.76 $Y=5.975
+ $X2=10.76 $Y2=6.36
r166 62 80 5.76222 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=8.51 $Y=5.865
+ $X2=8.4 $Y2=5.865
r167 61 81 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=10.65 $Y=5.865
+ $X2=10.76 $Y2=5.865
r168 61 62 112.101 $w=2.18e-07 $l=2.14e-06 $layer=LI1_cond $X=10.65 $Y=5.865
+ $X2=8.51 $Y2=5.865
r169 57 59 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=8.4 $Y=6.36 $X2=8.4
+ $Y2=7.04
r170 55 80 0.716491 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=8.4 $Y=5.975
+ $X2=8.4 $Y2=5.865
r171 55 57 20.1678 $w=2.18e-07 $l=3.85e-07 $layer=LI1_cond $X=8.4 $Y=5.975
+ $X2=8.4 $Y2=6.36
r172 54 78 0.716491 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=7.97 $Y=5.755
+ $X2=7.97 $Y2=5.865
r173 53 76 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=7.97 $Y=5.235
+ $X2=7.97 $Y2=5.07
r174 53 54 27.2396 $w=2.18e-07 $l=5.2e-07 $layer=LI1_cond $X=7.97 $Y=5.235
+ $X2=7.97 $Y2=5.755
r175 49 52 53.4314 $w=2.18e-07 $l=1.02e-06 $layer=LI1_cond $X=7.97 $Y=3 $X2=7.97
+ $Y2=4.02
r176 47 76 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=7.97 $Y=4.905
+ $X2=7.97 $Y2=5.07
r177 47 52 46.3596 $w=2.18e-07 $l=8.85e-07 $layer=LI1_cond $X=7.97 $Y=4.905
+ $X2=7.97 $Y2=4.02
r178 43 77 143.386 $w=3.3e-07 $l=8.2e-07 $layer=POLY_cond $X=7.05 $Y=5.07
+ $X2=7.87 $Y2=5.07
r179 43 44 28.4028 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=7.05 $Y=5.07
+ $X2=6.8 $Y2=5.07
r180 37 44 0.400124 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.8 $Y=4.905
+ $X2=6.8 $Y2=5.07
r181 37 39 139.108 $w=5e-07 $l=1.3e-06 $layer=POLY_cond $X=6.8 $Y=4.905 $X2=6.8
+ $Y2=3.605
r182 35 44 28.4028 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=6.55 $Y=5.07
+ $X2=6.8 $Y2=5.07
r183 35 36 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=6.55 $Y=5.07
+ $X2=6.115 $Y2=5.07
r184 34 36 29.0934 $w=3.3e-07 $l=2.09105e-07 $layer=POLY_cond $X=6.015 $Y=4.905
+ $X2=6.115 $Y2=5.07
r185 33 34 926.758 $w=2e-07 $l=2.795e-06 $layer=POLY_cond $X=6.015 $Y=2.11
+ $X2=6.015 $Y2=4.905
r186 32 42 60.25 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=5.48 $Y=2.01 $X2=5.23
+ $Y2=2.01
r187 31 33 26.9307 $w=2e-07 $l=1.41421e-07 $layer=POLY_cond $X=5.915 $Y=2.01
+ $X2=6.015 $Y2=2.11
r188 31 32 144.236 $w=2e-07 $l=4.35e-07 $layer=POLY_cond $X=5.915 $Y=2.01
+ $X2=5.48 $Y2=2.01
r189 27 42 9.64 $w=5e-07 $l=1e-07 $layer=POLY_cond $X=5.23 $Y=2.11 $X2=5.23
+ $Y2=2.01
r190 27 29 113.961 $w=5e-07 $l=1.065e-06 $layer=POLY_cond $X=5.23 $Y=2.11
+ $X2=5.23 $Y2=3.175
r191 23 42 9.64 $w=5e-07 $l=1e-07 $layer=POLY_cond $X=5.23 $Y=1.91 $X2=5.23
+ $Y2=2.01
r192 23 25 79.7194 $w=5e-07 $l=7.45e-07 $layer=POLY_cond $X=5.23 $Y=1.91
+ $X2=5.23 $Y2=1.165
r193 22 41 18.8672 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=4.7 $Y=2.01 $X2=4.45
+ $Y2=2.01
r194 21 42 60.25 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=4.98 $Y=2.01 $X2=5.23
+ $Y2=2.01
r195 21 22 92.8416 $w=2e-07 $l=2.8e-07 $layer=POLY_cond $X=4.98 $Y=2.01 $X2=4.7
+ $Y2=2.01
r196 17 41 9.03033 $w=5e-07 $l=1e-07 $layer=POLY_cond $X=4.45 $Y=2.11 $X2=4.45
+ $Y2=2.01
r197 17 19 113.961 $w=5e-07 $l=1.065e-06 $layer=POLY_cond $X=4.45 $Y=2.11
+ $X2=4.45 $Y2=3.175
r198 13 41 9.03033 $w=5e-07 $l=1e-07 $layer=POLY_cond $X=4.45 $Y=1.91 $X2=4.45
+ $Y2=2.01
r199 13 15 79.7194 $w=5e-07 $l=7.45e-07 $layer=POLY_cond $X=4.45 $Y=1.91
+ $X2=4.45 $Y2=1.165
r200 4 52 300 $w=1.7e-07 $l=1.23301e-06 $layer=licon1_PDIFF $count=2 $X=7.83
+ $Y=2.855 $X2=7.97 $Y2=4.02
r201 4 49 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.83
+ $Y=2.855 $X2=7.97 $Y2=3
r202 3 73 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=12.54
+ $Y=6.215 $X2=12.665 $Y2=6.36
r203 2 67 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1
+ $X=10.62 $Y=6.215 $X2=10.76 $Y2=7.04
r204 2 65 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1
+ $X=10.62 $Y=6.215 $X2=10.76 $Y2=6.36
r205 1 59 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1 $X=8.26
+ $Y=6.215 $X2=8.4 $Y2=7.04
r206 1 57 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.26
+ $Y=6.215 $X2=8.4 $Y2=6.36
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_362_1243# 1 2 3 4 15 17
+ 20 22 23 26 30 34 41 44 46 49 51
r92 50 51 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=6.04 $Y=5.865
+ $X2=6.41 $Y2=5.865
r93 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.83
+ $Y=2.35 $X2=6.83 $Y2=2.35
r94 44 46 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.52 $Y=2.35 $X2=6.83
+ $Y2=2.35
r95 41 43 53.4314 $w=2.18e-07 $l=1.02e-06 $layer=LI1_cond $X=6.41 $Y=3 $X2=6.41
+ $Y2=4.02
r96 39 51 0.716491 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=6.41 $Y=5.755
+ $X2=6.41 $Y2=5.865
r97 39 43 90.8858 $w=2.18e-07 $l=1.735e-06 $layer=LI1_cond $X=6.41 $Y=5.755
+ $X2=6.41 $Y2=4.02
r98 38 44 7.17723 $w=3.3e-07 $l=2.13014e-07 $layer=LI1_cond $X=6.41 $Y=2.515
+ $X2=6.52 $Y2=2.35
r99 38 41 25.4061 $w=2.18e-07 $l=4.85e-07 $layer=LI1_cond $X=6.41 $Y=2.515
+ $X2=6.41 $Y2=3
r100 34 36 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=6.04 $Y=6.36
+ $X2=6.04 $Y2=7.04
r101 32 50 0.716491 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=6.04 $Y=5.975
+ $X2=6.04 $Y2=5.865
r102 32 34 20.1678 $w=2.18e-07 $l=3.85e-07 $layer=LI1_cond $X=6.04 $Y=5.975
+ $X2=6.04 $Y2=6.36
r103 31 49 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=3.79 $Y=5.865
+ $X2=3.68 $Y2=5.865
r104 30 50 5.76222 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=5.93 $Y=5.865
+ $X2=6.04 $Y2=5.865
r105 30 31 112.101 $w=2.18e-07 $l=2.14e-06 $layer=LI1_cond $X=5.93 $Y=5.865
+ $X2=3.79 $Y2=5.865
r106 26 28 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=3.68 $Y=6.36
+ $X2=3.68 $Y2=7.04
r107 24 49 1.34256 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=3.68 $Y=5.975
+ $X2=3.68 $Y2=5.865
r108 24 26 20.1678 $w=2.18e-07 $l=3.85e-07 $layer=LI1_cond $X=3.68 $Y=5.975
+ $X2=3.68 $Y2=6.36
r109 22 49 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=3.57 $Y=5.865
+ $X2=3.68 $Y2=5.865
r110 22 23 79.0995 $w=2.18e-07 $l=1.51e-06 $layer=LI1_cond $X=3.57 $Y=5.865
+ $X2=2.06 $Y2=5.865
r111 18 23 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=1.95 $Y=5.975
+ $X2=2.06 $Y2=5.865
r112 18 20 20.1678 $w=2.18e-07 $l=3.85e-07 $layer=LI1_cond $X=1.95 $Y=5.975
+ $X2=1.95 $Y2=6.36
r113 17 47 87.4306 $w=3.3e-07 $l=5e-07 $layer=POLY_cond $X=7.33 $Y=2.35 $X2=6.83
+ $Y2=2.35
r114 13 17 28.4267 $w=3.3e-07 $l=3.22102e-07 $layer=POLY_cond $X=7.58 $Y=2.515
+ $X2=7.33 $Y2=2.35
r115 13 15 116.636 $w=5e-07 $l=1.09e-06 $layer=POLY_cond $X=7.58 $Y=2.515
+ $X2=7.58 $Y2=3.605
r116 4 43 300 $w=1.7e-07 $l=1.22591e-06 $layer=licon1_PDIFF $count=2 $X=6.285
+ $Y=2.855 $X2=6.41 $Y2=4.02
r117 4 41 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=6.285
+ $Y=2.855 $X2=6.41 $Y2=3
r118 3 36 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1 $X=5.9
+ $Y=6.215 $X2=6.04 $Y2=7.04
r119 3 34 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.9
+ $Y=6.215 $X2=6.04 $Y2=6.36
r120 2 28 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1 $X=3.54
+ $Y=6.215 $X2=3.68 $Y2=7.04
r121 2 26 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.54
+ $Y=6.215 $X2=3.68 $Y2=6.36
r122 1 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.81
+ $Y=6.215 $X2=1.95 $Y2=6.36
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_2092_381# 1 2 9 11 12 15
+ 17 21 23 27 31 33 34 36 37 40 44 48 50
c96 40 0 1.29889e-19 $X=13.595 $Y=5.59
r97 46 50 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=13.995 $Y=5.755
+ $X2=13.995 $Y2=5.59
r98 46 48 31.6922 $w=2.18e-07 $l=6.05e-07 $layer=LI1_cond $X=13.995 $Y=5.755
+ $X2=13.995 $Y2=6.36
r99 42 50 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=13.995 $Y=5.425
+ $X2=13.995 $Y2=5.59
r100 42 44 52.1219 $w=2.18e-07 $l=9.95e-07 $layer=LI1_cond $X=13.995 $Y=5.425
+ $X2=13.995 $Y2=4.43
r101 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.595
+ $Y=5.59 $X2=13.595 $Y2=5.59
r102 37 50 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=13.885 $Y=5.59
+ $X2=13.995 $Y2=5.59
r103 37 39 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=13.885 $Y=5.59
+ $X2=13.595 $Y2=5.59
r104 35 40 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=13.305 $Y=5.59
+ $X2=13.595 $Y2=5.59
r105 35 36 19.9095 $w=3.3e-07 $l=5.81679e-07 $layer=POLY_cond $X=13.305 $Y=5.59
+ $X2=12.8 $Y2=5.425
r106 29 36 5.72191 $w=5e-07 $l=4.39375e-07 $layer=POLY_cond $X=13.055 $Y=5.755
+ $X2=12.8 $Y2=5.425
r107 29 31 71.6939 $w=5e-07 $l=6.7e-07 $layer=POLY_cond $X=13.055 $Y=5.755
+ $X2=13.055 $Y2=6.425
r108 25 36 5.72191 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=13.05 $Y=5.425
+ $X2=12.8 $Y2=5.425
r109 25 27 202.241 $w=5e-07 $l=1.89e-06 $layer=POLY_cond $X=13.05 $Y=5.425
+ $X2=13.05 $Y2=3.535
r110 24 34 37.8846 $w=2.2e-07 $l=2.5e-07 $layer=POLY_cond $X=12.52 $Y=5.535
+ $X2=12.27 $Y2=5.535
r111 23 36 19.9095 $w=2.2e-07 $l=1.1e-07 $layer=POLY_cond $X=12.8 $Y=5.535
+ $X2=12.8 $Y2=5.425
r112 23 24 81.6729 $w=2.2e-07 $l=2.8e-07 $layer=POLY_cond $X=12.8 $Y=5.535
+ $X2=12.52 $Y2=5.535
r113 19 34 5.40546 $w=5e-07 $l=1.1e-07 $layer=POLY_cond $X=12.27 $Y=5.425
+ $X2=12.27 $Y2=5.535
r114 19 21 202.241 $w=5e-07 $l=1.89e-06 $layer=POLY_cond $X=12.27 $Y=5.425
+ $X2=12.27 $Y2=3.535
r115 18 33 37.8846 $w=2.2e-07 $l=2.5e-07 $layer=POLY_cond $X=11.74 $Y=5.535
+ $X2=11.49 $Y2=5.535
r116 17 34 37.8846 $w=2.2e-07 $l=2.5e-07 $layer=POLY_cond $X=12.02 $Y=5.535
+ $X2=12.27 $Y2=5.535
r117 17 18 81.6729 $w=2.2e-07 $l=2.8e-07 $layer=POLY_cond $X=12.02 $Y=5.535
+ $X2=11.74 $Y2=5.535
r118 13 33 5.40546 $w=5e-07 $l=1.1e-07 $layer=POLY_cond $X=11.49 $Y=5.425
+ $X2=11.49 $Y2=5.535
r119 13 15 202.241 $w=5e-07 $l=1.89e-06 $layer=POLY_cond $X=11.49 $Y=5.425
+ $X2=11.49 $Y2=3.535
r120 11 33 37.8846 $w=2.2e-07 $l=2.5e-07 $layer=POLY_cond $X=11.24 $Y=5.535
+ $X2=11.49 $Y2=5.535
r121 11 12 81.6729 $w=2.2e-07 $l=2.8e-07 $layer=POLY_cond $X=11.24 $Y=5.535
+ $X2=10.96 $Y2=5.535
r122 7 12 32.6025 $w=2.2e-07 $l=3e-07 $layer=POLY_cond $X=10.71 $Y=5.425
+ $X2=10.96 $Y2=5.535
r123 7 9 202.241 $w=5e-07 $l=1.89e-06 $layer=POLY_cond $X=10.71 $Y=5.425
+ $X2=10.71 $Y2=3.535
r124 2 44 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=13.87
+ $Y=4.285 $X2=13.995 $Y2=4.43
r125 1 48 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=13.87
+ $Y=6.215 $X2=13.995 $Y2=6.36
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_1472_1171# 1 2 3 4 15 17
+ 18 21 24 25 26 27 31 33 37 39 40 44 45 47 48 49 51 55 57 59 63 67 69 71 74 77
+ 79 80
c156 33 0 1.1883e-19 $X=10.9 $Y=5.955
r157 73 74 38.5818 $w=2.28e-07 $l=7.7e-07 $layer=LI1_cond $X=19.825 $Y=1.565
+ $X2=19.825 $Y2=2.335
r158 72 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.495 $Y=2.42
+ $X2=19.33 $Y2=2.42
r159 71 74 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=19.71 $Y=2.42
+ $X2=19.825 $Y2=2.335
r160 71 72 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=19.71 $Y=2.42
+ $X2=19.495 $Y2=2.42
r161 70 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.44 $Y=1.48
+ $X2=19.355 $Y2=1.48
r162 69 73 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=19.71 $Y=1.48
+ $X2=19.825 $Y2=1.565
r163 69 70 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=19.71 $Y=1.48
+ $X2=19.44 $Y2=1.48
r164 65 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.355 $Y=1.395
+ $X2=19.355 $Y2=1.48
r165 65 67 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=19.355 $Y=1.395
+ $X2=19.355 $Y2=0.96
r166 61 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=19.33 $Y=2.505
+ $X2=19.33 $Y2=2.42
r167 61 63 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=19.33 $Y=2.505
+ $X2=19.33 $Y2=3.2
r168 60 76 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.595 $Y=2.42
+ $X2=18.43 $Y2=2.42
r169 59 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.165 $Y=2.42
+ $X2=19.33 $Y2=2.42
r170 59 60 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=19.165 $Y=2.42
+ $X2=18.595 $Y2=2.42
r171 58 77 6.31926 $w=1.95e-07 $l=1.36931e-07 $layer=LI1_cond $X=18.53 $Y=1.48
+ $X2=18.405 $Y2=1.455
r172 57 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.27 $Y=1.48
+ $X2=19.355 $Y2=1.48
r173 57 58 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=19.27 $Y=1.48
+ $X2=18.53 $Y2=1.48
r174 53 77 0.465126 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=18.405 $Y=1.345
+ $X2=18.405 $Y2=1.455
r175 53 55 17.7476 $w=2.48e-07 $l=3.85e-07 $layer=LI1_cond $X=18.405 $Y=1.345
+ $X2=18.405 $Y2=0.96
r176 49 76 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.43 $Y=2.505
+ $X2=18.43 $Y2=2.42
r177 49 51 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=18.43 $Y=2.505
+ $X2=18.43 $Y2=3.2
r178 47 77 6.31926 $w=1.95e-07 $l=1.25e-07 $layer=LI1_cond $X=18.28 $Y=1.455
+ $X2=18.405 $Y2=1.455
r179 47 48 208.749 $w=2.18e-07 $l=3.985e-06 $layer=LI1_cond $X=18.28 $Y=1.455
+ $X2=14.295 $Y2=1.455
r180 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.13
+ $Y=1.78 $X2=14.13 $Y2=1.78
r181 42 48 7.17723 $w=2.2e-07 $l=2.13014e-07 $layer=LI1_cond $X=14.13 $Y=1.565
+ $X2=14.295 $Y2=1.455
r182 42 44 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=14.13 $Y=1.565
+ $X2=14.13 $Y2=1.78
r183 41 45 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=14.13 $Y=1.535
+ $X2=14.13 $Y2=1.78
r184 35 37 37.7059 $w=9e-07 $l=6.6e-07 $layer=POLY_cond $X=11.35 $Y=6.055
+ $X2=11.35 $Y2=6.715
r185 34 40 56.5239 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=10.62 $Y=5.955
+ $X2=10.17 $Y2=5.955
r186 33 35 44.5077 $w=2e-07 $l=4.97494e-07 $layer=POLY_cond $X=10.9 $Y=5.955
+ $X2=11.35 $Y2=6.055
r187 33 34 92.8416 $w=2e-07 $l=2.8e-07 $layer=POLY_cond $X=10.9 $Y=5.955
+ $X2=10.62 $Y2=5.955
r188 29 40 12.0272 $w=9e-07 $l=1e-07 $layer=POLY_cond $X=10.17 $Y=6.055
+ $X2=10.17 $Y2=5.955
r189 29 31 37.7059 $w=9e-07 $l=6.6e-07 $layer=POLY_cond $X=10.17 $Y=6.055
+ $X2=10.17 $Y2=6.715
r190 28 39 25.8713 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=9.44 $Y=5.955
+ $X2=8.99 $Y2=5.955
r191 27 40 56.5239 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=9.72 $Y=5.955
+ $X2=10.17 $Y2=5.955
r192 27 28 92.8416 $w=2e-07 $l=2.8e-07 $layer=POLY_cond $X=9.72 $Y=5.955
+ $X2=9.44 $Y2=5.955
r193 25 41 29.0934 $w=2e-07 $l=2.09105e-07 $layer=POLY_cond $X=13.965 $Y=1.435
+ $X2=14.13 $Y2=1.535
r194 25 26 1657.89 $w=2e-07 $l=5e-06 $layer=POLY_cond $X=13.965 $Y=1.435
+ $X2=8.965 $Y2=1.435
r195 24 39 2.4532 $w=2e-07 $l=1.67705e-07 $layer=POLY_cond $X=8.865 $Y=5.855
+ $X2=8.99 $Y2=5.955
r196 23 26 26.9307 $w=2e-07 $l=1.41421e-07 $layer=POLY_cond $X=8.865 $Y=1.535
+ $X2=8.965 $Y2=1.435
r197 23 24 1432.41 $w=2e-07 $l=4.32e-06 $layer=POLY_cond $X=8.865 $Y=1.535
+ $X2=8.865 $Y2=5.855
r198 19 39 2.4532 $w=9e-07 $l=1e-07 $layer=POLY_cond $X=8.99 $Y=6.055 $X2=8.99
+ $Y2=5.955
r199 19 21 37.7059 $w=9e-07 $l=6.6e-07 $layer=POLY_cond $X=8.99 $Y=6.055
+ $X2=8.99 $Y2=6.715
r200 17 39 25.8713 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=8.54 $Y=5.955
+ $X2=8.99 $Y2=5.955
r201 17 18 92.8416 $w=2e-07 $l=2.8e-07 $layer=POLY_cond $X=8.54 $Y=5.955
+ $X2=8.26 $Y2=5.955
r202 13 18 44.5077 $w=2e-07 $l=4.97494e-07 $layer=POLY_cond $X=7.81 $Y=6.055
+ $X2=8.26 $Y2=5.955
r203 13 15 37.7059 $w=9e-07 $l=6.6e-07 $layer=POLY_cond $X=7.81 $Y=6.055
+ $X2=7.81 $Y2=6.715
r204 4 79 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=19.18
+ $Y=2.225 $X2=19.33 $Y2=2.5
r205 4 63 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=19.18
+ $Y=2.225 $X2=19.33 $Y2=3.2
r206 3 76 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=18.28
+ $Y=2.225 $X2=18.43 $Y2=2.5
r207 3 51 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=18.28
+ $Y=2.225 $X2=18.43 $Y2=3.2
r208 2 67 91 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=2 $X=19.215
+ $Y=0.755 $X2=19.355 $Y2=0.96
r209 1 55 91 $w=1.7e-07 $l=2.80936e-07 $layer=licon1_NDIFF $count=2 $X=18.265
+ $Y=0.755 $X2=18.445 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%SLEEP_B 3 7 10 11 14 15
c29 15 0 1.29889e-19 $X=14.82 $Y=5.71
r30 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.82
+ $Y=5.71 $X2=14.82 $Y2=5.71
r31 11 15 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=14.65 $Y=5.71
+ $X2=14.82 $Y2=5.71
r32 9 14 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=14.635 $Y=5.71
+ $X2=14.82 $Y2=5.71
r33 9 10 11.3528 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=14.635 $Y=5.71
+ $X2=14.385 $Y2=5.71
r34 5 10 14.2643 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.385 $Y=5.875
+ $X2=14.385 $Y2=5.71
r35 5 7 76.5092 $w=5e-07 $l=7.15e-07 $layer=POLY_cond $X=14.385 $Y=5.875
+ $X2=14.385 $Y2=6.59
r36 1 10 14.2643 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.385 $Y=5.545
+ $X2=14.385 $Y2=5.71
r37 1 3 94.7002 $w=5e-07 $l=8.85e-07 $layer=POLY_cond $X=14.385 $Y=5.545
+ $X2=14.385 $Y2=4.66
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_3617_1198# 1 2 9 11 13
+ 16 18 20 23 25 27 28 30 33 35 43 47 55 57 58 59 68
c116 23 0 7.81328e-20 $X=19.07 $Y=7.015
c117 9 0 7.81328e-20 $X=18.16 $Y=7.015
r118 68 69 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=19.525 $Y=6.197
+ $X2=19.54 $Y2=6.197
r119 65 66 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=19.07 $Y=6.197
+ $X2=19.075 $Y2=6.197
r120 64 65 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=18.625 $Y=6.197
+ $X2=19.07 $Y2=6.197
r121 63 64 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=18.59 $Y=6.197
+ $X2=18.625 $Y2=6.197
r122 60 61 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=18.16 $Y=6.197
+ $X2=18.175 $Y2=6.197
r123 55 59 6.00814 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=20.78 $Y=6.79
+ $X2=20.78 $Y2=6.625
r124 51 58 4.14384 $w=2.85e-07 $l=1.1e-07 $layer=LI1_cond $X=20.757 $Y=6.405
+ $X2=20.757 $Y2=6.295
r125 51 59 8.89605 $w=2.83e-07 $l=2.2e-07 $layer=LI1_cond $X=20.757 $Y=6.405
+ $X2=20.757 $Y2=6.625
r126 47 50 33.5624 $w=2.83e-07 $l=8.3e-07 $layer=LI1_cond $X=20.757 $Y=4.94
+ $X2=20.757 $Y2=5.77
r127 45 58 4.14384 $w=2.85e-07 $l=1.1e-07 $layer=LI1_cond $X=20.757 $Y=6.185
+ $X2=20.757 $Y2=6.295
r128 45 50 16.7812 $w=2.83e-07 $l=4.15e-07 $layer=LI1_cond $X=20.757 $Y=6.185
+ $X2=20.757 $Y2=5.77
r129 43 58 2.28927 $w=2.2e-07 $l=1.42e-07 $layer=LI1_cond $X=20.615 $Y=6.295
+ $X2=20.757 $Y2=6.295
r130 43 57 35.359 $w=2.18e-07 $l=6.75e-07 $layer=LI1_cond $X=20.615 $Y=6.295
+ $X2=19.94 $Y2=6.295
r131 42 68 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=19.45 $Y=6.197
+ $X2=19.525 $Y2=6.197
r132 42 66 48.8514 $w=3.7e-07 $l=3.75e-07 $layer=POLY_cond $X=19.45 $Y=6.197
+ $X2=19.075 $Y2=6.197
r133 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=19.45
+ $Y=6.24 $X2=19.45 $Y2=6.24
r134 38 63 20.8432 $w=3.7e-07 $l=1.6e-07 $layer=POLY_cond $X=18.43 $Y=6.197
+ $X2=18.59 $Y2=6.197
r135 38 61 33.2189 $w=3.7e-07 $l=2.55e-07 $layer=POLY_cond $X=18.43 $Y=6.197
+ $X2=18.175 $Y2=6.197
r136 37 41 27.337 $w=4.28e-07 $l=1.02e-06 $layer=LI1_cond $X=18.43 $Y=6.19
+ $X2=19.45 $Y2=6.19
r137 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=18.43
+ $Y=6.24 $X2=18.43 $Y2=6.24
r138 35 57 8.50315 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=19.725 $Y=6.19
+ $X2=19.94 $Y2=6.19
r139 35 41 7.37028 $w=4.28e-07 $l=2.75e-07 $layer=LI1_cond $X=19.725 $Y=6.19
+ $X2=19.45 $Y2=6.19
r140 31 69 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=19.54 $Y=6.405
+ $X2=19.54 $Y2=6.197
r141 31 33 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=19.54 $Y=6.405
+ $X2=19.54 $Y2=7.015
r142 28 68 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=19.525 $Y=5.99
+ $X2=19.525 $Y2=6.197
r143 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=19.525 $Y=5.99
+ $X2=19.525 $Y2=5.355
r144 25 66 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=19.075 $Y=5.99
+ $X2=19.075 $Y2=6.197
r145 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=19.075 $Y=5.99
+ $X2=19.075 $Y2=5.355
r146 21 65 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=19.07 $Y=6.405
+ $X2=19.07 $Y2=6.197
r147 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=19.07 $Y=6.405
+ $X2=19.07 $Y2=7.015
r148 18 64 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=18.625 $Y=5.99
+ $X2=18.625 $Y2=6.197
r149 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=18.625 $Y=5.99
+ $X2=18.625 $Y2=5.355
r150 14 63 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=18.59 $Y=6.405
+ $X2=18.59 $Y2=6.197
r151 14 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=18.59 $Y=6.405
+ $X2=18.59 $Y2=7.015
r152 11 61 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=18.175 $Y=5.99
+ $X2=18.175 $Y2=6.197
r153 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=18.175 $Y=5.99
+ $X2=18.175 $Y2=5.355
r154 7 60 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=18.16 $Y=6.405
+ $X2=18.16 $Y2=6.197
r155 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=18.16 $Y=6.405
+ $X2=18.16 $Y2=7.015
r156 2 50 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=20.635
+ $Y=4.795 $X2=20.785 $Y2=5.77
r157 2 47 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=20.635
+ $Y=4.795 $X2=20.785 $Y2=4.94
r158 1 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=20.64
+ $Y=6.645 $X2=20.78 $Y2=6.79
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_528_1171# 1 2 3 4 15 17
+ 18 21 23 27 29 33 36 37 38 40 41 42 44 45 46 49 51 53 54 56 59 61 63 66 68 70
+ 73 75 76 77 79 80 85 88 89 91 92 94 95 98 102 104 106 108 110 114 116 118 119
+ 130
c255 94 0 7.44113e-20 $X=18.29 $Y=6.66
c256 73 0 7.81328e-20 $X=19.57 $Y=1.125
c257 59 0 7.81328e-20 $X=18.66 $Y=1.125
r258 130 131 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=19.555 $Y=1.942
+ $X2=19.57 $Y2=1.942
r259 127 128 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=19.105 $Y=1.942
+ $X2=19.14 $Y2=1.942
r260 126 127 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=18.66 $Y=1.942
+ $X2=19.105 $Y2=1.942
r261 125 126 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=18.655 $Y=1.942
+ $X2=18.66 $Y2=1.942
r262 122 123 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=18.19 $Y=1.942
+ $X2=18.205 $Y2=1.942
r263 112 114 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=19.325 $Y=6.745
+ $X2=19.325 $Y2=6.79
r264 108 121 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=19.3 $Y=5.635
+ $X2=19.3 $Y2=5.72
r265 108 110 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=19.3 $Y=5.635
+ $X2=19.3 $Y2=4.94
r266 107 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.565 $Y=5.72
+ $X2=18.4 $Y2=5.72
r267 106 121 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.135 $Y=5.72
+ $X2=19.3 $Y2=5.72
r268 106 107 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=19.135 $Y=5.72
+ $X2=18.565 $Y2=5.72
r269 105 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.46 $Y=6.66
+ $X2=18.375 $Y2=6.66
r270 104 112 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=19.2 $Y=6.66
+ $X2=19.325 $Y2=6.745
r271 104 105 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=19.2 $Y=6.66
+ $X2=18.46 $Y2=6.66
r272 100 119 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.375 $Y=6.745
+ $X2=18.375 $Y2=6.66
r273 100 102 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=18.375 $Y=6.745
+ $X2=18.375 $Y2=6.79
r274 96 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.4 $Y=5.635
+ $X2=18.4 $Y2=5.72
r275 96 98 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=18.4 $Y=5.635
+ $X2=18.4 $Y2=4.94
r276 94 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.29 $Y=6.66
+ $X2=18.375 $Y2=6.66
r277 94 95 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=18.29 $Y=6.66
+ $X2=18.02 $Y2=6.66
r278 93 116 5.91331 $w=1.95e-07 $l=1.26886e-07 $layer=LI1_cond $X=18.02 $Y=5.72
+ $X2=17.905 $Y2=5.745
r279 92 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.235 $Y=5.72
+ $X2=18.4 $Y2=5.72
r280 92 93 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=18.235 $Y=5.72
+ $X2=18.02 $Y2=5.72
r281 91 95 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=17.905 $Y=6.575
+ $X2=18.02 $Y2=6.66
r282 90 116 0.755422 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=17.905 $Y=5.855
+ $X2=17.905 $Y2=5.745
r283 90 91 36.0765 $w=2.28e-07 $l=7.2e-07 $layer=LI1_cond $X=17.905 $Y=5.855
+ $X2=17.905 $Y2=6.575
r284 88 116 5.91331 $w=1.95e-07 $l=1.15e-07 $layer=LI1_cond $X=17.79 $Y=5.745
+ $X2=17.905 $Y2=5.745
r285 88 89 21.4773 $w=2.18e-07 $l=4.1e-07 $layer=LI1_cond $X=17.79 $Y=5.745
+ $X2=17.38 $Y2=5.745
r286 86 130 33.2189 $w=3.7e-07 $l=2.55e-07 $layer=POLY_cond $X=19.3 $Y=1.942
+ $X2=19.555 $Y2=1.942
r287 86 128 20.8432 $w=3.7e-07 $l=1.6e-07 $layer=POLY_cond $X=19.3 $Y=1.942
+ $X2=19.14 $Y2=1.942
r288 85 86 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=19.3
+ $Y=1.9 $X2=19.3 $Y2=1.9
r289 83 125 48.8514 $w=3.7e-07 $l=3.75e-07 $layer=POLY_cond $X=18.28 $Y=1.942
+ $X2=18.655 $Y2=1.942
r290 83 123 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=18.28 $Y=1.942
+ $X2=18.205 $Y2=1.942
r291 82 85 27.337 $w=4.28e-07 $l=1.02e-06 $layer=LI1_cond $X=18.28 $Y=1.95
+ $X2=19.3 $Y2=1.95
r292 82 83 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=18.28
+ $Y=1.9 $X2=18.28 $Y2=1.9
r293 80 82 24.1209 $w=4.28e-07 $l=9e-07 $layer=LI1_cond $X=17.38 $Y=1.95
+ $X2=18.28 $Y2=1.95
r294 79 89 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=17.27 $Y=5.635
+ $X2=17.38 $Y2=5.745
r295 78 80 7.78542 $w=4.3e-07 $l=2.64339e-07 $layer=LI1_cond $X=17.27 $Y=2.165
+ $X2=17.38 $Y2=1.95
r296 78 79 181.772 $w=2.18e-07 $l=3.47e-06 $layer=LI1_cond $X=17.27 $Y=2.165
+ $X2=17.27 $Y2=5.635
r297 71 131 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=19.57 $Y=1.735
+ $X2=19.57 $Y2=1.942
r298 71 73 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=19.57 $Y=1.735
+ $X2=19.57 $Y2=1.125
r299 68 130 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=19.555 $Y=2.15
+ $X2=19.555 $Y2=1.942
r300 68 70 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=19.555 $Y=2.15
+ $X2=19.555 $Y2=2.785
r301 64 128 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=19.14 $Y=1.735
+ $X2=19.14 $Y2=1.942
r302 64 66 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=19.14 $Y=1.735
+ $X2=19.14 $Y2=1.125
r303 61 127 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=19.105 $Y=2.15
+ $X2=19.105 $Y2=1.942
r304 61 63 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=19.105 $Y=2.15
+ $X2=19.105 $Y2=2.785
r305 57 126 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=18.66 $Y=1.735
+ $X2=18.66 $Y2=1.942
r306 57 59 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=18.66 $Y=1.735
+ $X2=18.66 $Y2=1.125
r307 54 125 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=18.655 $Y=2.15
+ $X2=18.655 $Y2=1.942
r308 54 56 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=18.655 $Y=2.15
+ $X2=18.655 $Y2=2.785
r309 51 123 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=18.205 $Y=2.15
+ $X2=18.205 $Y2=1.942
r310 51 53 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=18.205 $Y=2.15
+ $X2=18.205 $Y2=2.785
r311 47 122 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=18.19 $Y=1.735
+ $X2=18.19 $Y2=1.942
r312 47 49 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=18.19 $Y=1.735
+ $X2=18.19 $Y2=1.125
r313 45 122 10.4461 $w=3.7e-07 $l=9.3675e-08 $layer=POLY_cond $X=18.115 $Y=1.9
+ $X2=18.19 $Y2=1.942
r314 45 46 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=18.115 $Y=1.9
+ $X2=17.665 $Y2=1.9
r315 44 46 29.0934 $w=3.3e-07 $l=2.09105e-07 $layer=POLY_cond $X=17.565 $Y=1.735
+ $X2=17.665 $Y2=1.9
r316 43 44 202.262 $w=2e-07 $l=6.1e-07 $layer=POLY_cond $X=17.565 $Y=1.125
+ $X2=17.565 $Y2=1.735
r317 41 43 26.9361 $w=2.05e-07 $l=1.44599e-07 $layer=POLY_cond $X=17.465
+ $Y=1.022 $X2=17.565 $Y2=1.125
r318 41 42 2911.41 $w=2.05e-07 $l=9e-06 $layer=POLY_cond $X=17.465 $Y=1.022
+ $X2=8.465 $Y2=1.022
r319 39 42 26.9361 $w=2.05e-07 $l=1.44599e-07 $layer=POLY_cond $X=8.365 $Y=1.125
+ $X2=8.465 $Y2=1.022
r320 39 40 1432.41 $w=2e-07 $l=4.32e-06 $layer=POLY_cond $X=8.365 $Y=1.125
+ $X2=8.365 $Y2=5.445
r321 37 40 26.9307 $w=2e-07 $l=1.41421e-07 $layer=POLY_cond $X=8.265 $Y=5.545
+ $X2=8.365 $Y2=5.445
r322 37 38 392.919 $w=2e-07 $l=1.185e-06 $layer=POLY_cond $X=8.265 $Y=5.545
+ $X2=7.08 $Y2=5.545
r323 36 77 8.2592 $w=5.5e-07 $l=3.96863e-07 $layer=POLY_cond $X=6.98 $Y=5.855
+ $X2=6.63 $Y2=5.955
r324 35 38 26.9307 $w=2e-07 $l=1.41421e-07 $layer=POLY_cond $X=6.98 $Y=5.645
+ $X2=7.08 $Y2=5.545
r325 35 36 69.6312 $w=2e-07 $l=2.1e-07 $layer=POLY_cond $X=6.98 $Y=5.645
+ $X2=6.98 $Y2=5.855
r326 31 77 8.2592 $w=5.5e-07 $l=1e-07 $layer=POLY_cond $X=6.63 $Y=6.055 $X2=6.63
+ $Y2=5.955
r327 31 33 37.7059 $w=9e-07 $l=6.6e-07 $layer=POLY_cond $X=6.63 $Y=6.055
+ $X2=6.63 $Y2=6.715
r328 30 76 56.5239 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=5.9 $Y=5.955 $X2=5.45
+ $Y2=5.955
r329 29 77 20.3121 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=6.18 $Y=5.955
+ $X2=6.63 $Y2=5.955
r330 29 30 92.8416 $w=2e-07 $l=2.8e-07 $layer=POLY_cond $X=6.18 $Y=5.955 $X2=5.9
+ $Y2=5.955
r331 25 76 12.0272 $w=9e-07 $l=1e-07 $layer=POLY_cond $X=5.45 $Y=6.055 $X2=5.45
+ $Y2=5.955
r332 25 27 37.7059 $w=9e-07 $l=6.6e-07 $layer=POLY_cond $X=5.45 $Y=6.055
+ $X2=5.45 $Y2=6.715
r333 24 75 56.5239 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=4.72 $Y=5.955
+ $X2=4.27 $Y2=5.955
r334 23 76 56.5239 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=5 $Y=5.955 $X2=5.45
+ $Y2=5.955
r335 23 24 92.8416 $w=2e-07 $l=2.8e-07 $layer=POLY_cond $X=5 $Y=5.955 $X2=4.72
+ $Y2=5.955
r336 19 75 12.0272 $w=9e-07 $l=1e-07 $layer=POLY_cond $X=4.27 $Y=6.055 $X2=4.27
+ $Y2=5.955
r337 19 21 37.7059 $w=9e-07 $l=6.6e-07 $layer=POLY_cond $X=4.27 $Y=6.055
+ $X2=4.27 $Y2=6.715
r338 17 75 56.5239 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=3.82 $Y=5.955
+ $X2=4.27 $Y2=5.955
r339 17 18 92.8416 $w=2e-07 $l=2.8e-07 $layer=POLY_cond $X=3.82 $Y=5.955
+ $X2=3.54 $Y2=5.955
r340 13 18 44.5077 $w=2e-07 $l=4.97494e-07 $layer=POLY_cond $X=3.09 $Y=6.055
+ $X2=3.54 $Y2=5.955
r341 13 15 37.7059 $w=9e-07 $l=6.6e-07 $layer=POLY_cond $X=3.09 $Y=6.055
+ $X2=3.09 $Y2=6.715
r342 4 121 400 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=19.15
+ $Y=4.795 $X2=19.3 $Y2=5.64
r343 4 110 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=19.15
+ $Y=4.795 $X2=19.3 $Y2=4.94
r344 3 118 400 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=18.25
+ $Y=4.795 $X2=18.4 $Y2=5.64
r345 3 98 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=18.25
+ $Y=4.795 $X2=18.4 $Y2=4.94
r346 2 114 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=19.145
+ $Y=6.645 $X2=19.285 $Y2=6.79
r347 1 102 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=18.235
+ $Y=6.645 $X2=18.375 $Y2=6.79
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A 1 2 3 5 8 10 12 14 16 18
+ 19 20
r53 23 25 11.0663 $w=3.92e-07 $l=9e-08 $layer=POLY_cond $X=21.16 $Y=6.29
+ $X2=21.16 $Y2=6.38
r54 20 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=21.235
+ $Y=6.29 $X2=21.235 $Y2=6.29
r55 16 23 56.0318 $w=3.92e-07 $l=3.67423e-07 $layer=POLY_cond $X=21.01 $Y=5.99
+ $X2=21.16 $Y2=6.29
r56 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=21.01 $Y=5.99
+ $X2=21.01 $Y2=5.355
r57 12 25 28.3659 $w=3.92e-07 $l=1.98997e-07 $layer=POLY_cond $X=20.995 $Y=6.455
+ $X2=21.16 $Y2=6.38
r58 12 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=20.995 $Y=6.455
+ $X2=20.995 $Y2=7.015
r59 11 19 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=20.65 $Y=6.38
+ $X2=20.56 $Y2=6.38
r60 10 25 25.3688 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=20.92 $Y=6.38
+ $X2=21.16 $Y2=6.38
r61 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=20.92 $Y=6.38
+ $X2=20.65 $Y2=6.38
r62 6 19 18.8402 $w=1.65e-07 $l=7.74597e-08 $layer=POLY_cond $X=20.565 $Y=6.455
+ $X2=20.56 $Y2=6.38
r63 6 8 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=20.565 $Y=6.455
+ $X2=20.565 $Y2=7.015
r64 3 5 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=20.56 $Y=5.99
+ $X2=20.56 $Y2=5.355
r65 2 19 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=20.56 $Y=6.305
+ $X2=20.56 $Y2=6.38
r66 1 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=20.56 $Y=6.08 $X2=20.56
+ $Y2=5.99
r67 1 2 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=20.56 $Y=6.08
+ $X2=20.56 $Y2=6.305
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%X 1 2 3 4 15 19 23 29 33
+ 34
c61 33 0 1.1774e-19 $X=2.73 $Y=2.03
r62 40 42 124.673 $w=2.18e-07 $l=2.38e-06 $layer=LI1_cond $X=1.17 $Y=2.57
+ $X2=1.17 $Y2=4.95
r63 34 37 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=1.17 $Y=2.03 $X2=1.17
+ $Y2=2.14
r64 34 40 22.2631 $w=2.18e-07 $l=4.25e-07 $layer=LI1_cond $X=1.17 $Y=2.145
+ $X2=1.17 $Y2=2.57
r65 34 37 0.261919 $w=2.18e-07 $l=5e-09 $layer=LI1_cond $X=1.17 $Y=2.145
+ $X2=1.17 $Y2=2.14
r66 29 31 124.673 $w=2.18e-07 $l=2.38e-06 $layer=LI1_cond $X=2.73 $Y=2.57
+ $X2=2.73 $Y2=4.95
r67 27 33 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=2.73 $Y=2.14 $X2=2.73
+ $Y2=2.03
r68 27 29 22.525 $w=2.18e-07 $l=4.3e-07 $layer=LI1_cond $X=2.73 $Y=2.14 $X2=2.73
+ $Y2=2.57
r69 23 26 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=2.73 $Y=0.81 $X2=2.73
+ $Y2=1.49
r70 21 33 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=2.73 $Y=1.92 $X2=2.73
+ $Y2=2.03
r71 21 26 22.525 $w=2.18e-07 $l=4.3e-07 $layer=LI1_cond $X=2.73 $Y=1.92 $X2=2.73
+ $Y2=1.49
r72 20 34 1.34256 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=1.28 $Y=2.03 $X2=1.17
+ $Y2=2.03
r73 19 33 1.34256 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=2.62 $Y=2.03 $X2=2.73
+ $Y2=2.03
r74 19 20 70.1943 $w=2.18e-07 $l=1.34e-06 $layer=LI1_cond $X=2.62 $Y=2.03
+ $X2=1.28 $Y2=2.03
r75 15 18 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=1.17 $Y=0.81 $X2=1.17
+ $Y2=1.49
r76 13 34 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=1.17 $Y=1.92 $X2=1.17
+ $Y2=2.03
r77 13 18 22.525 $w=2.18e-07 $l=4.3e-07 $layer=LI1_cond $X=1.17 $Y=1.92 $X2=1.17
+ $Y2=1.49
r78 4 31 150 $w=1.7e-07 $l=2.59406e-06 $layer=licon1_PDIFF $count=4 $X=2.59
+ $Y=2.425 $X2=2.73 $Y2=4.95
r79 4 29 150 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=4 $X=2.59
+ $Y=2.425 $X2=2.73 $Y2=2.57
r80 3 42 150 $w=1.7e-07 $l=2.58675e-06 $layer=licon1_PDIFF $count=4 $X=1.045
+ $Y=2.425 $X2=1.17 $Y2=4.95
r81 3 40 150 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=4 $X=1.045
+ $Y=2.425 $X2=1.17 $Y2=2.57
r82 2 26 121.333 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_NDIFF $count=1 $X=2.59
+ $Y=0.665 $X2=2.73 $Y2=1.49
r83 2 23 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.59
+ $Y=0.665 $X2=2.73 $Y2=0.81
r84 1 18 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.665 $X2=1.17 $Y2=1.49
r85 1 15 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.665 $X2=1.17 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%VPWR 1 2 3 4 5 6 7 24 32
+ 38 40 44 49 52 53 56 61 64 68 73 76 78 80 81 82 87 90 97 99 104 106 117 124
+ 131 132 136 142 152
c264 80 0 1.1883e-19 $X=11.88 $Y=5.145
r265 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.77 $Y=4.51
+ $X2=14.77 $Y2=4.51
r266 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.62 $Y=3.63
+ $X2=13.62 $Y2=3.63
r267 129 131 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=13.44 $Y=3.63
+ $X2=13.62 $Y2=3.63
r268 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.06 $Y=3.63
+ $X2=12.06 $Y2=3.63
r269 122 124 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=11.88 $Y=3.63
+ $X2=12.06 $Y2=3.63
r270 118 125 0.598892 $w=3.7e-07 $l=1.56e-06 $layer=MET1_cond $X=10.5 $Y=3.63
+ $X2=12.06 $Y2=3.63
r271 118 142 0.0422296 $w=3.7e-07 $l=1.1e-07 $layer=MET1_cond $X=10.5 $Y=3.63
+ $X2=10.39 $Y2=3.63
r272 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.5 $Y=3.63
+ $X2=10.5 $Y2=3.63
r273 115 117 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=10.32 $Y=3.63
+ $X2=10.5 $Y2=3.63
r274 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.835 $Y=3.63
+ $X2=4.835 $Y2=3.63
r275 107 152 2.50498 $w=3.7e-07 $l=6.525e-06 $layer=MET1_cond $X=3.69 $Y=4.51
+ $X2=10.215 $Y2=4.51
r276 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.69 $Y=4.51
+ $X2=3.69 $Y2=4.51
r277 104 106 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.51 $Y=4.51
+ $X2=3.69 $Y2=4.51
r278 100 107 0.598892 $w=3.7e-07 $l=1.56e-06 $layer=MET1_cond $X=2.13 $Y=4.51
+ $X2=3.69 $Y2=4.51
r279 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.13 $Y=4.51
+ $X2=2.13 $Y2=4.51
r280 97 99 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.95 $Y=4.51
+ $X2=2.13 $Y2=4.51
r281 93 136 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=14.41 $Y=4.51
+ $X2=14.77 $Y2=4.51
r282 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.41 $Y=4.51
+ $X2=14.41 $Y2=4.51
r283 90 135 3.40825 $w=2.3e-07 $l=1.43875e-07 $layer=LI1_cond $X=14.655 $Y=4.51
+ $X2=14.77 $Y2=4.445
r284 90 92 12.276 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=14.655 $Y=4.51
+ $X2=14.41 $Y2=4.51
r285 88 142 1.99439 $w=3.7e-07 $l=5.195e-06 $layer=MET1_cond $X=5.195 $Y=3.63
+ $X2=10.39 $Y2=3.63
r286 88 111 0.138206 $w=3.7e-07 $l=3.6e-07 $layer=MET1_cond $X=5.195 $Y=3.63
+ $X2=4.835 $Y2=3.63
r287 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.195 $Y=3.63
+ $X2=5.195 $Y2=3.63
r288 85 110 3.33769 $w=2.4e-07 $l=1.15e-07 $layer=LI1_cond $X=4.955 $Y=3.635
+ $X2=4.84 $Y2=3.635
r289 85 87 11.5244 $w=2.38e-07 $l=2.4e-07 $layer=LI1_cond $X=4.955 $Y=3.635
+ $X2=5.195 $Y2=3.635
r290 82 93 0.740937 $w=3.7e-07 $l=1.93e-06 $layer=MET1_cond $X=12.48 $Y=4.51
+ $X2=14.41 $Y2=4.51
r291 82 152 0.869546 $w=3.7e-07 $l=2.265e-06 $layer=MET1_cond $X=12.48 $Y=4.51
+ $X2=10.215 $Y2=4.51
r292 81 132 0.437652 $w=3.7e-07 $l=1.14e-06 $layer=MET1_cond $X=12.48 $Y=3.63
+ $X2=13.62 $Y2=3.63
r293 81 125 0.16124 $w=3.7e-07 $l=4.2e-07 $layer=MET1_cond $X=12.48 $Y=3.63
+ $X2=12.06 $Y2=3.63
r294 76 135 3.40825 $w=2.3e-07 $l=1.8e-07 $layer=LI1_cond $X=14.77 $Y=4.625
+ $X2=14.77 $Y2=4.445
r295 76 78 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=14.77 $Y=4.625
+ $X2=14.77 $Y2=4.77
r296 73 75 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=13.44 $Y=3.88
+ $X2=13.44 $Y2=4.56
r297 71 75 24.8823 $w=2.18e-07 $l=4.75e-07 $layer=LI1_cond $X=13.44 $Y=5.035
+ $X2=13.44 $Y2=4.56
r298 70 129 0.986088 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=13.44 $Y=3.745
+ $X2=13.44 $Y2=3.63
r299 70 73 7.07181 $w=2.18e-07 $l=1.35e-07 $layer=LI1_cond $X=13.44 $Y=3.745
+ $X2=13.44 $Y2=3.88
r300 66 129 0.986088 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=13.44 $Y=3.515
+ $X2=13.44 $Y2=3.63
r301 66 68 69.9323 $w=2.18e-07 $l=1.335e-06 $layer=LI1_cond $X=13.44 $Y=3.515
+ $X2=13.44 $Y2=2.18
r302 65 80 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=11.99 $Y=5.145
+ $X2=11.88 $Y2=5.145
r303 64 71 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=13.33 $Y=5.145
+ $X2=13.44 $Y2=5.035
r304 64 65 70.1943 $w=2.18e-07 $l=1.34e-06 $layer=LI1_cond $X=13.33 $Y=5.145
+ $X2=11.99 $Y2=5.145
r305 61 63 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=11.88 $Y=3.88
+ $X2=11.88 $Y2=4.56
r306 59 80 1.34256 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=11.88 $Y=5.035
+ $X2=11.88 $Y2=5.145
r307 59 63 24.8823 $w=2.18e-07 $l=4.75e-07 $layer=LI1_cond $X=11.88 $Y=5.035
+ $X2=11.88 $Y2=4.56
r308 58 122 0.986088 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=11.88 $Y=3.745
+ $X2=11.88 $Y2=3.63
r309 58 61 7.07181 $w=2.18e-07 $l=1.35e-07 $layer=LI1_cond $X=11.88 $Y=3.745
+ $X2=11.88 $Y2=3.88
r310 54 122 0.986088 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=11.88 $Y=3.515
+ $X2=11.88 $Y2=3.63
r311 54 56 69.9323 $w=2.18e-07 $l=1.335e-06 $layer=LI1_cond $X=11.88 $Y=3.515
+ $X2=11.88 $Y2=2.18
r312 52 80 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=11.77 $Y=5.145
+ $X2=11.88 $Y2=5.145
r313 52 53 70.1943 $w=2.18e-07 $l=1.34e-06 $layer=LI1_cond $X=11.77 $Y=5.145
+ $X2=10.43 $Y2=5.145
r314 49 51 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=10.32 $Y=3.88
+ $X2=10.32 $Y2=4.56
r315 47 53 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=10.32 $Y=5.035
+ $X2=10.43 $Y2=5.145
r316 47 51 24.8823 $w=2.18e-07 $l=4.75e-07 $layer=LI1_cond $X=10.32 $Y=5.035
+ $X2=10.32 $Y2=4.56
r317 46 115 0.986088 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=10.32 $Y=3.745
+ $X2=10.32 $Y2=3.63
r318 46 49 7.07181 $w=2.18e-07 $l=1.35e-07 $layer=LI1_cond $X=10.32 $Y=3.745
+ $X2=10.32 $Y2=3.88
r319 42 115 0.986088 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=10.32 $Y=3.515
+ $X2=10.32 $Y2=3.63
r320 42 44 69.9323 $w=2.18e-07 $l=1.335e-06 $layer=LI1_cond $X=10.32 $Y=3.515
+ $X2=10.32 $Y2=2.18
r321 38 110 3.48281 $w=2.3e-07 $l=1.2e-07 $layer=LI1_cond $X=4.84 $Y=3.515
+ $X2=4.84 $Y2=3.635
r322 38 40 47.3504 $w=2.28e-07 $l=9.45e-07 $layer=LI1_cond $X=4.84 $Y=3.515
+ $X2=4.84 $Y2=2.57
r323 32 35 85.1806 $w=2.28e-07 $l=1.7e-06 $layer=LI1_cond $X=3.51 $Y=2.57
+ $X2=3.51 $Y2=4.27
r324 30 104 0.716491 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=3.51 $Y=4.395
+ $X2=3.51 $Y2=4.51
r325 30 35 6.26328 $w=2.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.51 $Y=4.395
+ $X2=3.51 $Y2=4.27
r326 24 27 85.1806 $w=2.28e-07 $l=1.7e-06 $layer=LI1_cond $X=1.95 $Y=2.57
+ $X2=1.95 $Y2=4.27
r327 22 97 0.716491 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=1.95 $Y=4.395
+ $X2=1.95 $Y2=4.51
r328 22 27 6.26328 $w=2.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.95 $Y=4.395
+ $X2=1.95 $Y2=4.27
r329 7 135 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=14.635
+ $Y=4.285 $X2=14.775 $Y2=4.43
r330 7 78 600 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=1 $X=14.635
+ $Y=4.285 $X2=14.775 $Y2=4.77
r331 6 129 240 $w=1.7e-07 $l=1.57344e-06 $layer=licon1_PDIFF $count=2 $X=13.3
+ $Y=2.035 $X2=13.44 $Y2=3.54
r332 6 75 400 $w=1.7e-07 $l=2.59406e-06 $layer=licon1_PDIFF $count=1 $X=13.3
+ $Y=2.035 $X2=13.44 $Y2=4.56
r333 6 73 400 $w=1.7e-07 $l=1.91372e-06 $layer=licon1_PDIFF $count=1 $X=13.3
+ $Y=2.035 $X2=13.44 $Y2=3.88
r334 6 68 240 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=13.3
+ $Y=2.035 $X2=13.44 $Y2=2.18
r335 5 122 240 $w=1.7e-07 $l=1.57344e-06 $layer=licon1_PDIFF $count=2 $X=11.74
+ $Y=2.035 $X2=11.88 $Y2=3.54
r336 5 63 400 $w=1.7e-07 $l=2.59406e-06 $layer=licon1_PDIFF $count=1 $X=11.74
+ $Y=2.035 $X2=11.88 $Y2=4.56
r337 5 61 400 $w=1.7e-07 $l=1.91372e-06 $layer=licon1_PDIFF $count=1 $X=11.74
+ $Y=2.035 $X2=11.88 $Y2=3.88
r338 5 56 240 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=11.74
+ $Y=2.035 $X2=11.88 $Y2=2.18
r339 4 115 240 $w=1.7e-07 $l=1.56625e-06 $layer=licon1_PDIFF $count=2 $X=10.195
+ $Y=2.035 $X2=10.32 $Y2=3.54
r340 4 51 400 $w=1.7e-07 $l=2.58675e-06 $layer=licon1_PDIFF $count=1 $X=10.195
+ $Y=2.035 $X2=10.32 $Y2=4.56
r341 4 49 400 $w=1.7e-07 $l=1.90648e-06 $layer=licon1_PDIFF $count=1 $X=10.195
+ $Y=2.035 $X2=10.32 $Y2=3.88
r342 4 44 240 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=10.195
+ $Y=2.035 $X2=10.32 $Y2=2.18
r343 3 110 300 $w=1.7e-07 $l=1.23301e-06 $layer=licon1_PDIFF $count=2 $X=4.7
+ $Y=2.425 $X2=4.84 $Y2=3.59
r344 3 40 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.7
+ $Y=2.425 $X2=4.84 $Y2=2.57
r345 2 104 300 $w=1.7e-07 $l=2.25391e-06 $layer=licon1_PDIFF $count=2 $X=3.37
+ $Y=2.425 $X2=3.51 $Y2=4.61
r346 2 35 200 $w=1.7e-07 $l=1.91372e-06 $layer=licon1_PDIFF $count=3 $X=3.37
+ $Y=2.425 $X2=3.51 $Y2=4.27
r347 2 32 200 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=3 $X=3.37
+ $Y=2.425 $X2=3.51 $Y2=2.57
r348 1 97 300 $w=1.7e-07 $l=2.25391e-06 $layer=licon1_PDIFF $count=2 $X=1.81
+ $Y=2.425 $X2=1.95 $Y2=4.61
r349 1 27 200 $w=1.7e-07 $l=1.91372e-06 $layer=licon1_PDIFF $count=3 $X=1.81
+ $Y=2.425 $X2=1.95 $Y2=4.27
r350 1 24 200 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=3 $X=1.81
+ $Y=2.425 $X2=1.95 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_1410_571# 1 2 3 12 15 17
+ 18 19 22 26 30 37 41 43
r92 39 41 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.32 $Y=2.54
+ $X2=7.69 $Y2=2.54
r93 35 37 6.51381 $w=2.28e-07 $l=1.3e-07 $layer=LI1_cond $X=7.19 $Y=2.95
+ $X2=7.32 $Y2=2.95
r94 30 32 124.673 $w=2.18e-07 $l=2.38e-06 $layer=LI1_cond $X=12.66 $Y=2.18
+ $X2=12.66 $Y2=4.56
r95 28 30 19.6439 $w=2.18e-07 $l=3.75e-07 $layer=LI1_cond $X=12.66 $Y=1.805
+ $X2=12.66 $Y2=2.18
r96 27 43 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=11.21 $Y=1.695
+ $X2=11.1 $Y2=1.695
r97 26 28 6.81649 $w=2.2e-07 $l=1.55563e-07 $layer=LI1_cond $X=12.55 $Y=1.695
+ $X2=12.66 $Y2=1.805
r98 26 27 70.1943 $w=2.18e-07 $l=1.34e-06 $layer=LI1_cond $X=12.55 $Y=1.695
+ $X2=11.21 $Y2=1.695
r99 22 24 124.673 $w=2.18e-07 $l=2.38e-06 $layer=LI1_cond $X=11.1 $Y=2.18
+ $X2=11.1 $Y2=4.56
r100 20 43 1.34256 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=11.1 $Y=1.805
+ $X2=11.1 $Y2=1.695
r101 20 22 19.6439 $w=2.18e-07 $l=3.75e-07 $layer=LI1_cond $X=11.1 $Y=1.805
+ $X2=11.1 $Y2=2.18
r102 18 43 5.16603 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=10.99 $Y=1.695
+ $X2=11.1 $Y2=1.695
r103 18 19 166.842 $w=2.18e-07 $l=3.185e-06 $layer=LI1_cond $X=10.99 $Y=1.695
+ $X2=7.805 $Y2=1.695
r104 17 41 0.716491 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=7.69 $Y=2.425
+ $X2=7.69 $Y2=2.54
r105 16 19 6.82087 $w=2.2e-07 $l=1.60857e-07 $layer=LI1_cond $X=7.69 $Y=1.805
+ $X2=7.805 $Y2=1.695
r106 16 17 31.0659 $w=2.28e-07 $l=6.2e-07 $layer=LI1_cond $X=7.69 $Y=1.805
+ $X2=7.69 $Y2=2.425
r107 15 37 0.716491 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=7.32 $Y=2.835
+ $X2=7.32 $Y2=2.95
r108 14 39 0.716491 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=7.32 $Y=2.655
+ $X2=7.32 $Y2=2.54
r109 14 15 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=7.32 $Y=2.655
+ $X2=7.32 $Y2=2.835
r110 10 35 0.716491 $w=2.3e-07 $l=1.15e-07 $layer=LI1_cond $X=7.19 $Y=3.065
+ $X2=7.19 $Y2=2.95
r111 10 12 47.8514 $w=2.28e-07 $l=9.55e-07 $layer=LI1_cond $X=7.19 $Y=3.065
+ $X2=7.19 $Y2=4.02
r112 3 32 150 $w=1.7e-07 $l=2.59406e-06 $layer=licon1_PDIFF $count=4 $X=12.52
+ $Y=2.035 $X2=12.66 $Y2=4.56
r113 3 30 150 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=4 $X=12.52
+ $Y=2.035 $X2=12.66 $Y2=2.18
r114 2 24 150 $w=1.7e-07 $l=2.59406e-06 $layer=licon1_PDIFF $count=4 $X=10.96
+ $Y=2.035 $X2=11.1 $Y2=4.56
r115 2 22 150 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=4 $X=10.96
+ $Y=2.035 $X2=11.1 $Y2=2.18
r116 1 35 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.05
+ $Y=2.855 $X2=7.19 $Y2=3
r117 1 12 300 $w=1.7e-07 $l=1.23301e-06 $layer=licon1_PDIFF $count=2 $X=7.05
+ $Y=2.855 $X2=7.19 $Y2=4.02
.ends

