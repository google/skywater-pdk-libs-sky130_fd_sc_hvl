* File: sky130_fd_sc_hvl__and2_1.spice
* Created: Fri Aug 28 09:32:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__and2_1.pex.spice"
.subckt sky130_fd_sc_hvl__and2_1  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 A_183_107# N_A_M1005_g N_A_30_107#_M1005_s N_VNB_M1005_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=13.566 NRS=0 M=1 R=0.84 SA=250000
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g A_183_107# N_VNB_M1005_b NHV L=0.5 W=0.42
+ AD=0.157392 AS=0.0441 PD=1.12718 PS=0.63 NRD=86.7768 NRS=13.566 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1002 N_X_M1002_d N_A_30_107#_M1002_g N_VGND_M1004_d N_VNB_M1005_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.281058 PD=2.03 PS=2.01282 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1001 N_A_30_107#_M1001_d N_A_M1001_g N_VPWR_M1001_s N_VPB_M1001_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250002 A=0.21 P=1.84 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_A_30_107#_M1001_d N_VPB_M1001_b PHV L=0.5
+ W=0.42 AD=0.138075 AS=0.0588 PD=0.875 PS=0.7 NRD=52.2958 NRS=0 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1000 N_X_M1000_d N_A_30_107#_M1000_g N_VPWR_M1003_d N_VPB_M1001_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.493125 PD=3.57 PS=3.125 NRD=0 NRS=13.37 M=1 R=3 SA=250001
+ SB=250000 A=0.75 P=4 MULT=1
DX6_noxref N_VNB_M1005_b N_VPB_M1001_b NWDIODE A=10.452 P=13.24
*
.include "sky130_fd_sc_hvl__and2_1.pxi.spice"
*
.ends
*
*
