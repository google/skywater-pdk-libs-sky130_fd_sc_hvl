# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__dlrtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__dlrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.570000 1.930000 0.900000 2.600000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.735000 2.175000 9.475000 3.755000 ;
        RECT 9.140000 0.495000 9.475000 2.175000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.515000 0.810000 8.120000 1.780000 ;
        RECT 7.515000 1.780000 7.845000 1.855000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.175000 1.795000 1.400000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 9.600000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 9.600000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 9.600000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 9.600000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.985000 9.600000 4.155000 ;
      RECT 0.140000  0.495000 0.390000 1.580000 ;
      RECT 0.140000  1.580000 1.795000 1.675000 ;
      RECT 0.140000  1.675000 3.655000 1.750000 ;
      RECT 0.140000  1.750000 0.390000 3.610000 ;
      RECT 0.570000  0.365000 1.520000 0.995000 ;
      RECT 0.570000  2.780000 1.520000 3.705000 ;
      RECT 1.625000  1.750000 3.655000 1.845000 ;
      RECT 1.700000  0.495000 2.145000 0.995000 ;
      RECT 1.700000  2.025000 4.435000 2.195000 ;
      RECT 1.700000  2.195000 2.030000 3.610000 ;
      RECT 1.975000  0.995000 2.145000 1.325000 ;
      RECT 1.975000  1.325000 4.005000 1.495000 ;
      RECT 2.290000  2.375000 4.785000 2.545000 ;
      RECT 2.290000  2.545000 2.620000 3.245000 ;
      RECT 2.370000  0.495000 2.620000 0.975000 ;
      RECT 2.370000  0.975000 4.495000 1.145000 ;
      RECT 2.800000  0.365000 3.750000 0.795000 ;
      RECT 2.800000  2.725000 3.750000 3.705000 ;
      RECT 3.835000  1.495000 4.005000 1.605000 ;
      RECT 3.835000  1.605000 4.435000 2.025000 ;
      RECT 4.185000  1.145000 4.495000 1.225000 ;
      RECT 4.185000  1.225000 4.785000 1.395000 ;
      RECT 4.560000  2.725000 5.525000 2.895000 ;
      RECT 4.560000  2.895000 4.890000 3.245000 ;
      RECT 4.615000  1.395000 4.785000 1.965000 ;
      RECT 4.615000  1.965000 5.175000 2.295000 ;
      RECT 4.615000  2.295000 4.785000 2.375000 ;
      RECT 4.675000  0.495000 5.135000 0.995000 ;
      RECT 4.965000  0.995000 5.135000 1.175000 ;
      RECT 4.965000  1.175000 6.780000 1.345000 ;
      RECT 5.355000  1.345000 5.525000 2.725000 ;
      RECT 5.545000  0.365000 6.495000 0.995000 ;
      RECT 5.705000  2.255000 6.655000 3.705000 ;
      RECT 5.810000  1.525000 6.140000 1.905000 ;
      RECT 5.810000  1.905000 7.130000 2.035000 ;
      RECT 5.810000  2.035000 8.470000 2.075000 ;
      RECT 6.450000  1.345000 6.780000 1.725000 ;
      RECT 6.755000  0.495000 7.130000 0.995000 ;
      RECT 6.960000  0.995000 7.130000 1.905000 ;
      RECT 6.960000  2.075000 8.470000 2.205000 ;
      RECT 6.960000  2.205000 7.390000 3.005000 ;
      RECT 7.570000  2.385000 8.520000 3.755000 ;
      RECT 8.300000  0.365000 8.890000 1.325000 ;
      RECT 8.300000  1.665000 8.630000 1.995000 ;
      RECT 8.300000  1.995000 8.470000 2.035000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.600000  0.395000 0.770000 0.565000 ;
      RECT 0.600000  3.505000 0.770000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.960000  0.395000 1.130000 0.565000 ;
      RECT 0.960000  3.505000 1.130000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.320000  0.395000 1.490000 0.565000 ;
      RECT 1.320000  3.505000 1.490000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.830000  0.395000 3.000000 0.565000 ;
      RECT 2.830000  3.505000 3.000000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.190000  0.395000 3.360000 0.565000 ;
      RECT 3.190000  3.505000 3.360000 3.675000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.550000  0.395000 3.720000 0.565000 ;
      RECT 3.550000  3.505000 3.720000 3.675000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.985000 5.605000 4.155000 ;
      RECT 5.575000  0.395000 5.745000 0.565000 ;
      RECT 5.735000  3.505000 5.905000 3.675000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.985000 6.085000 4.155000 ;
      RECT 5.935000  0.395000 6.105000 0.565000 ;
      RECT 6.095000  3.505000 6.265000 3.675000 ;
      RECT 6.295000  0.395000 6.465000 0.565000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.985000 6.565000 4.155000 ;
      RECT 6.455000  3.505000 6.625000 3.675000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.985000 7.045000 4.155000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.600000  3.505000 7.770000 3.675000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 7.960000  3.505000 8.130000 3.675000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.985000 8.485000 4.155000 ;
      RECT 8.320000  3.505000 8.490000 3.675000 ;
      RECT 8.330000  0.395000 8.500000 0.565000 ;
      RECT 8.690000  0.395000 8.860000 0.565000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.985000 8.965000 4.155000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.985000 9.445000 4.155000 ;
  END
END sky130_fd_sc_hvl__dlrtp_1
