* File: sky130_fd_sc_hvl__o21a_1.pex.spice
* Created: Wed Sep  2 09:08:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__O21A_1%VNB 5 7 11 25
r33 7 25 2.89352e-05 $w=4.32e-06 $l=1e-09 $layer=MET1_cond $X=2.16 $Y=0.057
+ $X2=2.16 $Y2=0.058
r34 7 11 0.00164931 $w=4.32e-06 $l=5.7e-08 $layer=MET1_cond $X=2.16 $Y=0.057
+ $X2=2.16 $Y2=0
r35 5 11 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r36 5 11 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__O21A_1%VPB 4 6 14 21
r34 10 21 0.00164931 $w=4.32e-06 $l=5.7e-08 $layer=MET1_cond $X=2.16 $Y=4.07
+ $X2=2.16 $Y2=4.013
r35 10 14 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=4.07
+ $X2=4.08 $Y2=4.07
r36 9 14 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=4.08 $Y2=4.07
r37 9 10 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r38 6 21 2.89352e-05 $w=4.32e-06 $l=1e-09 $layer=MET1_cond $X=2.16 $Y=4.012
+ $X2=2.16 $Y2=4.013
r39 4 14 40.4444 $w=1.7e-07 $l=4.12228e-06 $layer=licon1_NTAP_notbjt $count=4
+ $X=0 $Y=3.985 $X2=4.08 $Y2=4.07
r40 4 9 40.4444 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=4
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__O21A_1%A_83_87# 1 2 9 13 15 19 21 25 29 33 35
c59 19 0 1.22012e-19 $X=1.66 $Y=0.66
r60 33 38 37.1177 $w=7.35e-07 $l=4.55e-07 $layer=POLY_cond $X=0.782 $Y=1.63
+ $X2=0.782 $Y2=2.085
r61 33 37 8.43598 $w=7.35e-07 $l=4.5e-08 $layer=POLY_cond $X=0.782 $Y=1.63
+ $X2=0.782 $Y2=1.585
r62 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.63 $X2=0.67 $Y2=1.63
r63 29 32 3.63929 $w=2.83e-07 $l=9e-08 $layer=LI1_cond $X=0.692 $Y=1.54
+ $X2=0.692 $Y2=1.63
r64 25 27 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.29 $Y=2.34
+ $X2=2.29 $Y2=3.59
r65 23 25 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.29 $Y=1.625
+ $X2=2.29 $Y2=2.34
r66 22 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=1.54
+ $X2=1.66 $Y2=1.54
r67 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.205 $Y=1.54
+ $X2=2.29 $Y2=1.625
r68 21 22 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.205 $Y=1.54
+ $X2=1.825 $Y2=1.54
r69 17 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=1.455
+ $X2=1.66 $Y2=1.54
r70 17 19 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=1.66 $Y=1.455
+ $X2=1.66 $Y2=0.66
r71 16 29 3.76007 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=0.835 $Y=1.54
+ $X2=0.692 $Y2=1.54
r72 15 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=1.54
+ $X2=1.66 $Y2=1.54
r73 15 16 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.495 $Y=1.54
+ $X2=0.835 $Y2=1.54
r74 13 38 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.9 $Y=2.965 $X2=0.9
+ $Y2=2.085
r75 9 37 69.0188 $w=5e-07 $l=6.45e-07 $layer=POLY_cond $X=0.665 $Y=0.94
+ $X2=0.665 $Y2=1.585
r76 2 27 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.15
+ $Y=2.215 $X2=2.29 $Y2=3.59
r77 2 25 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.15
+ $Y=2.215 $X2=2.29 $Y2=2.34
r78 1 19 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.515
+ $Y=0.535 $X2=1.66 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__O21A_1%B1 3 7 9 10 14 15
r36 14 17 19.0369 $w=6.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.975 $Y=1.89
+ $X2=1.975 $Y2=2.085
r37 14 16 42.0843 $w=6.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.975 $Y=1.89
+ $X2=1.975 $Y2=1.415
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.835
+ $Y=1.89 $X2=1.835 $Y2=1.89
r39 10 15 5.67075 $w=3.13e-07 $l=1.55e-07 $layer=LI1_cond $X=1.68 $Y=1.962
+ $X2=1.835 $Y2=1.962
r40 9 10 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.962 $X2=1.68
+ $Y2=1.962
r41 7 16 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.05 $Y=0.91 $X2=2.05
+ $Y2=1.415
r42 3 17 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.9 $Y=2.965 $X2=1.9
+ $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_HVL__O21A_1%A2 3 7 9 10 11 12 13 20
c35 20 0 1.22012e-19 $X=2.695 $Y=1.715
r36 20 23 19.7175 $w=5.7e-07 $l=2e-07 $layer=POLY_cond $X=2.795 $Y=1.715
+ $X2=2.795 $Y2=1.915
r37 20 22 29.104 $w=5.7e-07 $l=3e-07 $layer=POLY_cond $X=2.795 $Y=1.715
+ $X2=2.795 $Y2=1.415
r38 12 13 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.67 $Y=2.775
+ $X2=2.67 $Y2=3.145
r39 11 12 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.67 $Y=2.405
+ $X2=2.67 $Y2=2.775
r40 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.67 $Y=2.035
+ $X2=2.67 $Y2=2.405
r41 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.67 $Y=1.665
+ $X2=2.67 $Y2=2.035
r42 9 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.695
+ $Y=1.715 $X2=2.695 $Y2=1.715
r43 7 22 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.83 $Y=0.91 $X2=2.83
+ $Y2=1.415
r44 3 23 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.76 $Y=2.965 $X2=2.76
+ $Y2=1.915
.ends

.subckt PM_SKY130_FD_SC_HVL__O21A_1%A1 3 7 9 10 11 16
r26 16 19 39.0327 $w=5.9e-07 $l=4.15e-07 $layer=POLY_cond $X=3.585 $Y=1.67
+ $X2=3.585 $Y2=2.085
r27 16 18 24.5235 $w=5.9e-07 $l=2.55e-07 $layer=POLY_cond $X=3.585 $Y=1.67
+ $X2=3.585 $Y2=1.415
r28 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.475
+ $Y=1.67 $X2=3.475 $Y2=1.67
r29 10 11 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.67 $X2=4.08
+ $Y2=1.67
r30 10 17 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.6 $Y=1.67
+ $X2=3.475 $Y2=1.67
r31 9 17 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.12 $Y=1.67
+ $X2=3.475 $Y2=1.67
r32 7 18 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.63 $Y=0.91 $X2=3.63
+ $Y2=1.415
r33 3 19 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.54 $Y=2.965 $X2=3.54
+ $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_HVL__O21A_1%X 1 2 7 8 9 10 11 12 13 24 35 46
r19 46 47 4.01275 $w=4.68e-07 $l=6e-08 $layer=LI1_cond $X=0.36 $Y=2.035 $X2=0.36
+ $Y2=1.975
r20 33 35 3.3083 $w=4.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.36 $Y=2.21 $X2=0.36
+ $Y2=2.34
r21 13 43 11.3246 $w=4.68e-07 $l=4.45e-07 $layer=LI1_cond $X=0.36 $Y=3.145
+ $X2=0.36 $Y2=3.59
r22 12 13 9.41594 $w=4.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.36 $Y=2.775
+ $X2=0.36 $Y2=3.145
r23 11 12 9.41594 $w=4.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.36 $Y=2.405
+ $X2=0.36 $Y2=2.775
r24 11 35 1.65415 $w=4.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.36 $Y=2.405
+ $X2=0.36 $Y2=2.34
r25 10 33 4.1481 $w=4.68e-07 $l=1.63e-07 $layer=LI1_cond $X=0.36 $Y=2.047
+ $X2=0.36 $Y2=2.21
r26 10 46 0.305382 $w=4.68e-07 $l=1.2e-08 $layer=LI1_cond $X=0.36 $Y=2.047
+ $X2=0.36 $Y2=2.035
r27 10 47 0.58752 $w=2.53e-07 $l=1.3e-08 $layer=LI1_cond $X=0.252 $Y=1.962
+ $X2=0.252 $Y2=1.975
r28 9 10 13.4226 $w=2.53e-07 $l=2.97e-07 $layer=LI1_cond $X=0.252 $Y=1.665
+ $X2=0.252 $Y2=1.962
r29 8 9 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=1.295
+ $X2=0.252 $Y2=1.665
r30 7 8 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=0.925
+ $X2=0.252 $Y2=1.295
r31 7 24 9.71668 $w=2.53e-07 $l=2.15e-07 $layer=LI1_cond $X=0.252 $Y=0.925
+ $X2=0.252 $Y2=0.71
r32 2 43 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.365
+ $Y=2.215 $X2=0.51 $Y2=3.59
r33 2 35 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.365
+ $Y=2.215 $X2=0.51 $Y2=2.34
r34 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.565 $X2=0.275 $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_HVL__O21A_1%VPWR 1 2 7 10 20 27
r33 24 27 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=3.055 $Y=3.63
+ $X2=4.135 $Y2=3.63
r34 23 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.135 $Y=3.59
+ $X2=4.135 $Y2=3.59
r35 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.055 $Y=3.59
+ $X2=3.055 $Y2=3.59
r36 20 23 12.0553 $w=1.263e-06 $l=1.25e-06 $layer=LI1_cond $X=3.597 $Y=2.34
+ $X2=3.597 $Y2=3.59
r37 14 17 0.414618 $w=3.7e-07 $l=1.08e-06 $layer=MET1_cond $X=0.86 $Y=3.63
+ $X2=1.94 $Y2=3.63
r38 13 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.94 $Y=3.59
+ $X2=1.94 $Y2=3.59
r39 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.86 $Y=3.59
+ $X2=0.86 $Y2=3.59
r40 10 13 11.7608 $w=1.248e-06 $l=1.205e-06 $layer=LI1_cond $X=1.4 $Y=2.385
+ $X2=1.4 $Y2=3.59
r41 7 24 0.343595 $w=3.7e-07 $l=8.95e-07 $layer=MET1_cond $X=2.16 $Y=3.63
+ $X2=3.055 $Y2=3.63
r42 7 17 0.0844592 $w=3.7e-07 $l=2.2e-07 $layer=MET1_cond $X=2.16 $Y=3.63
+ $X2=1.94 $Y2=3.63
r43 2 23 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=3.79
+ $Y=2.215 $X2=3.93 $Y2=3.59
r44 2 20 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=3.79
+ $Y=2.215 $X2=3.93 $Y2=2.34
r45 1 13 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.15
+ $Y=2.215 $X2=1.29 $Y2=3.59
r46 1 10 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=1.15
+ $Y=2.215 $X2=1.29 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_HVL__O21A_1%VGND 1 2 7 10 17 21
r30 18 21 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.87 $Y=0.44
+ $X2=3.59 $Y2=0.44
r31 17 23 3.70112 $w=8.88e-07 $l=2.7e-07 $layer=LI1_cond $X=3.23 $Y=0.48
+ $X2=3.23 $Y2=0.75
r32 17 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.59 $Y=0.48
+ $X2=3.59 $Y2=0.48
r33 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.87 $Y=0.48
+ $X2=2.87 $Y2=0.48
r34 10 14 3.28335 $w=7.63e-07 $l=2.1e-07 $layer=LI1_cond $X=0.932 $Y=0.48
+ $X2=0.932 $Y2=0.69
r35 10 11 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.19 $Y=0.48
+ $X2=1.19 $Y2=0.48
r36 7 18 0.272573 $w=3.7e-07 $l=7.1e-07 $layer=MET1_cond $X=2.16 $Y=0.44
+ $X2=2.87 $Y2=0.44
r37 7 11 0.372388 $w=3.7e-07 $l=9.7e-07 $layer=MET1_cond $X=2.16 $Y=0.44
+ $X2=1.19 $Y2=0.44
r38 2 23 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=3.08
+ $Y=0.535 $X2=3.22 $Y2=0.75
r39 1 14 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.915
+ $Y=0.565 $X2=1.055 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HVL__O21A_1%A_460_107# 1 2 9 11 12 15
r27 13 15 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.02 $Y=1.105
+ $X2=4.02 $Y2=0.66
r28 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.855 $Y=1.19
+ $X2=4.02 $Y2=1.105
r29 11 12 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=3.855 $Y=1.19
+ $X2=2.605 $Y2=1.19
r30 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.44 $Y=1.105
+ $X2=2.605 $Y2=1.19
r31 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.44 $Y=1.105
+ $X2=2.44 $Y2=0.66
r32 2 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.88
+ $Y=0.535 $X2=4.02 $Y2=0.66
r33 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.3
+ $Y=0.535 $X2=2.44 $Y2=0.66
.ends

