* File: sky130_fd_sc_hvl__decap_4.spice
* Created: Wed Sep  2 09:04:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__decap_4.pex.spice"
.subckt sky130_fd_sc_hvl__decap_4  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_s N_VPWR_M1000_g N_VGND_M1000_s N_VNB_M1000_b NHV L=1 W=0.75
+ AD=0.21375 AS=0.19875 PD=2.07 PS=2.03 NRD=0 NRS=0 M=1 R=0.75 SA=500000
+ SB=500000 A=0.75 P=3.5 MULT=1
MM1001 N_VPWR_M1001_s N_VGND_M1001_g N_VPWR_M1001_s N_VPB_M1001_b PHV L=1 W=1
+ AD=0.285 AS=0.265 PD=2.57 PS=2.53 NRD=0 NRS=0 M=1 R=1 SA=500000 SB=500000 A=1
+ P=4 MULT=1
DX2_noxref N_VNB_M1000_b N_VPB_M1001_b NWDIODE A=6.708 P=10.36
*
.include "sky130_fd_sc_hvl__decap_4.pxi.spice"
*
.ends
*
*
