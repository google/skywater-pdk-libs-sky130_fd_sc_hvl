* File: sky130_fd_sc_hvl__or2_1.pex.spice
* Created: Fri Aug 28 09:39:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__OR2_1%VNB 5 7 11 25
r22 7 25 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0.058
r23 7 11 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=0.057
+ $X2=1.68 $Y2=0
r24 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r25 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__OR2_1%VPB 4 6 14 21
c19 4 0 1.73032e-19 $X=-0.33 $Y=1.885
r20 10 21 0.00212054 $w=3.36e-06 $l=5.7e-08 $layer=MET1_cond $X=1.68 $Y=4.07
+ $X2=1.68 $Y2=4.013
r21 10 14 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=4.07
+ $X2=3.12 $Y2=4.07
r22 9 14 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=3.12 $Y2=4.07
r23 9 10 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r24 6 21 3.72024e-05 $w=3.36e-06 $l=1e-09 $layer=MET1_cond $X=1.68 $Y=4.012
+ $X2=1.68 $Y2=4.013
r25 4 14 52 $w=1.7e-07 $l=3.16221e-06 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=3.12 $Y2=4.07
r26 4 9 52 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__OR2_1%B 3 7 9 12
r28 12 15 47.4652 $w=6.2e-07 $l=5.25e-07 $layer=POLY_cond $X=0.895 $Y=1.28
+ $X2=0.895 $Y2=1.805
r29 12 14 18.9878 $w=6.2e-07 $l=1.95e-07 $layer=POLY_cond $X=0.895 $Y=1.28
+ $X2=0.895 $Y2=1.085
r30 9 12 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.77 $Y=1.28
+ $X2=0.77 $Y2=1.28
r31 7 15 66.3437 $w=5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.955 $Y=2.425
+ $X2=0.955 $Y2=1.805
r32 3 14 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.955 $Y=0.745 $X2=0.955
+ $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_HVL__OR2_1%A 3 7 9 12
r29 12 15 50.2236 $w=5.7e-07 $l=5.25e-07 $layer=POLY_cond $X=1.7 $Y=1.28 $X2=1.7
+ $Y2=1.805
r30 12 14 19.2482 $w=5.7e-07 $l=1.95e-07 $layer=POLY_cond $X=1.7 $Y=1.28 $X2=1.7
+ $Y2=1.085
r31 9 12 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.695
+ $Y=1.28 $X2=1.695 $Y2=1.28
r32 7 14 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.735 $Y=0.745 $X2=1.735
+ $Y2=1.085
r33 3 15 66.3437 $w=5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.665 $Y=2.425
+ $X2=1.665 $Y2=1.805
.ends

.subckt PM_SKY130_FD_SC_HVL__OR2_1%A_84_443# 1 2 9 11 12 15 18 19 21 22 24 30 34
c57 18 0 1.73032e-19 $X=1.265 $Y=1.905
r58 25 34 115.031 $w=5e-07 $l=1.075e-06 $layer=POLY_cond $X=2.675 $Y=1.89
+ $X2=2.675 $Y2=2.965
r59 25 30 104.866 $w=5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.675 $Y=1.89
+ $X2=2.675 $Y2=0.91
r60 24 27 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.61 $Y=1.89 $X2=2.61
+ $Y2=1.99
r61 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.89 $X2=2.61 $Y2=1.89
r62 20 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=1.99
+ $X2=1.265 $Y2=1.99
r63 19 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=1.99
+ $X2=2.61 $Y2=1.99
r64 19 20 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=2.445 $Y=1.99
+ $X2=1.35 $Y2=1.99
r65 18 22 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=1.905
+ $X2=1.265 $Y2=1.99
r66 18 21 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=1.265 $Y=1.905
+ $X2=1.265 $Y2=0.995
r67 13 21 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=0.83
+ $X2=1.345 $Y2=0.995
r68 13 15 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.345 $Y=0.83
+ $X2=1.345 $Y2=0.745
r69 11 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=1.99
+ $X2=1.265 $Y2=1.99
r70 11 12 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.18 $Y=1.99
+ $X2=0.65 $Y2=1.99
r71 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.525 $Y=2.075
+ $X2=0.65 $Y2=1.99
r72 7 9 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=0.525 $Y=2.075
+ $X2=0.525 $Y2=2.425
r73 2 9 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.42
+ $Y=2.215 $X2=0.565 $Y2=2.425
r74 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.205
+ $Y=0.535 $X2=1.345 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__OR2_1%VPWR 1 4 7 16
r19 12 16 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.715 $Y=3.59
+ $X2=2.715 $Y2=3.59
r20 12 13 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.915 $Y=3.59
+ $X2=0.915 $Y2=3.59
r21 10 12 5.17107 $w=1.968e-06 $l=8.35e-07 $layer=LI1_cond $X=1.815 $Y=2.755
+ $X2=1.815 $Y2=3.59
r22 7 10 2.57005 $w=1.968e-06 $l=4.15e-07 $layer=LI1_cond $X=1.815 $Y=2.34
+ $X2=1.815 $Y2=2.755
r23 4 16 0.397342 $w=3.7e-07 $l=1.035e-06 $layer=MET1_cond $X=1.68 $Y=3.63
+ $X2=2.715 $Y2=3.63
r24 4 13 0.293688 $w=3.7e-07 $l=7.65e-07 $layer=MET1_cond $X=1.68 $Y=3.63
+ $X2=0.915 $Y2=3.63
r25 1 12 400 $w=1.7e-07 $l=1.54899e-06 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=2.215 $X2=2.285 $Y2=3.59
r26 1 10 400 $w=1.7e-07 $l=7.00999e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=2.215 $X2=2.285 $Y2=2.755
r27 1 7 600 $w=1.7e-07 $l=4.2796e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=2.215 $X2=2.285 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__OR2_1%X 1 2 7 8 9 10 11 12 13 22
r13 13 40 20.1113 $w=2.53e-07 $l=4.45e-07 $layer=LI1_cond $X=3.107 $Y=3.145
+ $X2=3.107 $Y2=3.59
r14 12 13 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.107 $Y=2.775
+ $X2=3.107 $Y2=3.145
r15 11 12 19.6593 $w=2.53e-07 $l=4.35e-07 $layer=LI1_cond $X=3.107 $Y=2.34
+ $X2=3.107 $Y2=2.775
r16 10 11 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=3.107 $Y=2.035
+ $X2=3.107 $Y2=2.34
r17 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.107 $Y=1.665
+ $X2=3.107 $Y2=2.035
r18 8 9 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.107 $Y=1.295
+ $X2=3.107 $Y2=1.665
r19 7 8 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.107 $Y=0.925
+ $X2=3.107 $Y2=1.295
r20 7 22 11.9764 $w=2.53e-07 $l=2.65e-07 $layer=LI1_cond $X=3.107 $Y=0.925
+ $X2=3.107 $Y2=0.66
r21 2 40 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.925
+ $Y=2.215 $X2=3.065 $Y2=3.59
r22 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.925
+ $Y=2.215 $X2=3.065 $Y2=2.34
r23 1 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.925
+ $Y=0.535 $X2=3.065 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__OR2_1%VGND 1 2 7 10 19 20
r26 23 25 10.1363 $w=5.88e-07 $l=5e-07 $layer=LI1_cond $X=2.335 $Y=0.66
+ $X2=2.335 $Y2=1.16
r27 19 23 3.64905 $w=5.88e-07 $l=1.8e-07 $layer=LI1_cond $X=2.335 $Y=0.48
+ $X2=2.335 $Y2=0.66
r28 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.515 $Y=0.48
+ $X2=2.515 $Y2=0.48
r29 11 14 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.185 $Y=0.44
+ $X2=0.905 $Y2=0.44
r30 10 16 3.55275 $w=9.08e-07 $l=2.65e-07 $layer=LI1_cond $X=0.545 $Y=0.48
+ $X2=0.545 $Y2=0.745
r31 10 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.905 $Y=0.48
+ $X2=0.905 $Y2=0.48
r32 10 11 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.185 $Y=0.48
+ $X2=0.185 $Y2=0.48
r33 7 20 0.320561 $w=3.7e-07 $l=8.35e-07 $layer=MET1_cond $X=1.68 $Y=0.44
+ $X2=2.515 $Y2=0.44
r34 7 14 0.297527 $w=3.7e-07 $l=7.75e-07 $layer=MET1_cond $X=1.68 $Y=0.44
+ $X2=0.905 $Y2=0.44
r35 2 25 182 $w=1.7e-07 $l=7.60345e-07 $layer=licon1_NDIFF $count=1 $X=1.985
+ $Y=0.535 $X2=2.285 $Y2=1.16
r36 2 23 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=1.985
+ $Y=0.535 $X2=2.285 $Y2=0.66
r37 1 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.42
+ $Y=0.535 $X2=0.565 $Y2=0.745
.ends

