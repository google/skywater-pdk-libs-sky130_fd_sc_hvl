# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__xor2_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__xor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  2.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.775000 3.235000 2.150000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.775000 1.510000 2.055000 ;
        RECT 1.340000 1.425000 3.585000 1.505000 ;
        RECT 1.340000 1.505000 3.715000 1.595000 ;
        RECT 1.340000 1.595000 1.510000 1.775000 ;
        RECT 3.415000 1.595000 3.715000 1.835000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.637500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.850000 0.495000 4.370000 1.325000 ;
        RECT 3.965000 1.325000 4.370000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.365000 0.680000 1.245000 ;
        RECT 1.340000 0.365000 3.670000 1.245000 ;
        RECT 4.550000 0.365000 5.140000 1.325000 ;
      LAYER mcon ;
        RECT 0.120000 0.395000 0.290000 0.565000 ;
        RECT 0.480000 0.395000 0.650000 0.565000 ;
        RECT 1.340000 0.395000 1.510000 0.565000 ;
        RECT 1.700000 0.395000 1.870000 0.565000 ;
        RECT 2.060000 0.395000 2.230000 0.565000 ;
        RECT 2.420000 0.395000 2.590000 0.565000 ;
        RECT 2.780000 0.395000 2.950000 0.565000 ;
        RECT 3.140000 0.395000 3.310000 0.565000 ;
        RECT 3.500000 0.395000 3.670000 0.565000 ;
        RECT 4.580000 0.395000 4.750000 0.565000 ;
        RECT 4.940000 0.395000 5.110000 0.565000 ;
      LAYER met1 ;
        RECT 0.000000 0.255000 5.280000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.115000 5.280000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 5.280000 4.155000 ;
      LAYER mcon ;
        RECT 0.155000 3.985000 0.325000 4.155000 ;
        RECT 0.635000 3.985000 0.805000 4.155000 ;
        RECT 1.115000 3.985000 1.285000 4.155000 ;
        RECT 1.595000 3.985000 1.765000 4.155000 ;
        RECT 2.075000 3.985000 2.245000 4.155000 ;
        RECT 2.555000 3.985000 2.725000 4.155000 ;
        RECT 3.035000 3.985000 3.205000 4.155000 ;
        RECT 3.515000 3.985000 3.685000 4.155000 ;
        RECT 3.995000 3.985000 4.165000 4.155000 ;
        RECT 4.475000 3.985000 4.645000 4.155000 ;
        RECT 4.955000 3.985000 5.125000 4.155000 ;
      LAYER met1 ;
        RECT 0.000000 3.955000 5.280000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.560000 2.785000 2.530000 3.755000 ;
        RECT 3.060000 3.305000 4.720000 3.755000 ;
      LAYER mcon ;
        RECT 0.560000 3.505000 0.730000 3.675000 ;
        RECT 0.920000 3.505000 1.090000 3.675000 ;
        RECT 1.280000 3.505000 1.450000 3.675000 ;
        RECT 1.640000 3.505000 1.810000 3.675000 ;
        RECT 2.000000 3.505000 2.170000 3.675000 ;
        RECT 2.360000 3.505000 2.530000 3.675000 ;
        RECT 3.085000 3.505000 3.255000 3.675000 ;
        RECT 3.445000 3.505000 3.615000 3.675000 ;
        RECT 3.805000 3.505000 3.975000 3.675000 ;
        RECT 4.165000 3.505000 4.335000 3.675000 ;
        RECT 4.525000 3.505000 4.695000 3.675000 ;
      LAYER met1 ;
        RECT 0.000000 3.445000 5.280000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.130000 1.425000 1.160000 1.595000 ;
      RECT 0.130000 1.595000 0.380000 2.435000 ;
      RECT 0.130000 2.435000 3.230000 2.605000 ;
      RECT 0.130000 2.605000 0.380000 3.755000 ;
      RECT 0.910000 0.495000 1.160000 1.425000 ;
      RECT 2.710000 2.785000 2.880000 2.955000 ;
      RECT 2.710000 2.955000 5.150000 3.125000 ;
      RECT 2.710000 3.125000 2.880000 3.755000 ;
      RECT 3.060000 2.605000 4.720000 2.775000 ;
      RECT 4.550000 1.665000 4.880000 1.995000 ;
      RECT 4.550000 1.995000 4.720000 2.605000 ;
      RECT 4.900000 2.175000 5.150000 2.955000 ;
      RECT 4.900000 3.125000 5.150000 3.755000 ;
  END
END sky130_fd_sc_hvl__xor2_1
