* File: sky130_fd_sc_hvl__dlclkp_1.spice
* Created: Fri Aug 28 09:34:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__dlclkp_1.pex.spice"
.subckt sky130_fd_sc_hvl__dlclkp_1  VNB VPB GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1002 A_189_159# N_GATE_M1002_g N_VGND_M1002_s N_VNB_M1002_b NHV L=0.5 W=0.42
+ AD=0.0525 AS=0.1239 PD=0.67 PS=1.43 NRD=18.9924 NRS=0 M=1 R=0.84 SA=250000
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1012 N_A_303_311#_M1012_d N_A_231_71#_M1012_g A_189_159# N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.0525 PD=1.37 PS=0.67 NRD=0 NRS=18.9924 M=1 R=0.84
+ SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1017 N_VGND_M1017_d N_A_231_71#_M1017_g N_A_239_419#_M1017_s N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1005 N_A_231_71#_M1005_d N_CLK_M1005_g N_VGND_M1017_d N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250001
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1004 A_1027_159# N_A_239_419#_M1004_g N_A_303_311#_M1004_s N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1009 N_VGND_M1009_d N_A_1069_133#_M1009_g A_1027_159# N_VNB_M1002_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1001 N_A_1069_133#_M1001_d N_A_303_311#_M1001_g N_VGND_M1009_d N_VNB_M1002_b
+ NHV L=0.5 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1015 A_1591_171# N_A_1069_133#_M1015_g N_A_1438_171#_M1015_s N_VNB_M1002_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=23.0622 NRS=0 M=1 R=0.84
+ SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1011 N_VGND_M1011_d N_CLK_M1011_g A_1591_171# N_VNB_M1002_b NHV L=0.5 W=0.42
+ AD=0.0826538 AS=0.0588 PD=0.782564 PS=0.7 NRD=16.2792 NRS=23.0622 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1010 N_GCLK_M1010_d N_A_1438_171#_M1010_g N_VGND_M1011_d N_VNB_M1002_b NHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.147596 PD=2.03 PS=1.39744 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1000 A_189_445# N_GATE_M1000_g N_VPWR_M1000_s N_VPB_M1000_b PHV L=0.5 W=0.75
+ AD=0.09375 AS=0.22125 PD=1 PS=2.09 NRD=17.8203 NRS=0 M=1 R=1.5 SA=250000
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1007 N_A_303_311#_M1007_d N_A_239_419#_M1007_g A_189_445# N_VPB_M1000_b PHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.09375 PD=2.03 PS=1 NRD=0 NRS=17.8203 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1018 N_VPWR_M1018_d N_A_231_71#_M1018_g N_A_239_419#_M1018_s N_VPB_M1000_b PHV
+ L=0.5 W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1006 N_A_231_71#_M1006_d N_CLK_M1006_g N_VPWR_M1018_d N_VPB_M1000_b PHV L=0.5
+ W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5 SA=250001
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1013 A_1027_457# N_A_231_71#_M1013_g N_A_303_311#_M1013_s N_VPB_M1000_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1014 N_VPWR_M1014_d N_A_1069_133#_M1014_g A_1027_457# N_VPB_M1000_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1008 N_A_1069_133#_M1008_d N_A_303_311#_M1008_g N_VPWR_M1014_d N_VPB_M1000_b
+ PHV L=0.5 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1003 N_A_1438_171#_M1003_d N_A_1069_133#_M1003_g N_VPWR_M1003_s N_VPB_M1000_b
+ PHV L=0.5 W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250002 A=0.375 P=2.5 MULT=1
MM1019 N_VPWR_M1019_d N_CLK_M1019_g N_A_1438_171#_M1003_d N_VPB_M1000_b PHV
+ L=0.5 W=0.75 AD=0.15125 AS=0.105 PD=1.22667 PS=1.03 NRD=15.2609 NRS=0 M=1
+ R=1.5 SA=250001 SB=250001 A=0.375 P=2.5 MULT=1
MM1016 N_GCLK_M1016_d N_A_1438_171#_M1016_g N_VPWR_M1019_d N_VPB_M1000_b PHV
+ L=0.5 W=1.5 AD=0.3975 AS=0.3025 PD=3.53 PS=2.45333 NRD=0 NRS=0 M=1 R=3
+ SA=250001 SB=250000 A=0.75 P=4 MULT=1
DX20_noxref N_VNB_M1002_b N_VPB_M1000_b NWDIODE A=27.924 P=26.68
*
.include "sky130_fd_sc_hvl__dlclkp_1.pxi.spice"
*
.ends
*
*
