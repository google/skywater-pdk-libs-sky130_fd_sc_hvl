* File: sky130_fd_sc_hvl__sdfsbp_1.pxi.spice
* Created: Fri Aug 28 09:39:59 2020
* 
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%VNB N_VNB_M1014_b VNB N_VNB_c_2_p
+ PM_SKY130_FD_SC_HVL__SDFSBP_1%VNB
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%VPB N_VPB_M1000_b VPB N_VPB_c_137_p
+ PM_SKY130_FD_SC_HVL__SDFSBP_1%VPB
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%SCE N_SCE_c_308_n N_SCE_M1000_g N_SCE_M1014_g
+ N_SCE_c_310_n N_SCE_M1012_g N_SCE_M1016_g N_SCE_c_300_n N_SCE_c_301_n
+ N_SCE_c_321_p N_SCE_c_341_p N_SCE_c_302_n SCE SCE SCE N_SCE_c_303_n
+ N_SCE_c_304_n N_SCE_c_306_n N_SCE_c_307_n PM_SKY130_FD_SC_HVL__SDFSBP_1%SCE
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%D N_D_M1029_g N_D_c_377_n N_D_M1015_g D
+ N_D_c_393_n PM_SKY130_FD_SC_HVL__SDFSBP_1%D
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%A_30_569# N_A_30_569#_M1014_s
+ N_A_30_569#_M1000_s N_A_30_569#_c_422_n N_A_30_569#_M1005_g
+ N_A_30_569#_c_415_n N_A_30_569#_c_417_n N_A_30_569#_c_426_n
+ N_A_30_569#_c_427_n N_A_30_569#_c_418_n N_A_30_569#_c_443_n
+ N_A_30_569#_c_419_n N_A_30_569#_c_428_n N_A_30_569#_M1028_g
+ PM_SKY130_FD_SC_HVL__SDFSBP_1%A_30_569#
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%SCD N_SCD_M1006_g N_SCD_c_496_n SCD SCD SCD SCD
+ N_SCD_M1017_g PM_SKY130_FD_SC_HVL__SDFSBP_1%SCD
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%CLK N_CLK_M1025_g N_CLK_M1001_g CLK CLK CLK
+ N_CLK_c_531_n PM_SKY130_FD_SC_HVL__SDFSBP_1%CLK
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%A_1243_116# N_A_1243_116#_M1022_d
+ N_A_1243_116#_M1011_d N_A_1243_116#_M1004_g N_A_1243_116#_M1041_g
+ N_A_1243_116#_c_586_n N_A_1243_116#_c_587_n N_A_1243_116#_M1020_g
+ N_A_1243_116#_c_588_n N_A_1243_116#_c_567_n N_A_1243_116#_c_589_n
+ N_A_1243_116#_c_590_n N_A_1243_116#_c_568_n N_A_1243_116#_c_570_n
+ N_A_1243_116#_c_572_n N_A_1243_116#_c_651_p N_A_1243_116#_c_574_n
+ N_A_1243_116#_c_575_n N_A_1243_116#_c_576_n N_A_1243_116#_c_577_n
+ N_A_1243_116#_c_578_n N_A_1243_116#_c_621_p N_A_1243_116#_c_592_n
+ N_A_1243_116#_c_580_n N_A_1243_116#_c_581_n N_A_1243_116#_c_629_p
+ N_A_1243_116#_c_582_n N_A_1243_116#_c_583_n N_A_1243_116#_M1023_g
+ N_A_1243_116#_c_595_n PM_SKY130_FD_SC_HVL__SDFSBP_1%A_1243_116#
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%A_972_569# N_A_972_569#_M1001_d
+ N_A_972_569#_M1025_d N_A_972_569#_M1022_g N_A_972_569#_M1011_g
+ N_A_972_569#_c_743_n N_A_972_569#_c_744_n N_A_972_569#_M1007_g
+ N_A_972_569#_c_745_n N_A_972_569#_c_746_n N_A_972_569#_M1030_g
+ N_A_972_569#_c_762_n N_A_972_569#_M1037_g N_A_972_569#_c_747_n
+ N_A_972_569#_M1008_g N_A_972_569#_c_766_n N_A_972_569#_c_749_n
+ N_A_972_569#_c_751_n N_A_972_569#_c_818_n N_A_972_569#_c_752_n
+ N_A_972_569#_c_768_n N_A_972_569#_c_849_p N_A_972_569#_c_769_n
+ N_A_972_569#_c_771_n N_A_972_569#_c_871_p N_A_972_569#_c_821_n
+ N_A_972_569#_c_824_n N_A_972_569#_c_773_n N_A_972_569#_c_774_n
+ N_A_972_569#_c_753_n N_A_972_569#_c_754_n N_A_972_569#_c_755_n
+ N_A_972_569#_c_837_n N_A_972_569#_c_777_n N_A_972_569#_c_779_n
+ PM_SKY130_FD_SC_HVL__SDFSBP_1%A_972_569#
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%A_1711_94# N_A_1711_94#_M1033_s
+ N_A_1711_94#_M1013_d N_A_1711_94#_M1040_g N_A_1711_94#_c_954_n
+ N_A_1711_94#_c_955_n N_A_1711_94#_c_960_n N_A_1711_94#_c_956_n
+ N_A_1711_94#_c_957_n N_A_1711_94#_c_980_n N_A_1711_94#_M1035_g
+ N_A_1711_94#_c_959_n PM_SKY130_FD_SC_HVL__SDFSBP_1%A_1711_94#
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%A_1513_120# N_A_1513_120#_M1007_d
+ N_A_1513_120#_M1004_d N_A_1513_120#_c_1005_n N_A_1513_120#_M1033_g
+ N_A_1513_120#_M1024_g N_A_1513_120#_c_1009_n N_A_1513_120#_c_1010_n
+ N_A_1513_120#_c_1014_n N_A_1513_120#_c_1015_n N_A_1513_120#_c_1011_n
+ N_A_1513_120#_c_1012_n N_A_1513_120#_c_1018_n N_A_1513_120#_c_1046_n
+ N_A_1513_120#_c_1019_n N_A_1513_120#_M1013_g N_A_1513_120#_M1021_g
+ PM_SKY130_FD_SC_HVL__SDFSBP_1%A_1513_120#
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%SET_B N_SET_B_M1018_g N_SET_B_c_1110_n
+ N_SET_B_c_1111_n N_SET_B_c_1113_n N_SET_B_c_1115_n N_SET_B_c_1160_p
+ N_SET_B_c_1116_n SET_B SET_B SET_B SET_B SET_B N_SET_B_M1038_g N_SET_B_M1010_g
+ N_SET_B_M1031_g N_SET_B_c_1119_n PM_SKY130_FD_SC_HVL__SDFSBP_1%SET_B
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%A_2729_463# N_A_2729_463#_M1027_s
+ N_A_2729_463#_M1002_s N_A_2729_463#_M1039_g N_A_2729_463#_c_1196_n
+ N_A_2729_463#_c_1197_n N_A_2729_463#_c_1194_n N_A_2729_463#_M1009_g
+ PM_SKY130_FD_SC_HVL__SDFSBP_1%A_2729_463#
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%A_2501_543# N_A_2501_543#_M1041_d
+ N_A_2501_543#_M1037_d N_A_2501_543#_M1031_d N_A_2501_543#_c_1238_n
+ N_A_2501_543#_M1027_g N_A_2501_543#_c_1251_n N_A_2501_543#_M1002_g
+ N_A_2501_543#_M1026_g N_A_2501_543#_c_1252_n N_A_2501_543#_M1036_g
+ N_A_2501_543#_c_1241_n N_A_2501_543#_c_1242_n N_A_2501_543#_M1034_g
+ N_A_2501_543#_M1032_g N_A_2501_543#_c_1244_n N_A_2501_543#_c_1245_n
+ N_A_2501_543#_c_1260_n N_A_2501_543#_c_1263_n N_A_2501_543#_c_1264_n
+ N_A_2501_543#_c_1246_n N_A_2501_543#_c_1247_n N_A_2501_543#_c_1265_n
+ N_A_2501_543#_c_1248_n N_A_2501_543#_c_1267_n N_A_2501_543#_c_1268_n
+ N_A_2501_543#_c_1327_n N_A_2501_543#_c_1308_n N_A_2501_543#_c_1249_n
+ N_A_2501_543#_c_1250_n N_A_2501_543#_c_1270_n
+ PM_SKY130_FD_SC_HVL__SDFSBP_1%A_2501_543#
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%A_3609_173# N_A_3609_173#_M1034_s
+ N_A_3609_173#_M1032_s N_A_3609_173#_c_1378_n N_A_3609_173#_c_1383_n
+ N_A_3609_173#_c_1379_n N_A_3609_173#_c_1380_n N_A_3609_173#_c_1398_n
+ N_A_3609_173#_M1003_g N_A_3609_173#_M1019_g
+ PM_SKY130_FD_SC_HVL__SDFSBP_1%A_3609_173#
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%VPWR N_VPWR_M1000_d N_VPWR_M1006_d
+ N_VPWR_M1011_s N_VPWR_M1035_d N_VPWR_M1018_d N_VPWR_M1039_d N_VPWR_M1002_d
+ N_VPWR_M1032_d VPWR N_VPWR_c_1419_n N_VPWR_c_1422_n N_VPWR_c_1425_n
+ N_VPWR_c_1428_n N_VPWR_c_1431_n N_VPWR_c_1434_n N_VPWR_c_1437_n
+ N_VPWR_c_1440_n N_VPWR_c_1443_n PM_SKY130_FD_SC_HVL__SDFSBP_1%VPWR
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%A_485_569# N_A_485_569#_M1028_d
+ N_A_485_569#_M1007_s N_A_485_569#_M1015_d N_A_485_569#_M1004_s
+ N_A_485_569#_c_1583_n N_A_485_569#_c_1537_n N_A_485_569#_c_1544_n
+ N_A_485_569#_c_1538_n N_A_485_569#_c_1546_n N_A_485_569#_c_1606_n
+ N_A_485_569#_c_1547_n N_A_485_569#_c_1550_n N_A_485_569#_c_1553_n
+ N_A_485_569#_c_1554_n N_A_485_569#_c_1555_n N_A_485_569#_c_1556_n
+ N_A_485_569#_c_1557_n N_A_485_569#_c_1560_n N_A_485_569#_c_1539_n
+ N_A_485_569#_c_1563_n N_A_485_569#_c_1564_n N_A_485_569#_c_1565_n
+ N_A_485_569#_c_1540_n N_A_485_569#_c_1566_n N_A_485_569#_c_1542_n
+ N_A_485_569#_c_1543_n PM_SKY130_FD_SC_HVL__SDFSBP_1%A_485_569#
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%Q_N N_Q_N_M1026_d N_Q_N_M1036_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_1685_n PM_SKY130_FD_SC_HVL__SDFSBP_1%Q_N
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%Q N_Q_M1003_d N_Q_M1019_d Q Q Q Q Q Q Q
+ N_Q_c_1704_n Q Q PM_SKY130_FD_SC_HVL__SDFSBP_1%Q
x_PM_SKY130_FD_SC_HVL__SDFSBP_1%VGND N_VGND_M1014_d N_VGND_M1017_d
+ N_VGND_M1022_s N_VGND_M1040_d N_VGND_M1038_d N_VGND_M1010_d N_VGND_M1027_d
+ N_VGND_M1034_d VGND N_VGND_c_1719_n N_VGND_c_1721_n N_VGND_c_1723_n
+ N_VGND_c_1725_n N_VGND_c_1727_n N_VGND_c_1729_n N_VGND_c_1731_n
+ N_VGND_c_1733_n N_VGND_c_1735_n PM_SKY130_FD_SC_HVL__SDFSBP_1%VGND
cc_1 N_VNB_M1014_b N_SCE_M1014_g 0.0472327f $X=-0.33 $Y=-0.265 $X2=0.71
+ $Y2=0.745
cc_2 N_VNB_c_2_p N_SCE_M1014_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.71 $Y2=0.745
cc_3 N_VNB_M1014_b N_SCE_c_300_n 0.0273407f $X=-0.33 $Y=-0.265 $X2=0.697
+ $Y2=1.347
cc_4 N_VNB_M1014_b N_SCE_c_301_n 0.0225519f $X=-0.33 $Y=-0.265 $X2=2.68 $Y2=1.58
cc_5 N_VNB_M1014_b N_SCE_c_302_n 0.0777083f $X=-0.33 $Y=-0.265 $X2=2.845
+ $Y2=1.26
cc_6 N_VNB_M1014_b N_SCE_c_303_n 0.0518864f $X=-0.33 $Y=-0.265 $X2=0.775
+ $Y2=1.66
cc_7 N_VNB_M1014_b N_SCE_c_304_n 0.0450892f $X=-0.33 $Y=-0.265 $X2=2.945
+ $Y2=1.075
cc_8 N_VNB_c_2_p N_SCE_c_304_n 0.0023273f $X=0.24 $Y=0 $X2=2.945 $Y2=1.075
cc_9 N_VNB_M1014_b N_SCE_c_306_n 0.0026855f $X=-0.33 $Y=-0.265 $X2=1.46 $Y2=1.83
cc_10 N_VNB_M1014_b N_SCE_c_307_n 0.0015457f $X=-0.33 $Y=-0.265 $X2=1.795
+ $Y2=1.83
cc_11 N_VNB_M1014_b N_D_M1029_g 0.0943246f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=3.055
cc_12 N_VNB_c_2_p N_D_M1029_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.685 $Y2=3.055
cc_13 N_VNB_M1014_b N_D_c_377_n 0.0478876f $X=-0.33 $Y=-0.265 $X2=0.71 $Y2=0.745
cc_14 N_VNB_M1014_b N_A_30_569#_c_415_n 0.0329725f $X=-0.33 $Y=-0.265 $X2=2.98
+ $Y2=0.745
cc_15 N_VNB_c_2_p N_A_30_569#_c_415_n 8.78606e-19 $X=0.24 $Y=0 $X2=2.98
+ $Y2=0.745
cc_16 N_VNB_M1014_b N_A_30_569#_c_417_n 0.0271312f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.527
cc_17 N_VNB_M1014_b N_A_30_569#_c_418_n 0.0098122f $X=-0.33 $Y=-0.265 $X2=2.817
+ $Y2=1.26
cc_18 N_VNB_M1014_b N_A_30_569#_c_419_n 0.0154754f $X=-0.33 $Y=-0.265 $X2=1.115
+ $Y2=1.58
cc_19 N_VNB_M1014_b N_A_30_569#_M1028_g 0.0914859f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_20 N_VNB_c_2_p N_A_30_569#_M1028_g 0.0023273f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_21 N_VNB_M1014_b N_SCD_M1017_g 0.126487f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_22 N_VNB_c_2_p N_SCD_M1017_g 0.00200614f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_23 N_VNB_M1014_b N_CLK_M1001_g 0.0830034f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_24 N_VNB_c_2_p N_CLK_M1001_g 5.86481e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_25 N_VNB_M1014_b CLK 0.0036886f $X=-0.33 $Y=-0.265 $X2=1.465 $Y2=3.055
cc_26 N_VNB_M1014_b N_CLK_c_531_n 0.0452313f $X=-0.33 $Y=-0.265 $X2=0.685
+ $Y2=2.527
cc_27 N_VNB_M1014_b N_A_1243_116#_M1041_g 0.0599235f $X=-0.33 $Y=-0.265 $X2=2.98
+ $Y2=0.745
cc_28 N_VNB_M1014_b N_A_1243_116#_c_567_n 0.00495813f $X=-0.33 $Y=-0.265
+ $X2=2.817 $Y2=1.495
cc_29 N_VNB_M1014_b N_A_1243_116#_c_568_n 0.0518925f $X=-0.33 $Y=-0.265
+ $X2=2.845 $Y2=1.6
cc_30 N_VNB_c_2_p N_A_1243_116#_c_568_n 0.00211002f $X=0.24 $Y=0 $X2=2.845
+ $Y2=1.6
cc_31 N_VNB_M1014_b N_A_1243_116#_c_570_n 0.0294281f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=1.58
cc_32 N_VNB_c_2_p N_A_1243_116#_c_570_n 0.00124361f $X=0.24 $Y=0 $X2=0.635
+ $Y2=1.58
cc_33 N_VNB_M1014_b N_A_1243_116#_c_572_n 0.0699225f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_c_2_p N_A_1243_116#_c_572_n 0.00289338f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_35 N_VNB_M1014_b N_A_1243_116#_c_574_n 0.00118725f $X=-0.33 $Y=-0.265
+ $X2=2.945 $Y2=1.075
cc_36 N_VNB_M1014_b N_A_1243_116#_c_575_n 0.00110987f $X=-0.33 $Y=-0.265
+ $X2=1.46 $Y2=1.83
cc_37 N_VNB_M1014_b N_A_1243_116#_c_576_n 0.0064362f $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=1.83
cc_38 N_VNB_M1014_b N_A_1243_116#_c_577_n 0.00408767f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_39 N_VNB_M1014_b N_A_1243_116#_c_578_n 0.0122675f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_c_2_p N_A_1243_116#_c_578_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_41 N_VNB_M1014_b N_A_1243_116#_c_580_n 7.39867e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_42 N_VNB_M1014_b N_A_1243_116#_c_581_n 5.63679e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_M1014_b N_A_1243_116#_c_582_n 0.0348534f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_44 N_VNB_M1014_b N_A_1243_116#_c_583_n 0.0334498f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_45 N_VNB_M1014_b N_A_1243_116#_M1023_g 0.0759563f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_c_2_p N_A_1243_116#_M1023_g 5.46696e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_47 N_VNB_M1014_b N_A_972_569#_M1022_g 0.0501079f $X=-0.33 $Y=-0.265 $X2=1.465
+ $Y2=3.055
cc_48 N_VNB_c_2_p N_A_972_569#_M1022_g 0.00102412f $X=0.24 $Y=0 $X2=1.465
+ $Y2=3.055
cc_49 N_VNB_M1014_b N_A_972_569#_c_743_n 0.069673f $X=-0.33 $Y=-0.265 $X2=0.697
+ $Y2=1.085
cc_50 N_VNB_M1014_b N_A_972_569#_c_744_n 0.0403719f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_51 N_VNB_M1014_b N_A_972_569#_c_745_n 0.0194796f $X=-0.33 $Y=-0.265 $X2=1.465
+ $Y2=2.527
cc_52 N_VNB_M1014_b N_A_972_569#_c_746_n 0.0208283f $X=-0.33 $Y=-0.265 $X2=2.68
+ $Y2=1.58
cc_53 N_VNB_M1014_b N_A_972_569#_c_747_n 0.0597329f $X=-0.33 $Y=-0.265 $X2=2.817
+ $Y2=1.63
cc_54 N_VNB_M1014_b N_A_972_569#_M1008_g 0.0403779f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_55 N_VNB_M1014_b N_A_972_569#_c_749_n 0.0321032f $X=-0.33 $Y=-0.265 $X2=1.46
+ $Y2=1.83
cc_56 N_VNB_c_2_p N_A_972_569#_c_749_n 5.64934e-19 $X=0.24 $Y=0 $X2=1.46
+ $Y2=1.83
cc_57 N_VNB_M1014_b N_A_972_569#_c_751_n 0.0288914f $X=-0.33 $Y=-0.265 $X2=1.2
+ $Y2=1.83
cc_58 N_VNB_M1014_b N_A_972_569#_c_752_n 0.0898492f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_59 N_VNB_M1014_b N_A_972_569#_c_753_n 0.0401812f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_60 N_VNB_M1014_b N_A_972_569#_c_754_n 3.99406e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_61 N_VNB_M1014_b N_A_972_569#_c_755_n 0.00369815f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_62 N_VNB_M1014_b N_A_1711_94#_c_954_n 0.00793101f $X=-0.33 $Y=-0.265
+ $X2=1.465 $Y2=3.055
cc_63 N_VNB_M1014_b N_A_1711_94#_c_955_n 0.0513454f $X=-0.33 $Y=-0.265 $X2=2.98
+ $Y2=0.745
cc_64 N_VNB_M1014_b N_A_1711_94#_c_956_n 0.0372385f $X=-0.33 $Y=-0.265 $X2=0.697
+ $Y2=2.527
cc_65 N_VNB_M1014_b N_A_1711_94#_c_957_n 0.0170417f $X=-0.33 $Y=-0.265 $X2=2.68
+ $Y2=1.58
cc_66 N_VNB_c_2_p N_A_1711_94#_c_957_n 7.98897e-19 $X=0.24 $Y=0 $X2=2.68
+ $Y2=1.58
cc_67 N_VNB_M1014_b N_A_1711_94#_c_959_n 0.0392201f $X=-0.33 $Y=-0.265 $X2=1.595
+ $Y2=1.58
cc_68 N_VNB_M1014_b N_A_1513_120#_c_1005_n 0.108933f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_69 N_VNB_c_2_p N_A_1513_120#_c_1005_n 0.0023273f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_70 N_VNB_M1014_b N_A_1513_120#_M1024_g 0.0889337f $X=-0.33 $Y=-0.265 $X2=2.98
+ $Y2=0.745
cc_71 N_VNB_c_2_p N_A_1513_120#_M1024_g 0.00221559f $X=0.24 $Y=0 $X2=2.98
+ $Y2=0.745
cc_72 N_VNB_M1014_b N_A_1513_120#_c_1009_n 0.00661095f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_73 N_VNB_M1014_b N_A_1513_120#_c_1010_n 0.00683f $X=-0.33 $Y=-0.265 $X2=1.795
+ $Y2=1.58
cc_74 N_VNB_M1014_b N_A_1513_120#_c_1011_n 0.0412199f $X=-0.33 $Y=-0.265
+ $X2=0.635 $Y2=1.58
cc_75 N_VNB_M1014_b N_A_1513_120#_c_1012_n 0.00219915f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_76 N_VNB_M1014_b N_SET_B_c_1110_n 0.055653f $X=-0.33 $Y=-0.265 $X2=0.71
+ $Y2=0.745
cc_77 N_VNB_M1014_b N_SET_B_c_1111_n 0.14282f $X=-0.33 $Y=-0.265 $X2=0.71
+ $Y2=0.745
cc_78 N_VNB_c_2_p N_SET_B_c_1111_n 0.00611967f $X=0.24 $Y=0 $X2=0.71 $Y2=0.745
cc_79 N_VNB_M1014_b N_SET_B_c_1113_n 0.0139229f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_80 N_VNB_c_2_p N_SET_B_c_1113_n 5.63772e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_81 N_VNB_M1014_b N_SET_B_c_1115_n 0.00594111f $X=-0.33 $Y=-0.265 $X2=1.465
+ $Y2=3.055
cc_82 N_VNB_M1014_b N_SET_B_c_1116_n 0.0056681f $X=-0.33 $Y=-0.265 $X2=2.98
+ $Y2=0.745
cc_83 N_VNB_M1014_b N_SET_B_M1038_g 0.0656929f $X=-0.33 $Y=-0.265 $X2=2.817
+ $Y2=1.63
cc_84 N_VNB_M1014_b N_SET_B_M1010_g 0.0811735f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_85 N_VNB_M1014_b N_SET_B_c_1119_n 0.0107167f $X=-0.33 $Y=-0.265 $X2=2.945
+ $Y2=1.26
cc_86 N_VNB_M1014_b N_A_2729_463#_c_1194_n 0.0158387f $X=-0.33 $Y=-0.265
+ $X2=1.465 $Y2=2.527
cc_87 N_VNB_M1014_b N_A_2729_463#_M1009_g 0.079029f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_88 N_VNB_M1014_b N_A_2501_543#_c_1238_n 0.046953f $X=-0.33 $Y=-0.265
+ $X2=1.465 $Y2=3.055
cc_89 N_VNB_M1014_b N_A_2501_543#_M1026_g 0.0686955f $X=-0.33 $Y=-0.265
+ $X2=0.697 $Y2=2.527
cc_90 N_VNB_c_2_p N_A_2501_543#_M1026_g 0.00112176f $X=0.24 $Y=0 $X2=0.697
+ $Y2=2.527
cc_91 N_VNB_M1014_b N_A_2501_543#_c_1241_n 0.0526127f $X=-0.33 $Y=-0.265
+ $X2=1.795 $Y2=1.58
cc_92 N_VNB_M1014_b N_A_2501_543#_c_1242_n 0.0653196f $X=-0.33 $Y=-0.265
+ $X2=2.817 $Y2=1.495
cc_93 N_VNB_M1014_b N_A_2501_543#_M1034_g 0.0657966f $X=-0.33 $Y=-0.265
+ $X2=2.845 $Y2=1.26
cc_94 N_VNB_M1014_b N_A_2501_543#_c_1244_n 0.0859505f $X=-0.33 $Y=-0.265
+ $X2=1.115 $Y2=1.58
cc_95 N_VNB_M1014_b N_A_2501_543#_c_1245_n 0.0218373f $X=-0.33 $Y=-0.265
+ $X2=0.697 $Y2=1.66
cc_96 N_VNB_M1014_b N_A_2501_543#_c_1246_n 0.00769091f $X=-0.33 $Y=-0.265
+ $X2=1.2 $Y2=1.83
cc_97 N_VNB_M1014_b N_A_2501_543#_c_1247_n 0.0109694f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_98 N_VNB_M1014_b N_A_2501_543#_c_1248_n 0.00623834f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_99 N_VNB_M1014_b N_A_2501_543#_c_1249_n 0.00710972f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_100 N_VNB_M1014_b N_A_2501_543#_c_1250_n 4.03932e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_101 N_VNB_M1014_b N_A_3609_173#_c_1378_n 0.0109308f $X=-0.33 $Y=-0.265
+ $X2=1.465 $Y2=3.055
cc_102 N_VNB_M1014_b N_A_3609_173#_c_1379_n 0.0174794f $X=-0.33 $Y=-0.265
+ $X2=0.697 $Y2=1.085
cc_103 N_VNB_M1014_b N_A_3609_173#_c_1380_n 7.73482e-19 $X=-0.33 $Y=-0.265
+ $X2=0.697 $Y2=2.32
cc_104 N_VNB_M1014_b N_A_3609_173#_M1003_g 0.0979482f $X=-0.33 $Y=-0.265
+ $X2=2.817 $Y2=1.495
cc_105 N_VNB_c_2_p N_A_3609_173#_M1003_g 0.00112176f $X=0.24 $Y=0 $X2=2.817
+ $Y2=1.495
cc_106 N_VNB_M1014_b N_A_485_569#_c_1537_n 0.00526154f $X=-0.33 $Y=-0.265
+ $X2=0.697 $Y2=1.085
cc_107 N_VNB_M1014_b N_A_485_569#_c_1538_n 0.00903674f $X=-0.33 $Y=-0.265
+ $X2=1.465 $Y2=2.527
cc_108 N_VNB_M1014_b N_A_485_569#_c_1539_n 0.00270968f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_109 N_VNB_M1014_b N_A_485_569#_c_1540_n 0.0109104f $X=-0.33 $Y=-0.265
+ $X2=1.68 $Y2=1.83
cc_110 N_VNB_c_2_p N_A_485_569#_c_1540_n 8.65969e-19 $X=0.24 $Y=0 $X2=1.68
+ $Y2=1.83
cc_111 N_VNB_M1014_b N_A_485_569#_c_1542_n 0.00201492f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_112 N_VNB_M1014_b N_A_485_569#_c_1543_n 0.00505244f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_113 N_VNB_M1014_b N_Q_N_c_1685_n 0.029591f $X=-0.33 $Y=-0.265 $X2=2.68
+ $Y2=1.58
cc_114 N_VNB_c_2_p N_Q_N_c_1685_n 9.37194e-19 $X=0.24 $Y=0 $X2=2.68 $Y2=1.58
cc_115 N_VNB_M1014_b Q 0.0377143f $X=-0.33 $Y=-0.265 $X2=1.465 $Y2=2.735
cc_116 N_VNB_M1014_b N_Q_c_1704_n 0.033699f $X=-0.33 $Y=-0.265 $X2=2.817
+ $Y2=1.26
cc_117 N_VNB_c_2_p N_Q_c_1704_n 8.31735e-19 $X=0.24 $Y=0 $X2=2.817 $Y2=1.26
cc_118 N_VNB_M1014_b N_VGND_c_1719_n 0.0468651f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_119 N_VNB_c_2_p N_VGND_c_1719_n 0.00269953f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_120 N_VNB_M1014_b N_VGND_c_1721_n 0.0618016f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_121 N_VNB_c_2_p N_VGND_c_1721_n 0.00252324f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_122 N_VNB_M1014_b N_VGND_c_1723_n 0.0501246f $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=1.83
cc_123 N_VNB_c_2_p N_VGND_c_1723_n 0.00166977f $X=0.24 $Y=0 $X2=0.72 $Y2=1.83
cc_124 N_VNB_M1014_b N_VGND_c_1725_n 0.0538695f $X=-0.33 $Y=-0.265 $X2=1.795
+ $Y2=1.83
cc_125 N_VNB_c_2_p N_VGND_c_1725_n 0.00269617f $X=0.24 $Y=0 $X2=1.795 $Y2=1.83
cc_126 N_VNB_M1014_b N_VGND_c_1727_n 0.0508653f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_127 N_VNB_c_2_p N_VGND_c_1727_n 0.00269144f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_128 N_VNB_M1014_b N_VGND_c_1729_n 0.0745564f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_129 N_VNB_c_2_p N_VGND_c_1729_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_130 N_VNB_M1014_b N_VGND_c_1731_n 0.0678664f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_131 N_VNB_c_2_p N_VGND_c_1731_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_132 N_VNB_M1014_b N_VGND_c_1733_n 0.0616735f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_133 N_VNB_c_2_p N_VGND_c_1733_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_134 N_VNB_M1014_b N_VGND_c_1735_n 0.292f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_135 N_VNB_c_2_p N_VGND_c_1735_n 2.15528f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_136 N_VPB_M1000_b N_SCE_c_308_n 0.0408982f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.735
cc_137 N_VPB_c_137_p N_SCE_c_308_n 0.00540119f $X=19.92 $Y=4.07 $X2=0.685
+ $Y2=2.735
cc_138 N_VPB_M1000_b N_SCE_c_310_n 0.128017f $X=-0.33 $Y=1.885 $X2=1.465
+ $Y2=2.735
cc_139 N_VPB_c_137_p N_SCE_c_310_n 0.00386003f $X=19.92 $Y=4.07 $X2=1.465
+ $Y2=2.735
cc_140 N_VPB_M1000_b N_SCE_c_303_n 0.0478111f $X=-0.33 $Y=1.885 $X2=0.775
+ $Y2=1.66
cc_141 N_VPB_M1000_b N_SCE_c_306_n 0.00400406f $X=-0.33 $Y=1.885 $X2=1.46
+ $Y2=1.83
cc_142 N_VPB_M1000_b N_SCE_c_307_n 0.00340924f $X=-0.33 $Y=1.885 $X2=1.795
+ $Y2=1.83
cc_143 N_VPB_M1000_b N_D_c_377_n 0.0502825f $X=-0.33 $Y=1.885 $X2=0.71 $Y2=0.745
cc_144 N_VPB_M1000_b N_D_M1015_g 0.0969052f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_145 N_VPB_c_137_p N_D_M1015_g 0.0110649f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_146 N_VPB_M1000_b N_A_30_569#_c_422_n 0.0750699f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_147 N_VPB_M1000_b N_A_30_569#_M1005_g 0.0396793f $X=-0.33 $Y=1.885 $X2=1.465
+ $Y2=3.055
cc_148 N_VPB_c_137_p N_A_30_569#_M1005_g 0.0110649f $X=19.92 $Y=4.07 $X2=1.465
+ $Y2=3.055
cc_149 N_VPB_M1000_b N_A_30_569#_c_417_n 0.0313698f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.527
cc_150 N_VPB_M1000_b N_A_30_569#_c_426_n 0.0272969f $X=-0.33 $Y=1.885 $X2=0.697
+ $Y2=2.32
cc_151 N_VPB_M1000_b N_A_30_569#_c_427_n 0.0186316f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_152 N_VPB_M1000_b N_A_30_569#_c_428_n 0.0132078f $X=-0.33 $Y=1.885 $X2=1.595
+ $Y2=1.58
cc_153 N_VPB_M1000_b N_SCD_M1006_g 0.0376534f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=3.055
cc_154 N_VPB_c_137_p N_SCD_M1006_g 0.00142985f $X=19.92 $Y=4.07 $X2=0.685
+ $Y2=3.055
cc_155 N_VPB_M1000_b N_SCD_c_496_n 0.0484164f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_156 N_VPB_M1000_b N_SCD_M1017_g 0.0328182f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_157 N_VPB_M1000_b N_CLK_M1025_g 0.0980712f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=3.055
cc_158 VPB N_CLK_M1025_g 6.42549e-19 $X=0 $Y=3.955 $X2=0.685 $Y2=3.055
cc_159 N_VPB_c_137_p N_CLK_M1025_g 0.00512665f $X=19.92 $Y=4.07 $X2=0.685
+ $Y2=3.055
cc_160 N_VPB_M1000_b N_CLK_c_531_n 0.0307829f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=2.527
cc_161 N_VPB_M1000_b N_A_1243_116#_c_586_n 0.0323755f $X=-0.33 $Y=1.885
+ $X2=0.697 $Y2=1.085
cc_162 N_VPB_M1000_b N_A_1243_116#_c_587_n 0.0409681f $X=-0.33 $Y=1.885
+ $X2=0.685 $Y2=2.527
cc_163 N_VPB_M1000_b N_A_1243_116#_c_588_n 0.051161f $X=-0.33 $Y=1.885 $X2=0.697
+ $Y2=2.32
cc_164 N_VPB_M1000_b N_A_1243_116#_c_589_n 0.00253218f $X=-0.33 $Y=1.885
+ $X2=2.845 $Y2=1.26
cc_165 N_VPB_M1000_b N_A_1243_116#_c_590_n 0.00220559f $X=-0.33 $Y=1.885
+ $X2=2.817 $Y2=1.63
cc_166 N_VPB_M1000_b N_A_1243_116#_c_577_n 0.00395637f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_167 N_VPB_M1000_b N_A_1243_116#_c_592_n 0.0513254f $X=-0.33 $Y=1.885 $X2=1.68
+ $Y2=1.83
cc_168 N_VPB_M1000_b N_A_1243_116#_c_580_n 0.00401866f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_169 N_VPB_M1000_b N_A_1243_116#_c_582_n 0.0115079f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_170 N_VPB_M1000_b N_A_1243_116#_c_595_n 0.0411753f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_171 N_VPB_c_137_p N_A_1243_116#_c_595_n 0.00980188f $X=19.92 $Y=4.07 $X2=0
+ $Y2=0
cc_172 N_VPB_M1000_b N_A_972_569#_M1011_g 0.0918482f $X=-0.33 $Y=1.885 $X2=2.98
+ $Y2=0.745
cc_173 N_VPB_c_137_p N_A_972_569#_M1011_g 0.00327509f $X=19.92 $Y=4.07 $X2=2.98
+ $Y2=0.745
cc_174 N_VPB_M1000_b N_A_972_569#_c_745_n 0.0179889f $X=-0.33 $Y=1.885 $X2=1.465
+ $Y2=2.527
cc_175 N_VPB_M1000_b N_A_972_569#_c_746_n 0.0702909f $X=-0.33 $Y=1.885 $X2=2.68
+ $Y2=1.58
cc_176 N_VPB_M1000_b N_A_972_569#_M1030_g 0.0406183f $X=-0.33 $Y=1.885 $X2=2.817
+ $Y2=1.495
cc_177 N_VPB_c_137_p N_A_972_569#_M1030_g 0.0102275f $X=19.92 $Y=4.07 $X2=2.817
+ $Y2=1.495
cc_178 N_VPB_M1000_b N_A_972_569#_c_762_n 0.0404996f $X=-0.33 $Y=1.885 $X2=2.845
+ $Y2=1.26
cc_179 VPB N_A_972_569#_c_762_n 0.00970178f $X=0 $Y=3.955 $X2=2.845 $Y2=1.26
cc_180 N_VPB_c_137_p N_A_972_569#_c_762_n 0.0196751f $X=19.92 $Y=4.07 $X2=2.845
+ $Y2=1.26
cc_181 N_VPB_M1000_b N_A_972_569#_c_747_n 0.023573f $X=-0.33 $Y=1.885 $X2=2.817
+ $Y2=1.63
cc_182 N_VPB_M1000_b N_A_972_569#_c_766_n 0.00942191f $X=-0.33 $Y=1.885
+ $X2=2.945 $Y2=1.26
cc_183 N_VPB_M1000_b N_A_972_569#_c_752_n 0.00599561f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_184 N_VPB_M1000_b N_A_972_569#_c_768_n 0.0148835f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_185 N_VPB_M1000_b N_A_972_569#_c_769_n 0.00805266f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_186 N_VPB_c_137_p N_A_972_569#_c_769_n 0.00784477f $X=19.92 $Y=4.07 $X2=0
+ $Y2=0
cc_187 N_VPB_M1000_b N_A_972_569#_c_771_n 0.00214089f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_188 N_VPB_c_137_p N_A_972_569#_c_771_n 0.00213938f $X=19.92 $Y=4.07 $X2=0
+ $Y2=0
cc_189 N_VPB_M1000_b N_A_972_569#_c_773_n 0.0150032f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_190 N_VPB_M1000_b N_A_972_569#_c_774_n 6.8562e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_191 N_VPB_M1000_b N_A_972_569#_c_753_n 0.0245168f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_192 N_VPB_M1000_b N_A_972_569#_c_754_n 0.0267789f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_193 N_VPB_M1000_b N_A_972_569#_c_777_n 0.00214493f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_194 N_VPB_c_137_p N_A_972_569#_c_777_n 0.00201067f $X=19.92 $Y=4.07 $X2=0
+ $Y2=0
cc_195 N_VPB_M1000_b N_A_972_569#_c_779_n 0.0473702f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_196 N_VPB_M1000_b N_A_1711_94#_c_960_n 0.00942425f $X=-0.33 $Y=1.885
+ $X2=0.697 $Y2=1.085
cc_197 N_VPB_M1000_b N_A_1711_94#_c_956_n 0.102285f $X=-0.33 $Y=1.885 $X2=0.697
+ $Y2=2.527
cc_198 N_VPB_c_137_p N_A_1711_94#_c_956_n 0.00127111f $X=19.92 $Y=4.07 $X2=0.697
+ $Y2=2.527
cc_199 N_VPB_M1000_b N_A_1513_120#_c_1009_n 0.0107304f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_200 N_VPB_M1000_b N_A_1513_120#_c_1014_n 0.0116445f $X=-0.33 $Y=1.885
+ $X2=2.845 $Y2=1.26
cc_201 N_VPB_M1000_b N_A_1513_120#_c_1015_n 0.0260132f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_202 N_VPB_M1000_b N_A_1513_120#_c_1011_n 0.104562f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=1.58
cc_203 N_VPB_c_137_p N_A_1513_120#_c_1011_n 0.00385519f $X=19.92 $Y=4.07
+ $X2=0.635 $Y2=1.58
cc_204 N_VPB_M1000_b N_A_1513_120#_c_1018_n 2.47659e-19 $X=-0.33 $Y=1.885
+ $X2=0.775 $Y2=1.66
cc_205 N_VPB_M1000_b N_A_1513_120#_c_1019_n 0.107619f $X=-0.33 $Y=1.885
+ $X2=2.945 $Y2=1.075
cc_206 VPB N_A_1513_120#_c_1019_n 0.00970178f $X=0 $Y=3.955 $X2=2.945 $Y2=1.075
cc_207 N_VPB_c_137_p N_A_1513_120#_c_1019_n 0.013715f $X=19.92 $Y=4.07 $X2=2.945
+ $Y2=1.075
cc_208 N_VPB_M1000_b N_SET_B_M1018_g 0.0840049f $X=-0.33 $Y=1.885 $X2=0.685
+ $Y2=3.055
cc_209 N_VPB_c_137_p N_SET_B_M1018_g 0.00385587f $X=19.92 $Y=4.07 $X2=0.685
+ $Y2=3.055
cc_210 N_VPB_M1000_b N_SET_B_c_1110_n 0.0375527f $X=-0.33 $Y=1.885 $X2=0.71
+ $Y2=0.745
cc_211 N_VPB_M1000_b N_SET_B_M1010_g 0.114759f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_212 N_VPB_M1000_b N_A_2729_463#_c_1196_n 0.0681922f $X=-0.33 $Y=1.885
+ $X2=2.98 $Y2=0.745
cc_213 N_VPB_M1000_b N_A_2729_463#_c_1197_n 0.0502656f $X=-0.33 $Y=1.885
+ $X2=2.98 $Y2=0.745
cc_214 N_VPB_M1000_b N_A_2729_463#_c_1194_n 0.00372075f $X=-0.33 $Y=1.885
+ $X2=1.465 $Y2=2.527
cc_215 N_VPB_M1000_b N_A_2729_463#_M1009_g 0.0364157f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_216 N_VPB_M1000_b N_A_2501_543#_c_1251_n 0.044232f $X=-0.33 $Y=1.885 $X2=2.98
+ $Y2=0.745
cc_217 N_VPB_M1000_b N_A_2501_543#_c_1252_n 0.0415295f $X=-0.33 $Y=1.885
+ $X2=1.465 $Y2=2.527
cc_218 VPB N_A_2501_543#_c_1252_n 0.00970178f $X=0 $Y=3.955 $X2=1.465 $Y2=2.527
cc_219 N_VPB_c_137_p N_A_2501_543#_c_1252_n 0.0163532f $X=19.92 $Y=4.07
+ $X2=1.465 $Y2=2.527
cc_220 N_VPB_M1000_b N_A_2501_543#_c_1241_n 0.0440107f $X=-0.33 $Y=1.885
+ $X2=1.795 $Y2=1.58
cc_221 N_VPB_M1000_b N_A_2501_543#_c_1242_n 0.0402317f $X=-0.33 $Y=1.885
+ $X2=2.817 $Y2=1.495
cc_222 N_VPB_M1000_b N_A_2501_543#_M1032_g 0.0608791f $X=-0.33 $Y=1.885
+ $X2=2.845 $Y2=1.6
cc_223 N_VPB_M1000_b N_A_2501_543#_c_1244_n 0.0430917f $X=-0.33 $Y=1.885
+ $X2=1.115 $Y2=1.58
cc_224 N_VPB_M1000_b N_A_2501_543#_c_1245_n 0.0162198f $X=-0.33 $Y=1.885
+ $X2=0.697 $Y2=1.66
cc_225 N_VPB_M1000_b N_A_2501_543#_c_1260_n 0.0103385f $X=-0.33 $Y=1.885
+ $X2=2.945 $Y2=1.26
cc_226 VPB N_A_2501_543#_c_1260_n 0.00100531f $X=0 $Y=3.955 $X2=2.945 $Y2=1.26
cc_227 N_VPB_c_137_p N_A_2501_543#_c_1260_n 0.0173323f $X=19.92 $Y=4.07
+ $X2=2.945 $Y2=1.26
cc_228 N_VPB_M1000_b N_A_2501_543#_c_1263_n 0.00810988f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_229 N_VPB_M1000_b N_A_2501_543#_c_1264_n 0.0027431f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_230 N_VPB_M1000_b N_A_2501_543#_c_1265_n 0.00686308f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_231 N_VPB_M1000_b N_A_2501_543#_c_1248_n 0.00418416f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_232 N_VPB_M1000_b N_A_2501_543#_c_1267_n 0.0126423f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_233 N_VPB_M1000_b N_A_2501_543#_c_1268_n 0.0228064f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_234 N_VPB_M1000_b N_A_2501_543#_c_1250_n 7.40541e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_235 N_VPB_M1000_b N_A_2501_543#_c_1270_n 5.73427e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_236 N_VPB_M1000_b N_A_3609_173#_c_1383_n 0.0146799f $X=-0.33 $Y=1.885
+ $X2=2.98 $Y2=0.745
cc_237 N_VPB_M1000_b N_A_3609_173#_M1003_g 0.0834912f $X=-0.33 $Y=1.885
+ $X2=2.817 $Y2=1.495
cc_238 VPB N_A_3609_173#_M1003_g 9.59033e-19 $X=0 $Y=3.955 $X2=2.817 $Y2=1.495
cc_239 N_VPB_c_137_p N_A_3609_173#_M1003_g 0.00514877f $X=19.92 $Y=4.07
+ $X2=2.817 $Y2=1.495
cc_240 N_VPB_M1000_b N_VPWR_c_1419_n 0.0203426f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1419_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_242 N_VPB_c_137_p N_VPWR_c_1419_n 0.0409968f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_243 N_VPB_M1000_b N_VPWR_c_1422_n 0.0187416f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1422_n 0.00252021f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_245 N_VPB_c_137_p N_VPWR_c_1422_n 0.0384021f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_246 N_VPB_M1000_b N_VPWR_c_1425_n 0.0137526f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1425_n 4.76796e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_248 N_VPB_c_137_p N_VPWR_c_1425_n 0.00726526f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_249 N_VPB_M1000_b N_VPWR_c_1428_n 0.031157f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1428_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_251 N_VPB_c_137_p N_VPWR_c_1428_n 0.0409968f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_252 N_VPB_M1000_b N_VPWR_c_1431_n 0.0116835f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1431_n 0.00368247f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_254 N_VPB_c_137_p N_VPWR_c_1431_n 0.0477532f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_255 N_VPB_M1000_b N_VPWR_c_1434_n 0.0342958f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1434_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_257 N_VPB_c_137_p N_VPWR_c_1434_n 0.0409968f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_258 N_VPB_M1000_b N_VPWR_c_1437_n 0.0583754f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1437_n 0.00319522f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_260 N_VPB_c_137_p N_VPWR_c_1437_n 0.0452257f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_261 N_VPB_M1000_b N_VPWR_c_1440_n 0.0385228f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1440_n 0.00269049f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_263 N_VPB_c_137_p N_VPWR_c_1440_n 0.0409968f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_264 N_VPB_M1000_b N_VPWR_c_1443_n 0.351209f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1443_n 2.15393f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_266 N_VPB_c_137_p N_VPWR_c_1443_n 0.111871f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_267 N_VPB_M1000_b N_A_485_569#_c_1544_n 0.00196932f $X=-0.33 $Y=1.885
+ $X2=0.697 $Y2=2.527
cc_268 N_VPB_M1000_b N_A_485_569#_c_1538_n 0.0101195f $X=-0.33 $Y=1.885
+ $X2=1.465 $Y2=2.527
cc_269 N_VPB_M1000_b N_A_485_569#_c_1546_n 0.0276167f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_270 N_VPB_M1000_b N_A_485_569#_c_1547_n 0.0109763f $X=-0.33 $Y=1.885
+ $X2=2.817 $Y2=1.26
cc_271 VPB N_A_485_569#_c_1547_n 0.00290046f $X=0 $Y=3.955 $X2=2.817 $Y2=1.26
cc_272 N_VPB_c_137_p N_A_485_569#_c_1547_n 0.0568137f $X=19.92 $Y=4.07 $X2=2.817
+ $Y2=1.26
cc_273 N_VPB_M1000_b N_A_485_569#_c_1550_n 0.00164055f $X=-0.33 $Y=1.885
+ $X2=2.845 $Y2=1.26
cc_274 VPB N_A_485_569#_c_1550_n 5.70856e-19 $X=0 $Y=3.955 $X2=2.845 $Y2=1.26
cc_275 N_VPB_c_137_p N_A_485_569#_c_1550_n 0.0114989f $X=19.92 $Y=4.07 $X2=2.845
+ $Y2=1.26
cc_276 N_VPB_M1000_b N_A_485_569#_c_1553_n 0.0298346f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_277 N_VPB_M1000_b N_A_485_569#_c_1554_n 0.0141789f $X=-0.33 $Y=1.885
+ $X2=2.817 $Y2=1.63
cc_278 N_VPB_M1000_b N_A_485_569#_c_1555_n 0.00394333f $X=-0.33 $Y=1.885
+ $X2=2.845 $Y2=1.6
cc_279 N_VPB_M1000_b N_A_485_569#_c_1556_n 0.00164977f $X=-0.33 $Y=1.885
+ $X2=0.635 $Y2=1.58
cc_280 N_VPB_M1000_b N_A_485_569#_c_1557_n 0.0270877f $X=-0.33 $Y=1.885
+ $X2=1.115 $Y2=1.58
cc_281 VPB N_A_485_569#_c_1557_n 0.00251245f $X=0 $Y=3.955 $X2=1.115 $Y2=1.58
cc_282 N_VPB_c_137_p N_A_485_569#_c_1557_n 0.0285427f $X=19.92 $Y=4.07 $X2=1.115
+ $Y2=1.58
cc_283 N_VPB_M1000_b N_A_485_569#_c_1560_n 0.00253372f $X=-0.33 $Y=1.885
+ $X2=1.595 $Y2=1.58
cc_284 VPB N_A_485_569#_c_1560_n 3.9e-19 $X=0 $Y=3.955 $X2=1.595 $Y2=1.58
cc_285 N_VPB_c_137_p N_A_485_569#_c_1560_n 0.00456541f $X=19.92 $Y=4.07
+ $X2=1.595 $Y2=1.58
cc_286 N_VPB_M1000_b N_A_485_569#_c_1563_n 0.00782245f $X=-0.33 $Y=1.885
+ $X2=2.945 $Y2=1.26
cc_287 N_VPB_M1000_b N_A_485_569#_c_1564_n 0.00913967f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_288 N_VPB_M1000_b N_A_485_569#_c_1565_n 0.00335007f $X=-0.33 $Y=1.885
+ $X2=1.46 $Y2=1.83
cc_289 N_VPB_M1000_b N_A_485_569#_c_1566_n 0.0028102f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_290 N_VPB_M1000_b N_A_485_569#_c_1543_n 0.0183242f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_291 N_VPB_M1000_b N_Q_N_c_1685_n 0.0242134f $X=-0.33 $Y=1.885 $X2=2.68
+ $Y2=1.58
cc_292 VPB N_Q_N_c_1685_n 0.00125715f $X=0 $Y=3.955 $X2=2.68 $Y2=1.58
cc_293 N_VPB_c_137_p N_Q_N_c_1685_n 0.01807f $X=19.92 $Y=4.07 $X2=2.68 $Y2=1.58
cc_294 N_VPB_M1000_b Q 0.0233716f $X=-0.33 $Y=1.885 $X2=1.465 $Y2=2.735
cc_295 N_VPB_M1000_b Q 0.038437f $X=-0.33 $Y=1.885 $X2=2.98 $Y2=0.745
cc_296 N_VPB_c_137_p Q 0.00532177f $X=19.92 $Y=4.07 $X2=2.98 $Y2=0.745
cc_297 N_VPB_M1000_b Q 0.00979711f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_298 N_SCE_M1014_g N_D_M1029_g 0.0325677f $X=0.71 $Y=0.745 $X2=0 $Y2=0
cc_299 N_SCE_c_306_n N_D_M1029_g 0.00955191f $X=1.46 $Y=1.83 $X2=0 $Y2=0
cc_300 N_SCE_c_307_n N_D_M1029_g 0.0138487f $X=1.795 $Y=1.83 $X2=0 $Y2=0
cc_301 N_SCE_c_310_n N_D_c_377_n 0.0315378f $X=1.465 $Y=2.735 $X2=-0.33
+ $Y2=-0.265
cc_302 N_SCE_c_300_n N_D_c_377_n 0.0325677f $X=0.697 $Y=1.347 $X2=-0.33
+ $Y2=-0.265
cc_303 N_SCE_c_301_n N_D_c_377_n 0.0112044f $X=2.68 $Y=1.58 $X2=-0.33 $Y2=-0.265
cc_304 N_SCE_c_321_p N_D_c_377_n 5.46209e-19 $X=2.817 $Y=1.495 $X2=-0.33
+ $Y2=-0.265
cc_305 N_SCE_c_302_n N_D_c_377_n 0.00647426f $X=2.845 $Y=1.26 $X2=-0.33
+ $Y2=-0.265
cc_306 N_SCE_c_306_n N_D_c_377_n 0.0143304f $X=1.46 $Y=1.83 $X2=-0.33 $Y2=-0.265
cc_307 N_SCE_c_307_n N_D_c_377_n 0.0278831f $X=1.795 $Y=1.83 $X2=-0.33
+ $Y2=-0.265
cc_308 N_SCE_c_310_n N_D_M1015_g 0.0792355f $X=1.465 $Y=2.735 $X2=0 $Y2=0
cc_309 N_SCE_c_307_n N_D_M1015_g 0.0014202f $X=1.795 $Y=1.83 $X2=0 $Y2=0
cc_310 N_SCE_c_310_n N_D_c_393_n 2.39089e-19 $X=1.465 $Y=2.735 $X2=0 $Y2=0
cc_311 N_SCE_c_301_n N_D_c_393_n 0.0245275f $X=2.68 $Y=1.58 $X2=0 $Y2=0
cc_312 N_SCE_c_307_n N_D_c_393_n 0.0245261f $X=1.795 $Y=1.83 $X2=0 $Y2=0
cc_313 N_SCE_c_321_p N_A_30_569#_c_422_n 0.0013231f $X=2.817 $Y=1.495 $X2=0
+ $Y2=0
cc_314 N_SCE_c_302_n N_A_30_569#_c_422_n 0.0376815f $X=2.845 $Y=1.26 $X2=0 $Y2=0
cc_315 N_SCE_M1014_g N_A_30_569#_c_415_n 0.0184667f $X=0.71 $Y=0.745 $X2=0 $Y2=0
cc_316 N_SCE_c_300_n N_A_30_569#_c_415_n 0.0012098f $X=0.697 $Y=1.347 $X2=0
+ $Y2=0
cc_317 N_SCE_c_303_n N_A_30_569#_c_417_n 0.0372171f $X=0.775 $Y=1.66 $X2=19.92
+ $Y2=0
cc_318 N_SCE_c_306_n N_A_30_569#_c_417_n 0.0343665f $X=1.46 $Y=1.83 $X2=19.92
+ $Y2=0
cc_319 N_SCE_c_308_n N_A_30_569#_c_426_n 0.0179965f $X=0.685 $Y=2.735 $X2=0
+ $Y2=0
cc_320 N_SCE_c_310_n N_A_30_569#_c_426_n 0.00203586f $X=1.465 $Y=2.735 $X2=0
+ $Y2=0
cc_321 N_SCE_c_310_n N_A_30_569#_c_427_n 0.0723975f $X=1.465 $Y=2.735 $X2=10.08
+ $Y2=0
cc_322 N_SCE_c_306_n N_A_30_569#_c_427_n 0.0523485f $X=1.46 $Y=1.83 $X2=10.08
+ $Y2=0
cc_323 N_SCE_c_300_n N_A_30_569#_c_418_n 0.0309403f $X=0.697 $Y=1.347 $X2=0
+ $Y2=0
cc_324 N_SCE_c_341_p N_A_30_569#_c_418_n 0.00897033f $X=2.845 $Y=1.26 $X2=0
+ $Y2=0
cc_325 N_SCE_c_302_n N_A_30_569#_c_418_n 6.74062e-19 $X=2.845 $Y=1.26 $X2=0
+ $Y2=0
cc_326 N_SCE_c_306_n N_A_30_569#_c_418_n 0.12666f $X=1.46 $Y=1.83 $X2=0 $Y2=0
cc_327 N_SCE_c_321_p N_A_30_569#_c_443_n 0.0126501f $X=2.817 $Y=1.495 $X2=0
+ $Y2=0
cc_328 N_SCE_c_302_n N_A_30_569#_c_443_n 9.51503e-19 $X=2.845 $Y=1.26 $X2=0
+ $Y2=0
cc_329 N_SCE_c_300_n N_A_30_569#_c_419_n 0.00802441f $X=0.697 $Y=1.347 $X2=0
+ $Y2=0
cc_330 N_SCE_c_310_n N_A_30_569#_c_428_n 0.00513266f $X=1.465 $Y=2.735 $X2=0
+ $Y2=0
cc_331 N_SCE_c_301_n N_A_30_569#_M1028_g 0.0070314f $X=2.68 $Y=1.58 $X2=0 $Y2=0
cc_332 N_SCE_c_341_p N_A_30_569#_M1028_g 0.00205769f $X=2.845 $Y=1.26 $X2=0
+ $Y2=0
cc_333 N_SCE_c_302_n N_A_30_569#_M1028_g 0.0284909f $X=2.845 $Y=1.26 $X2=0 $Y2=0
cc_334 N_SCE_c_304_n N_A_30_569#_M1028_g 0.0149364f $X=2.945 $Y=1.075 $X2=0
+ $Y2=0
cc_335 N_SCE_c_304_n SCD 9.80145e-19 $X=2.945 $Y=1.075 $X2=0 $Y2=0
cc_336 N_SCE_c_304_n N_SCD_M1017_g 0.091583f $X=2.945 $Y=1.075 $X2=19.92 $Y2=0
cc_337 N_SCE_c_308_n N_VPWR_c_1419_n 0.036572f $X=0.685 $Y=2.735 $X2=0 $Y2=0
cc_338 N_SCE_c_310_n N_VPWR_c_1419_n 0.0437251f $X=1.465 $Y=2.735 $X2=0 $Y2=0
cc_339 N_SCE_c_308_n N_VPWR_c_1443_n 0.00697248f $X=0.685 $Y=2.735 $X2=0 $Y2=0
cc_340 N_SCE_c_310_n N_VPWR_c_1443_n 0.00426472f $X=1.465 $Y=2.735 $X2=0 $Y2=0
cc_341 N_SCE_c_341_p N_A_485_569#_c_1537_n 0.0137411f $X=2.845 $Y=1.26 $X2=0
+ $Y2=0
cc_342 N_SCE_c_304_n N_A_485_569#_c_1537_n 0.0291876f $X=2.945 $Y=1.075 $X2=0
+ $Y2=0
cc_343 N_SCE_c_321_p N_A_485_569#_c_1538_n 0.0191228f $X=2.817 $Y=1.495 $X2=0
+ $Y2=0
cc_344 N_SCE_c_341_p N_A_485_569#_c_1538_n 0.0268555f $X=2.845 $Y=1.26 $X2=0
+ $Y2=0
cc_345 N_SCE_c_302_n N_A_485_569#_c_1538_n 0.0211219f $X=2.845 $Y=1.26 $X2=0
+ $Y2=0
cc_346 N_SCE_c_304_n N_A_485_569#_c_1538_n 0.00515904f $X=2.945 $Y=1.075 $X2=0
+ $Y2=0
cc_347 N_SCE_c_310_n N_A_485_569#_c_1565_n 0.0012815f $X=1.465 $Y=2.735 $X2=0
+ $Y2=0
cc_348 N_SCE_c_301_n N_A_485_569#_c_1540_n 0.00725234f $X=2.68 $Y=1.58 $X2=0
+ $Y2=0
cc_349 N_SCE_c_341_p N_A_485_569#_c_1540_n 0.00354615f $X=2.845 $Y=1.26 $X2=0
+ $Y2=0
cc_350 N_SCE_c_302_n N_A_485_569#_c_1540_n 0.00181045f $X=2.845 $Y=1.26 $X2=0
+ $Y2=0
cc_351 N_SCE_c_304_n N_A_485_569#_c_1540_n 0.00822988f $X=2.945 $Y=1.075 $X2=0
+ $Y2=0
cc_352 N_SCE_c_302_n N_A_485_569#_c_1566_n 2.25624e-19 $X=2.845 $Y=1.26 $X2=0
+ $Y2=0
cc_353 N_SCE_M1014_g N_VGND_c_1719_n 0.0317136f $X=0.71 $Y=0.745 $X2=0 $Y2=0
cc_354 N_SCE_c_304_n N_VGND_c_1721_n 0.0016019f $X=2.945 $Y=1.075 $X2=0 $Y2=0
cc_355 N_SCE_M1014_g N_VGND_c_1735_n 0.00595433f $X=0.71 $Y=0.745 $X2=0 $Y2=0
cc_356 N_SCE_c_341_p N_VGND_c_1735_n 7.27719e-19 $X=2.845 $Y=1.26 $X2=0 $Y2=0
cc_357 N_SCE_c_304_n N_VGND_c_1735_n 0.0151014f $X=2.945 $Y=1.075 $X2=0 $Y2=0
cc_358 N_D_c_377_n N_A_30_569#_c_422_n 0.0492808f $X=2.175 $Y=2.11 $X2=0 $Y2=0
cc_359 N_D_c_393_n N_A_30_569#_c_422_n 0.0011898f $X=2.14 $Y=1.93 $X2=0 $Y2=0
cc_360 N_D_M1015_g N_A_30_569#_M1005_g 0.0162433f $X=2.175 $Y=3.055 $X2=0 $Y2=0
cc_361 N_D_c_377_n N_A_30_569#_c_427_n 0.00468852f $X=2.175 $Y=2.11 $X2=10.08
+ $Y2=0
cc_362 N_D_M1015_g N_A_30_569#_c_427_n 0.0445849f $X=2.175 $Y=3.055 $X2=10.08
+ $Y2=0
cc_363 N_D_c_393_n N_A_30_569#_c_427_n 0.0232944f $X=2.14 $Y=1.93 $X2=10.08
+ $Y2=0
cc_364 N_D_M1029_g N_A_30_569#_c_418_n 0.0300401f $X=1.49 $Y=0.745 $X2=0 $Y2=0
cc_365 N_D_c_377_n N_A_30_569#_c_418_n 0.0013667f $X=2.175 $Y=2.11 $X2=0 $Y2=0
cc_366 N_D_c_377_n N_A_30_569#_c_443_n 0.00274965f $X=2.175 $Y=2.11 $X2=0 $Y2=0
cc_367 N_D_c_393_n N_A_30_569#_c_443_n 0.0146634f $X=2.14 $Y=1.93 $X2=0 $Y2=0
cc_368 N_D_M1029_g N_A_30_569#_M1028_g 0.0781539f $X=1.49 $Y=0.745 $X2=0 $Y2=0
cc_369 N_D_c_377_n N_A_30_569#_M1028_g 0.0312173f $X=2.175 $Y=2.11 $X2=0 $Y2=0
cc_370 N_D_M1015_g N_VPWR_c_1419_n 0.0028297f $X=2.175 $Y=3.055 $X2=0 $Y2=0
cc_371 N_D_M1015_g N_VPWR_c_1443_n 0.0169235f $X=2.175 $Y=3.055 $X2=0 $Y2=0
cc_372 N_D_M1015_g N_A_485_569#_c_1544_n 6.50221e-19 $X=2.175 $Y=3.055 $X2=0
+ $Y2=0
cc_373 N_D_M1015_g N_A_485_569#_c_1565_n 0.0115244f $X=2.175 $Y=3.055 $X2=0
+ $Y2=0
cc_374 N_D_M1029_g N_A_485_569#_c_1540_n 0.0014684f $X=1.49 $Y=0.745 $X2=0 $Y2=0
cc_375 N_D_M1029_g N_VGND_c_1719_n 0.0397166f $X=1.49 $Y=0.745 $X2=0 $Y2=0
cc_376 N_D_M1029_g N_VGND_c_1735_n 0.00445548f $X=1.49 $Y=0.745 $X2=0 $Y2=0
cc_377 N_A_30_569#_M1005_g N_SCD_M1006_g 0.0391387f $X=2.955 $Y=3.055 $X2=0
+ $Y2=0
cc_378 N_A_30_569#_c_422_n N_SCD_c_496_n 0.0391387f $X=2.955 $Y=2.715 $X2=0
+ $Y2=0
cc_379 N_A_30_569#_c_422_n N_SCD_M1017_g 0.00820229f $X=2.955 $Y=2.715 $X2=19.92
+ $Y2=0
cc_380 N_A_30_569#_c_426_n N_VPWR_c_1419_n 0.031873f $X=0.295 $Y=3.055 $X2=0
+ $Y2=0
cc_381 N_A_30_569#_c_427_n N_VPWR_c_1419_n 0.0647546f $X=2.635 $Y=2.62 $X2=0
+ $Y2=0
cc_382 N_A_30_569#_M1005_g N_VPWR_c_1422_n 0.00278711f $X=2.955 $Y=3.055 $X2=0
+ $Y2=0
cc_383 N_A_30_569#_M1005_g N_VPWR_c_1443_n 0.0169235f $X=2.955 $Y=3.055 $X2=0
+ $Y2=0
cc_384 N_A_30_569#_c_426_n N_VPWR_c_1443_n 0.0192871f $X=0.295 $Y=3.055 $X2=0
+ $Y2=0
cc_385 N_A_30_569#_M1005_g N_A_485_569#_c_1583_n 0.0274455f $X=2.955 $Y=3.055
+ $X2=0 $Y2=0
cc_386 N_A_30_569#_c_427_n N_A_485_569#_c_1583_n 0.0112889f $X=2.635 $Y=2.62
+ $X2=0 $Y2=0
cc_387 N_A_30_569#_c_422_n N_A_485_569#_c_1544_n 0.00261441f $X=2.955 $Y=2.715
+ $X2=0 $Y2=0
cc_388 N_A_30_569#_M1005_g N_A_485_569#_c_1544_n 0.00580641f $X=2.955 $Y=3.055
+ $X2=0 $Y2=0
cc_389 N_A_30_569#_c_427_n N_A_485_569#_c_1544_n 0.00578689f $X=2.635 $Y=2.62
+ $X2=0 $Y2=0
cc_390 N_A_30_569#_c_422_n N_A_485_569#_c_1538_n 0.0105143f $X=2.955 $Y=2.715
+ $X2=0 $Y2=0
cc_391 N_A_30_569#_c_443_n N_A_485_569#_c_1538_n 0.0233241f $X=2.8 $Y=2.18 $X2=0
+ $Y2=0
cc_392 N_A_30_569#_M1028_g N_A_485_569#_c_1538_n 6.33863e-19 $X=2.2 $Y=0.745
+ $X2=0 $Y2=0
cc_393 N_A_30_569#_c_422_n N_A_485_569#_c_1565_n 0.00173024f $X=2.955 $Y=2.715
+ $X2=0 $Y2=0
cc_394 N_A_30_569#_M1005_g N_A_485_569#_c_1565_n 0.00829232f $X=2.955 $Y=3.055
+ $X2=0 $Y2=0
cc_395 N_A_30_569#_c_427_n N_A_485_569#_c_1565_n 0.0205467f $X=2.635 $Y=2.62
+ $X2=0 $Y2=0
cc_396 N_A_30_569#_M1028_g N_A_485_569#_c_1540_n 0.0116951f $X=2.2 $Y=0.745
+ $X2=0 $Y2=0
cc_397 N_A_30_569#_c_422_n N_A_485_569#_c_1566_n 0.00787334f $X=2.955 $Y=2.715
+ $X2=0 $Y2=0
cc_398 N_A_30_569#_c_427_n N_A_485_569#_c_1566_n 0.00727324f $X=2.635 $Y=2.62
+ $X2=0 $Y2=0
cc_399 N_A_30_569#_c_443_n N_A_485_569#_c_1566_n 0.00594373f $X=2.8 $Y=2.18
+ $X2=0 $Y2=0
cc_400 N_A_30_569#_c_415_n N_VGND_c_1719_n 0.0301109f $X=0.32 $Y=0.745 $X2=0
+ $Y2=0
cc_401 N_A_30_569#_c_418_n N_VGND_c_1719_n 0.0630617f $X=2.135 $Y=1.23 $X2=0
+ $Y2=0
cc_402 N_A_30_569#_M1028_g N_VGND_c_1719_n 0.00362967f $X=2.2 $Y=0.745 $X2=0
+ $Y2=0
cc_403 N_A_30_569#_c_415_n N_VGND_c_1735_n 0.0347613f $X=0.32 $Y=0.745 $X2=0
+ $Y2=0
cc_404 N_A_30_569#_c_418_n N_VGND_c_1735_n 0.0321069f $X=2.135 $Y=1.23 $X2=0
+ $Y2=0
cc_405 N_A_30_569#_M1028_g N_VGND_c_1735_n 0.0212499f $X=2.2 $Y=0.745 $X2=0
+ $Y2=0
cc_406 N_SCD_M1006_g N_CLK_M1025_g 0.0116033f $X=3.665 $Y=3.055 $X2=0 $Y2=0
cc_407 N_SCD_c_496_n N_CLK_M1025_g 0.0207298f $X=3.677 $Y=2.715 $X2=0 $Y2=0
cc_408 SCD N_CLK_M1001_g 0.00146417f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_409 N_SCD_M1017_g N_CLK_M1001_g 0.0227727f $X=3.69 $Y=0.745 $X2=0 $Y2=0
cc_410 N_SCD_M1017_g CLK 0.00979424f $X=3.69 $Y=0.745 $X2=0 $Y2=0
cc_411 SCD N_CLK_c_531_n 0.00305125f $X=3.515 $Y=0.84 $X2=19.92 $Y2=0
cc_412 N_SCD_M1017_g N_CLK_c_531_n 0.0207298f $X=3.69 $Y=0.745 $X2=19.92 $Y2=0
cc_413 N_SCD_M1006_g N_VPWR_c_1422_n 0.0600545f $X=3.665 $Y=3.055 $X2=0 $Y2=0
cc_414 N_SCD_c_496_n N_VPWR_c_1422_n 7.54316e-19 $X=3.677 $Y=2.715 $X2=0 $Y2=0
cc_415 SCD N_A_485_569#_c_1537_n 0.00789052f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_416 N_SCD_M1017_g N_A_485_569#_c_1537_n 0.00152725f $X=3.69 $Y=0.745 $X2=0
+ $Y2=0
cc_417 N_SCD_c_496_n N_A_485_569#_c_1544_n 0.00402193f $X=3.677 $Y=2.715 $X2=0
+ $Y2=0
cc_418 N_SCD_c_496_n N_A_485_569#_c_1538_n 0.00535006f $X=3.677 $Y=2.715 $X2=0
+ $Y2=0
cc_419 SCD N_A_485_569#_c_1538_n 0.0856945f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_420 N_SCD_M1017_g N_A_485_569#_c_1538_n 0.0133535f $X=3.69 $Y=0.745 $X2=0
+ $Y2=0
cc_421 N_SCD_c_496_n N_A_485_569#_c_1546_n 0.0376868f $X=3.677 $Y=2.715
+ $X2=10.08 $Y2=0
cc_422 SCD N_A_485_569#_c_1546_n 0.00966847f $X=3.515 $Y=0.84 $X2=10.08 $Y2=0
cc_423 N_SCD_M1006_g N_A_485_569#_c_1606_n 8.57282e-19 $X=3.665 $Y=3.055 $X2=0
+ $Y2=0
cc_424 N_SCD_c_496_n N_A_485_569#_c_1606_n 4.84789e-19 $X=3.677 $Y=2.715 $X2=0
+ $Y2=0
cc_425 N_SCD_M1006_g N_A_485_569#_c_1565_n 7.66324e-19 $X=3.665 $Y=3.055 $X2=0
+ $Y2=0
cc_426 N_SCD_M1017_g N_A_485_569#_c_1540_n 9.53229e-19 $X=3.69 $Y=0.745 $X2=0
+ $Y2=0
cc_427 SCD N_VGND_c_1721_n 0.0135724f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_428 N_SCD_M1017_g N_VGND_c_1721_n 0.0235381f $X=3.69 $Y=0.745 $X2=0 $Y2=0
cc_429 SCD N_VGND_c_1735_n 0.00983628f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_430 N_SCD_M1017_g N_VGND_c_1735_n 0.0211862f $X=3.69 $Y=0.745 $X2=0 $Y2=0
cc_431 N_CLK_M1025_g N_A_972_569#_c_766_n 0.0131739f $X=4.61 $Y=3.22 $X2=0 $Y2=0
cc_432 N_CLK_c_531_n N_A_972_569#_c_766_n 7.39111e-19 $X=4.545 $Y=1.645 $X2=0
+ $Y2=0
cc_433 N_CLK_M1001_g N_A_972_569#_c_749_n 0.0262096f $X=4.635 $Y=0.745 $X2=0
+ $Y2=0
cc_434 CLK N_A_972_569#_c_749_n 0.0320463f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_435 N_CLK_M1025_g N_A_972_569#_c_754_n 0.0229226f $X=4.61 $Y=3.22 $X2=0 $Y2=0
cc_436 CLK N_A_972_569#_c_754_n 0.0171139f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_437 N_CLK_c_531_n N_A_972_569#_c_754_n 0.00915386f $X=4.545 $Y=1.645 $X2=0
+ $Y2=0
cc_438 CLK N_A_972_569#_c_755_n 0.0114322f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_439 N_CLK_c_531_n N_A_972_569#_c_755_n 0.00520216f $X=4.545 $Y=1.645 $X2=0
+ $Y2=0
cc_440 N_CLK_M1025_g N_VPWR_c_1422_n 0.00404099f $X=4.61 $Y=3.22 $X2=0 $Y2=0
cc_441 N_CLK_M1025_g N_VPWR_c_1443_n 0.0183107f $X=4.61 $Y=3.22 $X2=0 $Y2=0
cc_442 N_CLK_M1025_g N_A_485_569#_c_1546_n 0.0213774f $X=4.61 $Y=3.22 $X2=10.08
+ $Y2=0
cc_443 CLK N_A_485_569#_c_1546_n 0.0139107f $X=4.475 $Y=1.21 $X2=10.08 $Y2=0
cc_444 N_CLK_M1025_g N_A_485_569#_c_1606_n 0.0404712f $X=4.61 $Y=3.22 $X2=0
+ $Y2=0
cc_445 N_CLK_M1025_g N_A_485_569#_c_1547_n 0.0115404f $X=4.61 $Y=3.22 $X2=0
+ $Y2=0
cc_446 N_CLK_M1025_g N_A_485_569#_c_1550_n 0.00484464f $X=4.61 $Y=3.22 $X2=0
+ $Y2=0
cc_447 N_CLK_M1025_g N_A_485_569#_c_1553_n 0.00297941f $X=4.61 $Y=3.22 $X2=0
+ $Y2=0
cc_448 N_CLK_M1001_g N_VGND_c_1721_n 0.0487113f $X=4.635 $Y=0.745 $X2=0 $Y2=0
cc_449 CLK N_VGND_c_1721_n 0.0248918f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_450 N_CLK_c_531_n N_VGND_c_1721_n 7.3375e-19 $X=4.545 $Y=1.645 $X2=0 $Y2=0
cc_451 N_CLK_M1001_g N_VGND_c_1723_n 0.00207769f $X=4.635 $Y=0.745 $X2=0 $Y2=0
cc_452 N_CLK_M1001_g N_VGND_c_1735_n 0.00936553f $X=4.635 $Y=0.745 $X2=0 $Y2=0
cc_453 CLK N_VGND_c_1735_n 0.00120566f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_454 N_A_1243_116#_c_567_n N_A_972_569#_M1022_g 0.00951227f $X=6.355 $Y=0.79
+ $X2=0 $Y2=0
cc_455 N_A_1243_116#_c_576_n N_A_972_569#_M1022_g 0.00549407f $X=6.377 $Y=1.02
+ $X2=0 $Y2=0
cc_456 N_A_1243_116#_c_577_n N_A_972_569#_M1022_g 0.0042676f $X=6.52 $Y=2.29
+ $X2=0 $Y2=0
cc_457 N_A_1243_116#_c_589_n N_A_972_569#_M1011_g 0.00442926f $X=6.52 $Y=2.415
+ $X2=0 $Y2=0
cc_458 N_A_1243_116#_c_590_n N_A_972_569#_M1011_g 0.0154166f $X=6.56 $Y=2.585
+ $X2=0 $Y2=0
cc_459 N_A_1243_116#_c_577_n N_A_972_569#_M1011_g 0.0170393f $X=6.52 $Y=2.29
+ $X2=0 $Y2=0
cc_460 N_A_1243_116#_c_589_n N_A_972_569#_c_743_n 0.00221357f $X=6.52 $Y=2.415
+ $X2=0 $Y2=0
cc_461 N_A_1243_116#_c_568_n N_A_972_569#_c_743_n 0.00393368f $X=7.19 $Y=0.35
+ $X2=0 $Y2=0
cc_462 N_A_1243_116#_c_577_n N_A_972_569#_c_743_n 0.0205239f $X=6.52 $Y=2.29
+ $X2=0 $Y2=0
cc_463 N_A_1243_116#_c_567_n N_A_972_569#_c_744_n 0.00247818f $X=6.355 $Y=0.79
+ $X2=19.92 $Y2=0
cc_464 N_A_1243_116#_c_568_n N_A_972_569#_c_744_n 0.00473366f $X=7.19 $Y=0.35
+ $X2=19.92 $Y2=0
cc_465 N_A_1243_116#_c_572_n N_A_972_569#_c_744_n 0.00742959f $X=8.05 $Y=0.35
+ $X2=19.92 $Y2=0
cc_466 N_A_1243_116#_c_580_n N_A_972_569#_c_744_n 0.0297463f $X=7.355 $Y=2.29
+ $X2=19.92 $Y2=0
cc_467 N_A_1243_116#_c_581_n N_A_972_569#_c_744_n 0.0011518f $X=8.187 $Y=1.15
+ $X2=19.92 $Y2=0
cc_468 N_A_1243_116#_M1023_g N_A_972_569#_c_744_n 0.0299511f $X=8.095 $Y=0.81
+ $X2=19.92 $Y2=0
cc_469 N_A_1243_116#_M1023_g N_A_972_569#_c_745_n 0.0344742f $X=8.095 $Y=0.81
+ $X2=0 $Y2=0
cc_470 N_A_1243_116#_c_575_n N_A_972_569#_c_746_n 0.00742147f $X=8.325 $Y=1.645
+ $X2=0 $Y2=0
cc_471 N_A_1243_116#_c_592_n N_A_972_569#_c_746_n 0.0204877f $X=7.355 $Y=2.455
+ $X2=0 $Y2=0
cc_472 N_A_1243_116#_c_580_n N_A_972_569#_c_746_n 4.18249e-19 $X=7.355 $Y=2.29
+ $X2=0 $Y2=0
cc_473 N_A_1243_116#_c_583_n N_A_972_569#_c_746_n 0.00628961f $X=12.2 $Y=1.717
+ $X2=0 $Y2=0
cc_474 N_A_1243_116#_c_592_n N_A_972_569#_M1030_g 0.0141933f $X=7.355 $Y=2.455
+ $X2=0 $Y2=0
cc_475 N_A_1243_116#_c_587_n N_A_972_569#_c_762_n 0.00863239f $X=13.185 $Y=2.605
+ $X2=0 $Y2=0
cc_476 N_A_1243_116#_c_588_n N_A_972_569#_c_762_n 0.00127578f $X=12.78 $Y=2.45
+ $X2=0 $Y2=0
cc_477 N_A_1243_116#_c_582_n N_A_972_569#_c_762_n 7.65899e-19 $X=12.365 $Y=1.71
+ $X2=0 $Y2=0
cc_478 N_A_1243_116#_c_621_p N_A_972_569#_c_747_n 0.00117034f $X=7.355 $Y=2.455
+ $X2=0 $Y2=0
cc_479 N_A_1243_116#_c_592_n N_A_972_569#_c_747_n 0.0439072f $X=7.355 $Y=2.455
+ $X2=0 $Y2=0
cc_480 N_A_1243_116#_c_580_n N_A_972_569#_c_747_n 0.0421991f $X=7.355 $Y=2.29
+ $X2=0 $Y2=0
cc_481 N_A_1243_116#_M1041_g N_A_972_569#_M1008_g 0.0131401f $X=12.43 $Y=0.91
+ $X2=0 $Y2=0
cc_482 N_A_1243_116#_c_577_n N_A_972_569#_c_751_n 0.00759532f $X=6.52 $Y=2.29
+ $X2=0 $Y2=0
cc_483 N_A_1243_116#_c_577_n N_A_972_569#_c_818_n 0.0209681f $X=6.52 $Y=2.29
+ $X2=0 $Y2=0
cc_484 N_A_1243_116#_c_576_n N_A_972_569#_c_752_n 0.0046479f $X=6.377 $Y=1.02
+ $X2=0 $Y2=0
cc_485 N_A_1243_116#_c_577_n N_A_972_569#_c_752_n 0.0229141f $X=6.52 $Y=2.29
+ $X2=0 $Y2=0
cc_486 N_A_1243_116#_c_629_p N_A_972_569#_c_821_n 0.00787995f $X=12.365 $Y=1.71
+ $X2=0 $Y2=0
cc_487 N_A_1243_116#_c_582_n N_A_972_569#_c_821_n 6.20123e-19 $X=12.365 $Y=1.71
+ $X2=0 $Y2=0
cc_488 N_A_1243_116#_c_583_n N_A_972_569#_c_821_n 0.00731768f $X=12.2 $Y=1.717
+ $X2=0 $Y2=0
cc_489 N_A_1243_116#_c_588_n N_A_972_569#_c_824_n 0.00144777f $X=12.78 $Y=2.45
+ $X2=0 $Y2=0
cc_490 N_A_1243_116#_c_586_n N_A_972_569#_c_773_n 0.0240419f $X=12.78 $Y=2.295
+ $X2=0 $Y2=0
cc_491 N_A_1243_116#_c_588_n N_A_972_569#_c_773_n 0.00989353f $X=12.78 $Y=2.45
+ $X2=0 $Y2=0
cc_492 N_A_1243_116#_c_629_p N_A_972_569#_c_773_n 0.0105165f $X=12.365 $Y=1.71
+ $X2=0 $Y2=0
cc_493 N_A_1243_116#_c_582_n N_A_972_569#_c_773_n 0.0064933f $X=12.365 $Y=1.71
+ $X2=0 $Y2=0
cc_494 N_A_1243_116#_M1041_g N_A_972_569#_c_774_n 0.00116628f $X=12.43 $Y=0.91
+ $X2=0 $Y2=0
cc_495 N_A_1243_116#_c_586_n N_A_972_569#_c_774_n 0.00136783f $X=12.78 $Y=2.295
+ $X2=0 $Y2=0
cc_496 N_A_1243_116#_c_629_p N_A_972_569#_c_774_n 0.007903f $X=12.365 $Y=1.71
+ $X2=0 $Y2=0
cc_497 N_A_1243_116#_c_582_n N_A_972_569#_c_774_n 0.0024675f $X=12.365 $Y=1.71
+ $X2=0 $Y2=0
cc_498 N_A_1243_116#_M1041_g N_A_972_569#_c_753_n 0.00663239f $X=12.43 $Y=0.91
+ $X2=0 $Y2=0
cc_499 N_A_1243_116#_c_588_n N_A_972_569#_c_753_n 0.0210361f $X=12.78 $Y=2.45
+ $X2=0 $Y2=0
cc_500 N_A_1243_116#_c_629_p N_A_972_569#_c_753_n 7.64902e-19 $X=12.365 $Y=1.71
+ $X2=0 $Y2=0
cc_501 N_A_1243_116#_c_582_n N_A_972_569#_c_753_n 0.0322829f $X=12.365 $Y=1.71
+ $X2=0 $Y2=0
cc_502 N_A_1243_116#_c_592_n N_A_972_569#_c_837_n 3.35508e-19 $X=7.355 $Y=2.455
+ $X2=0 $Y2=0
cc_503 N_A_1243_116#_c_586_n N_A_972_569#_c_779_n 0.0184567f $X=12.78 $Y=2.295
+ $X2=0 $Y2=0
cc_504 N_A_1243_116#_c_588_n N_A_972_569#_c_779_n 0.0110899f $X=12.78 $Y=2.45
+ $X2=0 $Y2=0
cc_505 N_A_1243_116#_c_629_p N_A_972_569#_c_779_n 9.51312e-19 $X=12.365 $Y=1.71
+ $X2=0 $Y2=0
cc_506 N_A_1243_116#_c_582_n N_A_972_569#_c_779_n 0.01799f $X=12.365 $Y=1.71
+ $X2=0 $Y2=0
cc_507 N_A_1243_116#_c_583_n N_A_972_569#_c_779_n 0.0042382f $X=12.2 $Y=1.717
+ $X2=0 $Y2=0
cc_508 N_A_1243_116#_c_651_p N_A_1711_94#_c_954_n 0.00646527f $X=8.187 $Y=1.287
+ $X2=0.24 $Y2=0
cc_509 N_A_1243_116#_c_583_n N_A_1711_94#_c_954_n 0.0713053f $X=12.2 $Y=1.717
+ $X2=0.24 $Y2=0
cc_510 N_A_1243_116#_M1023_g N_A_1711_94#_c_954_n 5.42624e-19 $X=8.095 $Y=0.81
+ $X2=0.24 $Y2=0
cc_511 N_A_1243_116#_c_651_p N_A_1711_94#_c_955_n 0.00195983f $X=8.187 $Y=1.287
+ $X2=0 $Y2=0
cc_512 N_A_1243_116#_c_583_n N_A_1711_94#_c_955_n 0.00723311f $X=12.2 $Y=1.717
+ $X2=0 $Y2=0
cc_513 N_A_1243_116#_c_574_n N_A_1711_94#_c_956_n 0.00185606f $X=8.16 $Y=1.315
+ $X2=0 $Y2=0
cc_514 N_A_1243_116#_c_583_n N_A_1711_94#_c_956_n 0.0301731f $X=12.2 $Y=1.717
+ $X2=0 $Y2=0
cc_515 N_A_1243_116#_c_581_n N_A_1711_94#_c_959_n 0.00153271f $X=8.187 $Y=1.15
+ $X2=0 $Y2=0
cc_516 N_A_1243_116#_M1023_g N_A_1711_94#_c_959_n 0.0711191f $X=8.095 $Y=0.81
+ $X2=0 $Y2=0
cc_517 N_A_1243_116#_c_583_n N_A_1513_120#_c_1005_n 0.00882775f $X=12.2 $Y=1.717
+ $X2=0 $Y2=0
cc_518 N_A_1243_116#_M1041_g N_A_1513_120#_M1024_g 0.0529822f $X=12.43 $Y=0.91
+ $X2=0 $Y2=0
cc_519 N_A_1243_116#_c_629_p N_A_1513_120#_M1024_g 0.00101821f $X=12.365 $Y=1.71
+ $X2=0 $Y2=0
cc_520 N_A_1243_116#_c_583_n N_A_1513_120#_M1024_g 0.0348653f $X=12.2 $Y=1.717
+ $X2=0 $Y2=0
cc_521 N_A_1243_116#_c_582_n N_A_1513_120#_c_1009_n 0.0529822f $X=12.365 $Y=1.71
+ $X2=10.08 $Y2=0
cc_522 N_A_1243_116#_c_583_n N_A_1513_120#_c_1009_n 0.00482482f $X=12.2 $Y=1.717
+ $X2=10.08 $Y2=0
cc_523 N_A_1243_116#_c_651_p N_A_1513_120#_c_1010_n 0.0311855f $X=8.187 $Y=1.287
+ $X2=10.08 $Y2=0.057
cc_524 N_A_1243_116#_c_575_n N_A_1513_120#_c_1010_n 0.0136205f $X=8.325 $Y=1.645
+ $X2=10.08 $Y2=0.057
cc_525 N_A_1243_116#_c_580_n N_A_1513_120#_c_1010_n 0.0354597f $X=7.355 $Y=2.29
+ $X2=10.08 $Y2=0.057
cc_526 N_A_1243_116#_M1023_g N_A_1513_120#_c_1010_n 0.0104444f $X=8.095 $Y=0.81
+ $X2=10.08 $Y2=0.057
cc_527 N_A_1243_116#_c_621_p N_A_1513_120#_c_1014_n 0.0191896f $X=7.355 $Y=2.455
+ $X2=0 $Y2=0
cc_528 N_A_1243_116#_c_592_n N_A_1513_120#_c_1014_n 0.0156988f $X=7.355 $Y=2.455
+ $X2=0 $Y2=0
cc_529 N_A_1243_116#_c_580_n N_A_1513_120#_c_1014_n 0.0100111f $X=7.355 $Y=2.29
+ $X2=0 $Y2=0
cc_530 N_A_1243_116#_c_595_n N_A_1513_120#_c_1014_n 0.0207126f $X=7.47 $Y=2.67
+ $X2=0 $Y2=0
cc_531 N_A_1243_116#_c_575_n N_A_1513_120#_c_1015_n 0.0199042f $X=8.325 $Y=1.645
+ $X2=0 $Y2=0
cc_532 N_A_1243_116#_c_583_n N_A_1513_120#_c_1015_n 0.201936f $X=12.2 $Y=1.717
+ $X2=0 $Y2=0
cc_533 N_A_1243_116#_M1023_g N_A_1513_120#_c_1015_n 4.56806e-19 $X=8.095 $Y=0.81
+ $X2=0 $Y2=0
cc_534 N_A_1243_116#_c_583_n N_A_1513_120#_c_1011_n 0.0332717f $X=12.2 $Y=1.717
+ $X2=0 $Y2=0
cc_535 N_A_1243_116#_c_572_n N_A_1513_120#_c_1012_n 0.0152699f $X=8.05 $Y=0.35
+ $X2=0 $Y2=0
cc_536 N_A_1243_116#_c_580_n N_A_1513_120#_c_1012_n 0.0286495f $X=7.355 $Y=2.29
+ $X2=0 $Y2=0
cc_537 N_A_1243_116#_c_581_n N_A_1513_120#_c_1012_n 0.0311855f $X=8.187 $Y=1.15
+ $X2=0 $Y2=0
cc_538 N_A_1243_116#_M1023_g N_A_1513_120#_c_1012_n 0.00774158f $X=8.095 $Y=0.81
+ $X2=0 $Y2=0
cc_539 N_A_1243_116#_c_580_n N_A_1513_120#_c_1018_n 0.00758407f $X=7.355 $Y=2.29
+ $X2=0 $Y2=0
cc_540 N_A_1243_116#_M1023_g N_A_1513_120#_c_1018_n 6.24248e-19 $X=8.095 $Y=0.81
+ $X2=0 $Y2=0
cc_541 N_A_1243_116#_c_583_n N_A_1513_120#_c_1046_n 0.0244834f $X=12.2 $Y=1.717
+ $X2=0 $Y2=0
cc_542 N_A_1243_116#_c_583_n N_SET_B_c_1110_n 0.0342516f $X=12.2 $Y=1.717
+ $X2=-0.33 $Y2=-0.265
cc_543 N_A_1243_116#_M1041_g N_SET_B_c_1111_n 0.014545f $X=12.43 $Y=0.91 $X2=0
+ $Y2=0
cc_544 N_A_1243_116#_M1041_g N_SET_B_c_1113_n 0.00389575f $X=12.43 $Y=0.91 $X2=0
+ $Y2=0
cc_545 N_A_1243_116#_M1041_g SET_B 0.0474815f $X=12.43 $Y=0.91 $X2=0 $Y2=0
cc_546 N_A_1243_116#_c_583_n SET_B 0.0128343f $X=12.2 $Y=1.717 $X2=0 $Y2=0
cc_547 N_A_1243_116#_M1041_g N_SET_B_c_1119_n 0.00159657f $X=12.43 $Y=0.91 $X2=0
+ $Y2=0
cc_548 N_A_1243_116#_c_583_n N_SET_B_c_1119_n 0.134866f $X=12.2 $Y=1.717 $X2=0
+ $Y2=0
cc_549 N_A_1243_116#_c_587_n N_A_2729_463#_c_1196_n 0.0320532f $X=13.185
+ $Y=2.605 $X2=0 $Y2=0
cc_550 N_A_1243_116#_c_588_n N_A_2729_463#_c_1196_n 0.0320532f $X=12.78 $Y=2.45
+ $X2=0 $Y2=0
cc_551 N_A_1243_116#_c_588_n N_A_2729_463#_M1009_g 6.14537e-19 $X=12.78 $Y=2.45
+ $X2=0 $Y2=0
cc_552 N_A_1243_116#_c_587_n N_A_2501_543#_c_1260_n 0.0118782f $X=13.185
+ $Y=2.605 $X2=0 $Y2=0
cc_553 N_A_1243_116#_c_587_n N_A_2501_543#_c_1263_n 0.0274055f $X=13.185
+ $Y=2.605 $X2=0 $Y2=0
cc_554 N_A_1243_116#_c_588_n N_A_2501_543#_c_1263_n 0.0147283f $X=12.78 $Y=2.45
+ $X2=0 $Y2=0
cc_555 N_A_1243_116#_c_588_n N_A_2501_543#_c_1264_n 0.00898293f $X=12.78 $Y=2.45
+ $X2=0 $Y2=0
cc_556 N_A_1243_116#_c_586_n N_A_2501_543#_c_1265_n 4.97229e-19 $X=12.78
+ $Y=2.295 $X2=0 $Y2=0
cc_557 N_A_1243_116#_c_588_n N_A_2501_543#_c_1265_n 0.00498254f $X=12.78 $Y=2.45
+ $X2=0 $Y2=0
cc_558 N_A_1243_116#_M1041_g N_A_2501_543#_c_1249_n 0.0175525f $X=12.43 $Y=0.91
+ $X2=0 $Y2=0
cc_559 N_A_1243_116#_c_582_n N_A_2501_543#_c_1249_n 0.00966982f $X=12.365
+ $Y=1.71 $X2=0 $Y2=0
cc_560 N_A_1243_116#_c_587_n N_VPWR_c_1434_n 0.00626054f $X=13.185 $Y=2.605
+ $X2=0 $Y2=0
cc_561 N_A_1243_116#_c_587_n N_VPWR_c_1443_n 0.0156697f $X=13.185 $Y=2.605 $X2=0
+ $Y2=0
cc_562 N_A_1243_116#_c_590_n N_VPWR_c_1443_n 0.00179277f $X=6.56 $Y=2.585 $X2=0
+ $Y2=0
cc_563 N_A_1243_116#_c_595_n N_VPWR_c_1443_n 0.0154875f $X=7.47 $Y=2.67 $X2=0
+ $Y2=0
cc_564 N_A_1243_116#_c_577_n N_A_485_569#_c_1554_n 0.0123662f $X=6.52 $Y=2.29
+ $X2=0 $Y2=0
cc_565 N_A_1243_116#_c_577_n N_A_485_569#_c_1556_n 0.0658156f $X=6.52 $Y=2.29
+ $X2=0 $Y2=0
cc_566 N_A_1243_116#_c_590_n N_A_485_569#_c_1557_n 0.0180295f $X=6.56 $Y=2.585
+ $X2=0 $Y2=0
cc_567 N_A_1243_116#_c_567_n N_A_485_569#_c_1539_n 0.0164405f $X=6.355 $Y=0.79
+ $X2=0 $Y2=0
cc_568 N_A_1243_116#_c_568_n N_A_485_569#_c_1539_n 0.0166151f $X=7.19 $Y=0.35
+ $X2=0 $Y2=0
cc_569 N_A_1243_116#_c_580_n N_A_485_569#_c_1539_n 0.0592845f $X=7.355 $Y=2.29
+ $X2=0 $Y2=0
cc_570 N_A_1243_116#_c_590_n N_A_485_569#_c_1563_n 0.0330779f $X=6.56 $Y=2.585
+ $X2=0 $Y2=0
cc_571 N_A_1243_116#_c_621_p N_A_485_569#_c_1563_n 0.00868214f $X=7.355 $Y=2.455
+ $X2=0 $Y2=0
cc_572 N_A_1243_116#_c_592_n N_A_485_569#_c_1563_n 0.00323554f $X=7.355 $Y=2.455
+ $X2=0 $Y2=0
cc_573 N_A_1243_116#_c_595_n N_A_485_569#_c_1563_n 0.00727565f $X=7.47 $Y=2.67
+ $X2=0 $Y2=0
cc_574 N_A_1243_116#_c_595_n N_A_485_569#_c_1564_n 0.0148631f $X=7.47 $Y=2.67
+ $X2=0 $Y2=0
cc_575 N_A_1243_116#_c_576_n N_A_485_569#_c_1542_n 0.0164405f $X=6.377 $Y=1.02
+ $X2=0 $Y2=0
cc_576 N_A_1243_116#_c_621_p N_A_485_569#_c_1542_n 0.0592845f $X=7.355 $Y=2.455
+ $X2=0 $Y2=0
cc_577 N_A_1243_116#_c_589_n N_A_485_569#_c_1543_n 0.0330779f $X=6.52 $Y=2.415
+ $X2=0 $Y2=0
cc_578 N_A_1243_116#_c_577_n N_A_485_569#_c_1543_n 0.0623722f $X=6.52 $Y=2.29
+ $X2=0 $Y2=0
cc_579 N_A_1243_116#_c_592_n N_A_485_569#_c_1543_n 0.0119859f $X=7.355 $Y=2.455
+ $X2=0 $Y2=0
cc_580 N_A_1243_116#_c_595_n N_A_485_569#_c_1543_n 0.00247963f $X=7.47 $Y=2.67
+ $X2=0 $Y2=0
cc_581 N_A_1243_116#_c_567_n N_VGND_c_1723_n 0.0335251f $X=6.355 $Y=0.79 $X2=0
+ $Y2=0
cc_582 N_A_1243_116#_c_570_n N_VGND_c_1723_n 0.00384269f $X=6.565 $Y=0.35 $X2=0
+ $Y2=0
cc_583 N_A_1243_116#_c_572_n N_VGND_c_1725_n 0.00464341f $X=8.05 $Y=0.35 $X2=0
+ $Y2=0
cc_584 N_A_1243_116#_c_581_n N_VGND_c_1725_n 0.0359171f $X=8.187 $Y=1.15 $X2=0
+ $Y2=0
cc_585 N_A_1243_116#_c_583_n N_VGND_c_1725_n 0.0138504f $X=12.2 $Y=1.717 $X2=0
+ $Y2=0
cc_586 N_A_1243_116#_M1023_g N_VGND_c_1725_n 0.0037704f $X=8.095 $Y=0.81 $X2=0
+ $Y2=0
cc_587 N_A_1243_116#_M1041_g N_VGND_c_1727_n 0.00227306f $X=12.43 $Y=0.91 $X2=0
+ $Y2=0
cc_588 N_A_1243_116#_M1041_g N_VGND_c_1735_n 0.0168464f $X=12.43 $Y=0.91 $X2=0
+ $Y2=0
cc_589 N_A_1243_116#_c_567_n N_VGND_c_1735_n 0.0284984f $X=6.355 $Y=0.79 $X2=0
+ $Y2=0
cc_590 N_A_1243_116#_c_568_n N_VGND_c_1735_n 0.0259067f $X=7.19 $Y=0.35 $X2=0
+ $Y2=0
cc_591 N_A_1243_116#_c_570_n N_VGND_c_1735_n 0.0122262f $X=6.565 $Y=0.35 $X2=0
+ $Y2=0
cc_592 N_A_1243_116#_c_572_n N_VGND_c_1735_n 0.0350673f $X=8.05 $Y=0.35 $X2=0
+ $Y2=0
cc_593 N_A_1243_116#_c_651_p N_VGND_c_1735_n 0.00338714f $X=8.187 $Y=1.287 $X2=0
+ $Y2=0
cc_594 N_A_1243_116#_c_578_n N_VGND_c_1735_n 0.00355762f $X=7.275 $Y=0.35 $X2=0
+ $Y2=0
cc_595 N_A_1243_116#_c_580_n N_VGND_c_1735_n 0.0228228f $X=7.355 $Y=2.29 $X2=0
+ $Y2=0
cc_596 N_A_1243_116#_c_581_n N_VGND_c_1735_n 0.0205068f $X=8.187 $Y=1.15 $X2=0
+ $Y2=0
cc_597 N_A_1243_116#_M1023_g N_VGND_c_1735_n 0.016818f $X=8.095 $Y=0.81 $X2=0
+ $Y2=0
cc_598 N_A_972_569#_c_769_n N_A_1711_94#_M1013_d 0.00180746f $X=10.605 $Y=3.255
+ $X2=0 $Y2=0
cc_599 N_A_972_569#_c_746_n N_A_1711_94#_c_960_n 5.80236e-19 $X=8.3 $Y=2.65
+ $X2=0 $Y2=0
cc_600 N_A_972_569#_c_768_n N_A_1711_94#_c_960_n 0.0691251f $X=9.745 $Y=2.695
+ $X2=0 $Y2=0
cc_601 N_A_972_569#_c_837_n N_A_1711_94#_c_960_n 0.00579499f $X=8.365 $Y=2.455
+ $X2=0 $Y2=0
cc_602 N_A_972_569#_c_746_n N_A_1711_94#_c_956_n 0.110794f $X=8.3 $Y=2.65 $X2=0
+ $Y2=0
cc_603 N_A_972_569#_c_768_n N_A_1711_94#_c_956_n 0.0276729f $X=9.745 $Y=2.695
+ $X2=0 $Y2=0
cc_604 N_A_972_569#_c_849_p N_A_1711_94#_c_956_n 6.90313e-19 $X=9.83 $Y=3.17
+ $X2=0 $Y2=0
cc_605 N_A_972_569#_c_837_n N_A_1711_94#_c_956_n 0.00194047f $X=8.365 $Y=2.455
+ $X2=0 $Y2=0
cc_606 N_A_972_569#_c_768_n N_A_1711_94#_c_980_n 0.0129587f $X=9.745 $Y=2.695
+ $X2=0 $Y2=0
cc_607 N_A_972_569#_c_849_p N_A_1711_94#_c_980_n 0.0142924f $X=9.83 $Y=3.17
+ $X2=0 $Y2=0
cc_608 N_A_972_569#_c_769_n N_A_1711_94#_c_980_n 0.0155034f $X=10.605 $Y=3.255
+ $X2=0 $Y2=0
cc_609 N_A_972_569#_c_744_n N_A_1513_120#_c_1010_n 0.0101706f $X=7.315 $Y=1.13
+ $X2=10.08 $Y2=0.057
cc_610 N_A_972_569#_c_745_n N_A_1513_120#_c_1010_n 0.0188034f $X=8.01 $Y=1.885
+ $X2=10.08 $Y2=0.057
cc_611 N_A_972_569#_c_746_n N_A_1513_120#_c_1014_n 0.0134673f $X=8.3 $Y=2.65
+ $X2=0 $Y2=0
cc_612 N_A_972_569#_M1030_g N_A_1513_120#_c_1014_n 0.0019534f $X=8.3 $Y=2.99
+ $X2=0 $Y2=0
cc_613 N_A_972_569#_c_837_n N_A_1513_120#_c_1014_n 0.0333303f $X=8.365 $Y=2.455
+ $X2=0 $Y2=0
cc_614 N_A_972_569#_c_745_n N_A_1513_120#_c_1015_n 5.66483e-19 $X=8.01 $Y=1.885
+ $X2=0 $Y2=0
cc_615 N_A_972_569#_c_746_n N_A_1513_120#_c_1015_n 0.0315224f $X=8.3 $Y=2.65
+ $X2=0 $Y2=0
cc_616 N_A_972_569#_c_768_n N_A_1513_120#_c_1015_n 0.011736f $X=9.745 $Y=2.695
+ $X2=0 $Y2=0
cc_617 N_A_972_569#_c_837_n N_A_1513_120#_c_1015_n 0.0205132f $X=8.365 $Y=2.455
+ $X2=0 $Y2=0
cc_618 N_A_972_569#_c_768_n N_A_1513_120#_c_1011_n 0.0190377f $X=9.745 $Y=2.695
+ $X2=0 $Y2=0
cc_619 N_A_972_569#_c_849_p N_A_1513_120#_c_1011_n 0.0164678f $X=9.83 $Y=3.17
+ $X2=0 $Y2=0
cc_620 N_A_972_569#_c_769_n N_A_1513_120#_c_1011_n 0.0160918f $X=10.605 $Y=3.255
+ $X2=0 $Y2=0
cc_621 N_A_972_569#_c_771_n N_A_1513_120#_c_1011_n 0.00626001f $X=9.915 $Y=3.255
+ $X2=0 $Y2=0
cc_622 N_A_972_569#_c_777_n N_A_1513_120#_c_1011_n 6.40009e-19 $X=10.69 $Y=3.085
+ $X2=0 $Y2=0
cc_623 N_A_972_569#_c_744_n N_A_1513_120#_c_1012_n 0.00906789f $X=7.315 $Y=1.13
+ $X2=0 $Y2=0
cc_624 N_A_972_569#_c_745_n N_A_1513_120#_c_1012_n 0.00343421f $X=8.01 $Y=1.885
+ $X2=0 $Y2=0
cc_625 N_A_972_569#_c_745_n N_A_1513_120#_c_1018_n 0.0157779f $X=8.01 $Y=1.885
+ $X2=0 $Y2=0
cc_626 N_A_972_569#_c_871_p N_A_1513_120#_c_1046_n 0.01138f $X=12.025 $Y=3.085
+ $X2=0 $Y2=0
cc_627 N_A_972_569#_c_821_n N_A_1513_120#_c_1046_n 0.00708731f $X=12.18 $Y=2.295
+ $X2=0 $Y2=0
cc_628 N_A_972_569#_c_824_n N_A_1513_120#_c_1046_n 0.0101484f $X=12.18 $Y=3
+ $X2=0 $Y2=0
cc_629 N_A_972_569#_c_779_n N_A_1513_120#_c_1046_n 0.0013755f $X=12.19 $Y=2.29
+ $X2=0 $Y2=0
cc_630 N_A_972_569#_c_871_p N_A_1513_120#_c_1019_n 0.0341337f $X=12.025 $Y=3.085
+ $X2=0 $Y2=0
cc_631 N_A_972_569#_c_821_n N_A_1513_120#_c_1019_n 6.79994e-19 $X=12.18 $Y=2.295
+ $X2=0 $Y2=0
cc_632 N_A_972_569#_c_824_n N_A_1513_120#_c_1019_n 0.00417591f $X=12.18 $Y=3
+ $X2=0 $Y2=0
cc_633 N_A_972_569#_c_777_n N_A_1513_120#_c_1019_n 9.01456e-19 $X=10.69 $Y=3.085
+ $X2=0 $Y2=0
cc_634 N_A_972_569#_c_779_n N_A_1513_120#_c_1019_n 0.121345f $X=12.19 $Y=2.29
+ $X2=0 $Y2=0
cc_635 N_A_972_569#_c_849_p N_SET_B_M1018_g 5.99284e-19 $X=9.83 $Y=3.17 $X2=0
+ $Y2=0
cc_636 N_A_972_569#_c_769_n N_SET_B_M1018_g 0.0171342f $X=10.605 $Y=3.255 $X2=0
+ $Y2=0
cc_637 N_A_972_569#_c_871_p N_SET_B_M1018_g 0.0130244f $X=12.025 $Y=3.085 $X2=0
+ $Y2=0
cc_638 N_A_972_569#_c_777_n N_SET_B_M1018_g 0.0220842f $X=10.69 $Y=3.085 $X2=0
+ $Y2=0
cc_639 N_A_972_569#_M1008_g N_SET_B_c_1111_n 0.00231099f $X=13.325 $Y=1.075
+ $X2=0 $Y2=0
cc_640 N_A_972_569#_M1008_g N_SET_B_c_1115_n 2.81388e-19 $X=13.325 $Y=1.075
+ $X2=0 $Y2=0
cc_641 N_A_972_569#_M1008_g N_A_2729_463#_M1009_g 0.0839752f $X=13.325 $Y=1.075
+ $X2=0 $Y2=0
cc_642 N_A_972_569#_c_774_n N_A_2729_463#_M1009_g 2.80576e-19 $X=13.285 $Y=1.58
+ $X2=0 $Y2=0
cc_643 N_A_972_569#_c_762_n N_A_2501_543#_c_1260_n 0.00256916f $X=12.255
+ $Y=2.835 $X2=0 $Y2=0
cc_644 N_A_972_569#_c_824_n N_A_2501_543#_c_1260_n 0.0114757f $X=12.18 $Y=3
+ $X2=0 $Y2=0
cc_645 N_A_972_569#_c_773_n N_A_2501_543#_c_1263_n 0.0322925f $X=13.165 $Y=2.21
+ $X2=0 $Y2=0
cc_646 N_A_972_569#_c_753_n N_A_2501_543#_c_1263_n 0.00469089f $X=13.285 $Y=1.58
+ $X2=0 $Y2=0
cc_647 N_A_972_569#_c_762_n N_A_2501_543#_c_1264_n 0.00137633f $X=12.255
+ $Y=2.835 $X2=0 $Y2=0
cc_648 N_A_972_569#_c_824_n N_A_2501_543#_c_1264_n 0.0136361f $X=12.18 $Y=3
+ $X2=0 $Y2=0
cc_649 N_A_972_569#_c_773_n N_A_2501_543#_c_1264_n 0.0211749f $X=13.165 $Y=2.21
+ $X2=0 $Y2=0
cc_650 N_A_972_569#_c_779_n N_A_2501_543#_c_1264_n 5.33628e-19 $X=12.19 $Y=2.29
+ $X2=0 $Y2=0
cc_651 N_A_972_569#_M1008_g N_A_2501_543#_c_1246_n 0.0298896f $X=13.325 $Y=1.075
+ $X2=0 $Y2=0
cc_652 N_A_972_569#_c_774_n N_A_2501_543#_c_1246_n 0.00608615f $X=13.285 $Y=1.58
+ $X2=0 $Y2=0
cc_653 N_A_972_569#_M1008_g N_A_2501_543#_c_1247_n 0.00906909f $X=13.325
+ $Y=1.075 $X2=0 $Y2=0
cc_654 N_A_972_569#_c_774_n N_A_2501_543#_c_1247_n 0.0287393f $X=13.285 $Y=1.58
+ $X2=0 $Y2=0
cc_655 N_A_972_569#_c_773_n N_A_2501_543#_c_1265_n 0.0137873f $X=13.165 $Y=2.21
+ $X2=0 $Y2=0
cc_656 N_A_972_569#_c_774_n N_A_2501_543#_c_1265_n 0.00922058f $X=13.285 $Y=1.58
+ $X2=0 $Y2=0
cc_657 N_A_972_569#_c_753_n N_A_2501_543#_c_1265_n 7.01845e-19 $X=13.285 $Y=1.58
+ $X2=0 $Y2=0
cc_658 N_A_972_569#_M1008_g N_A_2501_543#_c_1249_n 0.0085184f $X=13.325 $Y=1.075
+ $X2=0 $Y2=0
cc_659 N_A_972_569#_c_774_n N_A_2501_543#_c_1250_n 0.0134383f $X=13.285 $Y=1.58
+ $X2=0 $Y2=0
cc_660 N_A_972_569#_c_753_n N_A_2501_543#_c_1250_n 0.00154707f $X=13.285 $Y=1.58
+ $X2=0 $Y2=0
cc_661 N_A_972_569#_c_871_p N_VPWR_M1018_d 0.0139121f $X=12.025 $Y=3.085
+ $X2=-0.33 $Y2=-0.265
cc_662 N_A_972_569#_M1011_g N_VPWR_c_1425_n 0.00755044f $X=6.17 $Y=2.815 $X2=0
+ $Y2=0
cc_663 N_A_972_569#_M1030_g N_VPWR_c_1428_n 0.00717777f $X=8.3 $Y=2.99 $X2=0
+ $Y2=0
cc_664 N_A_972_569#_c_768_n N_VPWR_c_1428_n 0.0669162f $X=9.745 $Y=2.695 $X2=0
+ $Y2=0
cc_665 N_A_972_569#_c_771_n N_VPWR_c_1428_n 0.0131067f $X=9.915 $Y=3.255 $X2=0
+ $Y2=0
cc_666 N_A_972_569#_c_762_n N_VPWR_c_1431_n 0.00454985f $X=12.255 $Y=2.835 $X2=0
+ $Y2=0
cc_667 N_A_972_569#_c_871_p N_VPWR_c_1431_n 0.0551186f $X=12.025 $Y=3.085 $X2=0
+ $Y2=0
cc_668 N_A_972_569#_M1011_g N_VPWR_c_1443_n 0.0040826f $X=6.17 $Y=2.815 $X2=0
+ $Y2=0
cc_669 N_A_972_569#_M1030_g N_VPWR_c_1443_n 0.0162837f $X=8.3 $Y=2.99 $X2=0
+ $Y2=0
cc_670 N_A_972_569#_c_762_n N_VPWR_c_1443_n 0.0227462f $X=12.255 $Y=2.835 $X2=0
+ $Y2=0
cc_671 N_A_972_569#_c_766_n N_VPWR_c_1443_n 0.0227753f $X=5 $Y=2.97 $X2=0 $Y2=0
cc_672 N_A_972_569#_c_769_n N_VPWR_c_1443_n 0.0269931f $X=10.605 $Y=3.255 $X2=0
+ $Y2=0
cc_673 N_A_972_569#_c_771_n N_VPWR_c_1443_n 0.00720935f $X=9.915 $Y=3.255 $X2=0
+ $Y2=0
cc_674 N_A_972_569#_c_871_p N_VPWR_c_1443_n 0.0317371f $X=12.025 $Y=3.085 $X2=0
+ $Y2=0
cc_675 N_A_972_569#_c_777_n N_VPWR_c_1443_n 0.00683654f $X=10.69 $Y=3.085 $X2=0
+ $Y2=0
cc_676 N_A_972_569#_c_754_n N_A_485_569#_c_1546_n 0.00939604f $X=5 $Y=2.805
+ $X2=10.08 $Y2=0
cc_677 N_A_972_569#_c_766_n N_A_485_569#_c_1606_n 0.0442312f $X=5 $Y=2.97 $X2=0
+ $Y2=0
cc_678 N_A_972_569#_c_754_n N_A_485_569#_c_1606_n 0.00891586f $X=5 $Y=2.805
+ $X2=0 $Y2=0
cc_679 N_A_972_569#_c_766_n N_A_485_569#_c_1547_n 0.0209757f $X=5 $Y=2.97 $X2=0
+ $Y2=0
cc_680 N_A_972_569#_M1011_g N_A_485_569#_c_1553_n 0.00518663f $X=6.17 $Y=2.815
+ $X2=0 $Y2=0
cc_681 N_A_972_569#_c_754_n N_A_485_569#_c_1553_n 0.0925296f $X=5 $Y=2.805 $X2=0
+ $Y2=0
cc_682 N_A_972_569#_M1011_g N_A_485_569#_c_1554_n 0.0264158f $X=6.17 $Y=2.815
+ $X2=0 $Y2=0
cc_683 N_A_972_569#_c_751_n N_A_485_569#_c_1554_n 0.0405691f $X=5.735 $Y=1.785
+ $X2=0 $Y2=0
cc_684 N_A_972_569#_c_752_n N_A_485_569#_c_1554_n 0.00548941f $X=5.9 $Y=1.365
+ $X2=0 $Y2=0
cc_685 N_A_972_569#_c_751_n N_A_485_569#_c_1555_n 0.0137879f $X=5.735 $Y=1.785
+ $X2=0 $Y2=0
cc_686 N_A_972_569#_c_754_n N_A_485_569#_c_1555_n 0.0140562f $X=5 $Y=2.805 $X2=0
+ $Y2=0
cc_687 N_A_972_569#_M1011_g N_A_485_569#_c_1556_n 0.0479987f $X=6.17 $Y=2.815
+ $X2=0 $Y2=0
cc_688 N_A_972_569#_M1011_g N_A_485_569#_c_1557_n 0.0090724f $X=6.17 $Y=2.815
+ $X2=0 $Y2=0
cc_689 N_A_972_569#_M1022_g N_A_485_569#_c_1539_n 6.22112e-19 $X=5.965 $Y=0.79
+ $X2=0 $Y2=0
cc_690 N_A_972_569#_c_744_n N_A_485_569#_c_1539_n 0.00365685f $X=7.315 $Y=1.13
+ $X2=0 $Y2=0
cc_691 N_A_972_569#_M1011_g N_A_485_569#_c_1563_n 0.00232834f $X=6.17 $Y=2.815
+ $X2=0 $Y2=0
cc_692 N_A_972_569#_c_747_n N_A_485_569#_c_1563_n 0.00304434f $X=7.315 $Y=1.38
+ $X2=0 $Y2=0
cc_693 N_A_972_569#_M1011_g N_A_485_569#_c_1564_n 0.00247913f $X=6.17 $Y=2.815
+ $X2=0 $Y2=0
cc_694 N_A_972_569#_c_743_n N_A_485_569#_c_1542_n 0.0038708f $X=7.065 $Y=1.38
+ $X2=0 $Y2=0
cc_695 N_A_972_569#_c_743_n N_A_485_569#_c_1543_n 0.0301945f $X=7.065 $Y=1.38
+ $X2=0 $Y2=0
cc_696 N_A_972_569#_c_747_n N_A_485_569#_c_1543_n 0.00631092f $X=7.315 $Y=1.38
+ $X2=0 $Y2=0
cc_697 N_A_972_569#_c_752_n N_A_485_569#_c_1543_n 0.00232834f $X=5.9 $Y=1.365
+ $X2=0 $Y2=0
cc_698 N_A_972_569#_c_871_p A_2359_543# 0.00482642f $X=12.025 $Y=3.085 $X2=0
+ $Y2=0
cc_699 N_A_972_569#_c_749_n N_VGND_c_1721_n 0.0218749f $X=5.025 $Y=0.745 $X2=0
+ $Y2=0
cc_700 N_A_972_569#_M1022_g N_VGND_c_1723_n 0.0335463f $X=5.965 $Y=0.79 $X2=0
+ $Y2=0
cc_701 N_A_972_569#_c_749_n N_VGND_c_1723_n 0.0399118f $X=5.025 $Y=0.745 $X2=0
+ $Y2=0
cc_702 N_A_972_569#_c_818_n N_VGND_c_1723_n 0.0173987f $X=5.9 $Y=1.365 $X2=0
+ $Y2=0
cc_703 N_A_972_569#_M1001_d N_VGND_c_1735_n 0.00221032f $X=4.885 $Y=0.535 $X2=0
+ $Y2=0
cc_704 N_A_972_569#_M1022_g N_VGND_c_1735_n 0.0102145f $X=5.965 $Y=0.79 $X2=0
+ $Y2=0
cc_705 N_A_972_569#_c_744_n N_VGND_c_1735_n 0.0217693f $X=7.315 $Y=1.13 $X2=0
+ $Y2=0
cc_706 N_A_972_569#_c_749_n N_VGND_c_1735_n 0.0236764f $X=5.025 $Y=0.745 $X2=0
+ $Y2=0
cc_707 N_A_972_569#_c_818_n N_VGND_c_1735_n 0.00408083f $X=5.9 $Y=1.365 $X2=0
+ $Y2=0
cc_708 N_A_972_569#_c_752_n N_VGND_c_1735_n 0.00483051f $X=5.9 $Y=1.365 $X2=0
+ $Y2=0
cc_709 N_A_1711_94#_c_954_n N_A_1513_120#_c_1005_n 0.0192419f $X=9.58 $Y=1.26
+ $X2=0 $Y2=0
cc_710 N_A_1711_94#_c_955_n N_A_1513_120#_c_1005_n 0.0395435f $X=9.075 $Y=1.295
+ $X2=0 $Y2=0
cc_711 N_A_1711_94#_c_957_n N_A_1513_120#_c_1005_n 0.0272023f $X=9.745 $Y=0.745
+ $X2=0 $Y2=0
cc_712 N_A_1711_94#_c_959_n N_A_1513_120#_c_1005_n 0.00111541f $X=8.907 $Y=1.13
+ $X2=0 $Y2=0
cc_713 N_A_1711_94#_c_960_n N_A_1513_120#_c_1015_n 0.105766f $X=10.095 $Y=2.345
+ $X2=0 $Y2=0
cc_714 N_A_1711_94#_c_956_n N_A_1513_120#_c_1015_n 0.0279376f $X=9.075 $Y=2.345
+ $X2=0 $Y2=0
cc_715 N_A_1711_94#_c_960_n N_A_1513_120#_c_1011_n 0.0314781f $X=10.095 $Y=2.345
+ $X2=0 $Y2=0
cc_716 N_A_1711_94#_c_956_n N_A_1513_120#_c_1011_n 0.0395435f $X=9.075 $Y=2.345
+ $X2=0 $Y2=0
cc_717 N_A_1711_94#_c_980_n N_A_1513_120#_c_1011_n 0.0192173f $X=10.26 $Y=2.905
+ $X2=0 $Y2=0
cc_718 N_A_1711_94#_c_960_n N_SET_B_M1018_g 0.0110581f $X=10.095 $Y=2.345 $X2=0
+ $Y2=0
cc_719 N_A_1711_94#_c_980_n N_SET_B_M1018_g 0.0307595f $X=10.26 $Y=2.905 $X2=0
+ $Y2=0
cc_720 N_A_1711_94#_c_954_n N_SET_B_M1038_g 2.83782e-19 $X=9.58 $Y=1.26 $X2=0
+ $Y2=0
cc_721 N_A_1711_94#_c_957_n N_SET_B_M1038_g 7.35212e-19 $X=9.745 $Y=0.745 $X2=0
+ $Y2=0
cc_722 N_A_1711_94#_c_954_n N_SET_B_c_1119_n 0.00911601f $X=9.58 $Y=1.26 $X2=0
+ $Y2=0
cc_723 N_A_1711_94#_c_956_n N_VPWR_c_1428_n 0.0390539f $X=9.075 $Y=2.345 $X2=0
+ $Y2=0
cc_724 N_A_1711_94#_c_954_n N_VGND_c_1725_n 0.0307349f $X=9.58 $Y=1.26 $X2=0
+ $Y2=0
cc_725 N_A_1711_94#_c_955_n N_VGND_c_1725_n 0.00541478f $X=9.075 $Y=1.295 $X2=0
+ $Y2=0
cc_726 N_A_1711_94#_c_957_n N_VGND_c_1725_n 0.030862f $X=9.745 $Y=0.745 $X2=0
+ $Y2=0
cc_727 N_A_1711_94#_c_959_n N_VGND_c_1725_n 0.0484313f $X=8.907 $Y=1.13 $X2=0
+ $Y2=0
cc_728 N_A_1711_94#_c_957_n N_VGND_c_1727_n 0.00748247f $X=9.745 $Y=0.745 $X2=0
+ $Y2=0
cc_729 N_A_1711_94#_c_954_n N_VGND_c_1735_n 0.00980819f $X=9.58 $Y=1.26 $X2=0
+ $Y2=0
cc_730 N_A_1711_94#_c_957_n N_VGND_c_1735_n 0.0247997f $X=9.745 $Y=0.745 $X2=0
+ $Y2=0
cc_731 N_A_1513_120#_c_1046_n N_SET_B_M1018_g 0.00258367f $X=11.48 $Y=2.05 $X2=0
+ $Y2=0
cc_732 N_A_1513_120#_c_1019_n N_SET_B_M1018_g 0.0456328f $X=11.48 $Y=2.05 $X2=0
+ $Y2=0
cc_733 N_A_1513_120#_c_1005_n N_SET_B_c_1110_n 0.0358536f $X=10.135 $Y=1.065
+ $X2=-0.33 $Y2=-0.265
cc_734 N_A_1513_120#_M1024_g N_SET_B_c_1110_n 0.00853893f $X=11.72 $Y=0.91
+ $X2=-0.33 $Y2=-0.265
cc_735 N_A_1513_120#_c_1009_n N_SET_B_c_1110_n 0.0203277f $X=11.632 $Y=1.895
+ $X2=-0.33 $Y2=-0.265
cc_736 N_A_1513_120#_c_1015_n N_SET_B_c_1110_n 0.0523892f $X=11.315 $Y=1.995
+ $X2=-0.33 $Y2=-0.265
cc_737 N_A_1513_120#_c_1011_n N_SET_B_c_1110_n 0.0744154f $X=9.935 $Y=1.995
+ $X2=-0.33 $Y2=-0.265
cc_738 N_A_1513_120#_c_1046_n N_SET_B_c_1110_n 5.42421e-19 $X=11.48 $Y=2.05
+ $X2=-0.33 $Y2=-0.265
cc_739 N_A_1513_120#_M1024_g N_SET_B_c_1113_n 3.52271e-19 $X=11.72 $Y=0.91 $X2=0
+ $Y2=0
cc_740 N_A_1513_120#_M1024_g SET_B 0.00632123f $X=11.72 $Y=0.91 $X2=0 $Y2=0
cc_741 N_A_1513_120#_c_1005_n N_SET_B_M1038_g 0.0358536f $X=10.135 $Y=1.065
+ $X2=0 $Y2=0
cc_742 N_A_1513_120#_M1024_g N_SET_B_M1038_g 0.0382739f $X=11.72 $Y=0.91 $X2=0
+ $Y2=0
cc_743 N_A_1513_120#_c_1005_n N_SET_B_c_1119_n 0.0132437f $X=10.135 $Y=1.065
+ $X2=0 $Y2=0
cc_744 N_A_1513_120#_M1024_g N_SET_B_c_1119_n 0.0306909f $X=11.72 $Y=0.91 $X2=0
+ $Y2=0
cc_745 N_A_1513_120#_c_1014_n N_VPWR_c_1428_n 0.00540781f $X=7.91 $Y=2.99 $X2=0
+ $Y2=0
cc_746 N_A_1513_120#_c_1011_n N_VPWR_c_1428_n 0.00307109f $X=9.935 $Y=1.995
+ $X2=0 $Y2=0
cc_747 N_A_1513_120#_c_1019_n N_VPWR_c_1431_n 0.0314063f $X=11.48 $Y=2.05 $X2=0
+ $Y2=0
cc_748 N_A_1513_120#_c_1014_n N_VPWR_c_1443_n 0.0159378f $X=7.91 $Y=2.99 $X2=0
+ $Y2=0
cc_749 N_A_1513_120#_c_1011_n N_VPWR_c_1443_n 0.00408888f $X=9.935 $Y=1.995
+ $X2=0 $Y2=0
cc_750 N_A_1513_120#_c_1019_n N_VPWR_c_1443_n 0.00250239f $X=11.48 $Y=2.05 $X2=0
+ $Y2=0
cc_751 N_A_1513_120#_c_1014_n N_A_485_569#_c_1563_n 0.0189282f $X=7.91 $Y=2.99
+ $X2=0 $Y2=0
cc_752 N_A_1513_120#_c_1005_n N_VGND_c_1725_n 0.00279295f $X=10.135 $Y=1.065
+ $X2=0 $Y2=0
cc_753 N_A_1513_120#_c_1005_n N_VGND_c_1727_n 0.00490519f $X=10.135 $Y=1.065
+ $X2=0 $Y2=0
cc_754 N_A_1513_120#_M1024_g N_VGND_c_1727_n 0.0203225f $X=11.72 $Y=0.91 $X2=0
+ $Y2=0
cc_755 N_A_1513_120#_M1007_d N_VGND_c_1735_n 0.00217792f $X=7.565 $Y=0.6 $X2=0
+ $Y2=0
cc_756 N_A_1513_120#_c_1005_n N_VGND_c_1735_n 0.0281424f $X=10.135 $Y=1.065
+ $X2=0 $Y2=0
cc_757 N_A_1513_120#_M1024_g N_VGND_c_1735_n 0.0174135f $X=11.72 $Y=0.91 $X2=0
+ $Y2=0
cc_758 N_A_1513_120#_c_1012_n N_VGND_c_1735_n 0.0119593f $X=7.705 $Y=0.81 $X2=0
+ $Y2=0
cc_759 N_SET_B_M1010_g N_A_2729_463#_c_1196_n 0.0179898f $X=14.745 $Y=1.075
+ $X2=0 $Y2=0
cc_760 N_SET_B_M1010_g N_A_2729_463#_c_1197_n 0.0329547f $X=14.745 $Y=1.075
+ $X2=0 $Y2=0
cc_761 N_SET_B_c_1111_n N_A_2729_463#_M1009_g 0.00684422f $X=14 $Y=0.35 $X2=0
+ $Y2=0
cc_762 N_SET_B_c_1115_n N_A_2729_463#_M1009_g 0.0290723f $X=14.085 $Y=1.425
+ $X2=0 $Y2=0
cc_763 N_SET_B_c_1160_p N_A_2729_463#_M1009_g 0.00857737f $X=14.17 $Y=1.535
+ $X2=0 $Y2=0
cc_764 N_SET_B_c_1116_n N_A_2729_463#_M1009_g 0.01115f $X=14.68 $Y=1.56 $X2=0
+ $Y2=0
cc_765 N_SET_B_M1010_g N_A_2729_463#_M1009_g 0.130538f $X=14.745 $Y=1.075 $X2=0
+ $Y2=0
cc_766 N_SET_B_c_1116_n N_A_2501_543#_c_1244_n 6.99872e-19 $X=14.68 $Y=1.56
+ $X2=0 $Y2=0
cc_767 N_SET_B_M1010_g N_A_2501_543#_c_1244_n 0.0502318f $X=14.745 $Y=1.075
+ $X2=0 $Y2=0
cc_768 N_SET_B_c_1111_n N_A_2501_543#_c_1246_n 0.0515588f $X=14 $Y=0.35 $X2=0
+ $Y2=0
cc_769 N_SET_B_c_1115_n N_A_2501_543#_c_1246_n 0.0107699f $X=14.085 $Y=1.425
+ $X2=0 $Y2=0
cc_770 N_SET_B_c_1115_n N_A_2501_543#_c_1247_n 0.022494f $X=14.085 $Y=1.425
+ $X2=0 $Y2=0
cc_771 N_SET_B_c_1160_p N_A_2501_543#_c_1247_n 0.013338f $X=14.17 $Y=1.535 $X2=0
+ $Y2=0
cc_772 N_SET_B_c_1160_p N_A_2501_543#_c_1248_n 0.0122858f $X=14.17 $Y=1.535
+ $X2=0 $Y2=0
cc_773 N_SET_B_c_1116_n N_A_2501_543#_c_1248_n 0.0461731f $X=14.68 $Y=1.56 $X2=0
+ $Y2=0
cc_774 N_SET_B_M1010_g N_A_2501_543#_c_1248_n 0.0269771f $X=14.745 $Y=1.075
+ $X2=0 $Y2=0
cc_775 N_SET_B_M1010_g N_A_2501_543#_c_1267_n 0.0403919f $X=14.745 $Y=1.075
+ $X2=0 $Y2=0
cc_776 N_SET_B_M1010_g N_A_2501_543#_c_1268_n 0.0181155f $X=14.745 $Y=1.075
+ $X2=0 $Y2=0
cc_777 N_SET_B_c_1116_n N_A_2501_543#_c_1308_n 0.0092914f $X=14.68 $Y=1.56 $X2=0
+ $Y2=0
cc_778 N_SET_B_M1010_g N_A_2501_543#_c_1308_n 0.00220264f $X=14.745 $Y=1.075
+ $X2=0 $Y2=0
cc_779 N_SET_B_c_1111_n N_A_2501_543#_c_1249_n 0.0211167f $X=14 $Y=0.35 $X2=0
+ $Y2=0
cc_780 SET_B N_A_2501_543#_c_1249_n 0.0331062f $X=12.155 $Y=1.21 $X2=0 $Y2=0
cc_781 N_SET_B_M1010_g N_VPWR_c_1434_n 0.00557214f $X=14.745 $Y=1.075 $X2=0
+ $Y2=0
cc_782 N_SET_B_M1018_g N_VPWR_c_1443_n 0.00413607f $X=10.65 $Y=2.99 $X2=0 $Y2=0
cc_783 N_SET_B_M1010_g N_VPWR_c_1443_n 0.0156697f $X=14.745 $Y=1.075 $X2=0 $Y2=0
cc_784 N_SET_B_c_1119_n N_VGND_M1038_d 0.00229266f $X=12.185 $Y=1.295 $X2=-0.33
+ $Y2=-0.265
cc_785 N_SET_B_M1038_g N_VGND_c_1727_n 0.0553397f $X=10.845 $Y=0.745 $X2=0 $Y2=0
cc_786 N_SET_B_c_1119_n N_VGND_c_1727_n 0.0653018f $X=12.185 $Y=1.295 $X2=0
+ $Y2=0
cc_787 N_SET_B_c_1111_n N_VGND_c_1729_n 0.00489946f $X=14 $Y=0.35 $X2=0 $Y2=0
cc_788 N_SET_B_c_1115_n N_VGND_c_1729_n 0.0603749f $X=14.085 $Y=1.425 $X2=0
+ $Y2=0
cc_789 N_SET_B_c_1116_n N_VGND_c_1729_n 0.0350984f $X=14.68 $Y=1.56 $X2=0 $Y2=0
cc_790 N_SET_B_M1010_g N_VGND_c_1729_n 0.0497567f $X=14.745 $Y=1.075 $X2=0 $Y2=0
cc_791 N_SET_B_c_1111_n N_VGND_c_1735_n 0.0652481f $X=14 $Y=0.35 $X2=0 $Y2=0
cc_792 N_SET_B_c_1113_n N_VGND_c_1735_n 0.00923655f $X=12.355 $Y=0.35 $X2=0
+ $Y2=0
cc_793 N_SET_B_c_1115_n N_VGND_c_1735_n 0.0164973f $X=14.085 $Y=1.425 $X2=0
+ $Y2=0
cc_794 SET_B N_VGND_c_1735_n 0.023215f $X=12.155 $Y=1.21 $X2=0 $Y2=0
cc_795 N_SET_B_c_1119_n N_VGND_c_1735_n 0.0332178f $X=12.185 $Y=1.295 $X2=0
+ $Y2=0
cc_796 N_SET_B_c_1119_n A_2394_107# 0.00191361f $X=12.185 $Y=1.295 $X2=0 $Y2=0
cc_797 N_A_2729_463#_c_1194_n N_A_2501_543#_c_1238_n 0.0155952f $X=15.895
+ $Y=1.075 $X2=0.24 $Y2=0
cc_798 N_A_2729_463#_c_1194_n N_A_2501_543#_c_1251_n 0.0172717f $X=15.895
+ $Y=1.075 $X2=0 $Y2=0
cc_799 N_A_2729_463#_c_1194_n N_A_2501_543#_c_1242_n 0.0349723f $X=15.895
+ $Y=1.075 $X2=0 $Y2=0
cc_800 N_A_2729_463#_c_1197_n N_A_2501_543#_c_1244_n 0.018576f $X=15.685 $Y=2.26
+ $X2=0 $Y2=0
cc_801 N_A_2729_463#_c_1194_n N_A_2501_543#_c_1244_n 0.0482003f $X=15.895
+ $Y=1.075 $X2=0 $Y2=0
cc_802 N_A_2729_463#_M1009_g N_A_2501_543#_c_1246_n 5.09458e-19 $X=14.035
+ $Y=1.075 $X2=0 $Y2=0
cc_803 N_A_2729_463#_M1009_g N_A_2501_543#_c_1247_n 0.0100864f $X=14.035
+ $Y=1.075 $X2=0 $Y2=0
cc_804 N_A_2729_463#_c_1196_n N_A_2501_543#_c_1265_n 0.0135019f $X=13.965
+ $Y=2.605 $X2=0 $Y2=0
cc_805 N_A_2729_463#_c_1197_n N_A_2501_543#_c_1265_n 0.0127031f $X=15.685
+ $Y=2.26 $X2=0 $Y2=0
cc_806 N_A_2729_463#_M1009_g N_A_2501_543#_c_1265_n 0.0100466f $X=14.035
+ $Y=1.075 $X2=0 $Y2=0
cc_807 N_A_2729_463#_c_1196_n N_A_2501_543#_c_1248_n 7.48832e-19 $X=13.965
+ $Y=2.605 $X2=0 $Y2=0
cc_808 N_A_2729_463#_c_1197_n N_A_2501_543#_c_1248_n 0.0860625f $X=15.685
+ $Y=2.26 $X2=0 $Y2=0
cc_809 N_A_2729_463#_M1009_g N_A_2501_543#_c_1248_n 0.0327315f $X=14.035
+ $Y=1.075 $X2=0 $Y2=0
cc_810 N_A_2729_463#_c_1196_n N_A_2501_543#_c_1267_n 0.0260497f $X=13.965
+ $Y=2.605 $X2=0 $Y2=0
cc_811 N_A_2729_463#_c_1197_n N_A_2501_543#_c_1267_n 0.102622f $X=15.685 $Y=2.26
+ $X2=0 $Y2=0
cc_812 N_A_2729_463#_c_1197_n N_A_2501_543#_c_1327_n 0.0248971f $X=15.685
+ $Y=2.26 $X2=0 $Y2=0
cc_813 N_A_2729_463#_c_1194_n N_A_2501_543#_c_1327_n 0.0126759f $X=15.895
+ $Y=1.075 $X2=0 $Y2=0
cc_814 N_A_2729_463#_c_1194_n N_A_2501_543#_c_1308_n 0.0280159f $X=15.895
+ $Y=1.075 $X2=0 $Y2=0
cc_815 N_A_2729_463#_c_1196_n N_A_2501_543#_c_1270_n 0.00493352f $X=13.965
+ $Y=2.605 $X2=0 $Y2=0
cc_816 N_A_2729_463#_c_1196_n N_VPWR_c_1434_n 0.0411583f $X=13.965 $Y=2.605
+ $X2=0 $Y2=0
cc_817 N_A_2729_463#_c_1197_n N_VPWR_c_1437_n 0.0215853f $X=15.685 $Y=2.26 $X2=0
+ $Y2=0
cc_818 N_A_2729_463#_c_1194_n N_VGND_c_1729_n 0.019489f $X=15.895 $Y=1.075 $X2=0
+ $Y2=0
cc_819 N_A_2729_463#_M1009_g N_VGND_c_1729_n 0.00417503f $X=14.035 $Y=1.075
+ $X2=0 $Y2=0
cc_820 N_A_2729_463#_c_1194_n N_VGND_c_1731_n 0.0379441f $X=15.895 $Y=1.075
+ $X2=0 $Y2=0
cc_821 N_A_2729_463#_c_1194_n N_VGND_c_1735_n 0.0181496f $X=15.895 $Y=1.075
+ $X2=0 $Y2=0
cc_822 N_A_2729_463#_M1009_g N_VGND_c_1735_n 0.0108445f $X=14.035 $Y=1.075 $X2=0
+ $Y2=0
cc_823 N_A_2501_543#_M1026_g N_A_3609_173#_c_1378_n 0.00174457f $X=17.18 $Y=0.91
+ $X2=0 $Y2=0
cc_824 N_A_2501_543#_M1034_g N_A_3609_173#_c_1378_n 0.0229914f $X=18.58 $Y=1.075
+ $X2=0 $Y2=0
cc_825 N_A_2501_543#_c_1252_n N_A_3609_173#_c_1383_n 0.00224645f $X=17.23
+ $Y=2.095 $X2=0 $Y2=0
cc_826 N_A_2501_543#_c_1241_n N_A_3609_173#_c_1383_n 0.0243753f $X=18.33
+ $Y=1.845 $X2=0 $Y2=0
cc_827 N_A_2501_543#_M1032_g N_A_3609_173#_c_1383_n 0.0354815f $X=18.58 $Y=2.77
+ $X2=0 $Y2=0
cc_828 N_A_2501_543#_c_1245_n N_A_3609_173#_c_1383_n 0.019714f $X=18.58 $Y=1.845
+ $X2=0 $Y2=0
cc_829 N_A_2501_543#_M1034_g N_A_3609_173#_c_1379_n 0.0173827f $X=18.58 $Y=1.075
+ $X2=0 $Y2=0
cc_830 N_A_2501_543#_c_1245_n N_A_3609_173#_c_1379_n 0.0257198f $X=18.58
+ $Y=1.845 $X2=0 $Y2=0
cc_831 N_A_2501_543#_M1026_g N_A_3609_173#_c_1380_n 3.47071e-19 $X=17.18 $Y=0.91
+ $X2=0 $Y2=0
cc_832 N_A_2501_543#_c_1241_n N_A_3609_173#_c_1380_n 0.00903649f $X=18.33
+ $Y=1.845 $X2=0 $Y2=0
cc_833 N_A_2501_543#_M1034_g N_A_3609_173#_c_1380_n 0.00200762f $X=18.58
+ $Y=1.075 $X2=0 $Y2=0
cc_834 N_A_2501_543#_c_1245_n N_A_3609_173#_c_1398_n 0.00336651f $X=18.58
+ $Y=1.845 $X2=10.08 $Y2=0
cc_835 N_A_2501_543#_M1034_g N_A_3609_173#_M1003_g 0.0642893f $X=18.58 $Y=1.075
+ $X2=0 $Y2=0
cc_836 N_A_2501_543#_c_1260_n N_VPWR_c_1431_n 0.005385f $X=12.68 $Y=2.84 $X2=0
+ $Y2=0
cc_837 N_A_2501_543#_c_1260_n N_VPWR_c_1434_n 0.0224808f $X=12.68 $Y=2.84 $X2=0
+ $Y2=0
cc_838 N_A_2501_543#_c_1263_n N_VPWR_c_1434_n 0.00662568f $X=13.585 $Y=2.61
+ $X2=0 $Y2=0
cc_839 N_A_2501_543#_c_1267_n N_VPWR_c_1434_n 0.0494826f $X=14.97 $Y=2.61 $X2=0
+ $Y2=0
cc_840 N_A_2501_543#_c_1268_n N_VPWR_c_1434_n 0.00533851f $X=15.135 $Y=2.925
+ $X2=0 $Y2=0
cc_841 N_A_2501_543#_c_1270_n N_VPWR_c_1434_n 0.0117176f $X=13.67 $Y=2.61 $X2=0
+ $Y2=0
cc_842 N_A_2501_543#_c_1251_n N_VPWR_c_1437_n 0.0645116f $X=16.355 $Y=2.095
+ $X2=0 $Y2=0
cc_843 N_A_2501_543#_c_1252_n N_VPWR_c_1437_n 0.0671556f $X=17.23 $Y=2.095 $X2=0
+ $Y2=0
cc_844 N_A_2501_543#_c_1242_n N_VPWR_c_1437_n 0.00987893f $X=17.48 $Y=1.845
+ $X2=0 $Y2=0
cc_845 N_A_2501_543#_M1032_g N_VPWR_c_1440_n 0.0779387f $X=18.58 $Y=2.77 $X2=0
+ $Y2=0
cc_846 N_A_2501_543#_M1037_d N_VPWR_c_1443_n 3.33633e-19 $X=12.505 $Y=2.715
+ $X2=0 $Y2=0
cc_847 N_A_2501_543#_c_1252_n N_VPWR_c_1443_n 0.0138762f $X=17.23 $Y=2.095 $X2=0
+ $Y2=0
cc_848 N_A_2501_543#_M1032_g N_VPWR_c_1443_n 0.00649418f $X=18.58 $Y=2.77 $X2=0
+ $Y2=0
cc_849 N_A_2501_543#_c_1260_n N_VPWR_c_1443_n 0.0481068f $X=12.68 $Y=2.84 $X2=0
+ $Y2=0
cc_850 N_A_2501_543#_c_1268_n N_VPWR_c_1443_n 0.0168517f $X=15.135 $Y=2.925
+ $X2=0 $Y2=0
cc_851 N_A_2501_543#_M1026_g N_Q_N_c_1685_n 0.0368755f $X=17.18 $Y=0.91 $X2=0
+ $Y2=0
cc_852 N_A_2501_543#_c_1252_n N_Q_N_c_1685_n 0.0425437f $X=17.23 $Y=2.095 $X2=0
+ $Y2=0
cc_853 N_A_2501_543#_c_1241_n N_Q_N_c_1685_n 0.0346906f $X=18.33 $Y=1.845 $X2=0
+ $Y2=0
cc_854 N_A_2501_543#_c_1242_n N_Q_N_c_1685_n 0.0277525f $X=17.48 $Y=1.845 $X2=0
+ $Y2=0
cc_855 N_A_2501_543#_M1034_g N_Q_N_c_1685_n 0.00483836f $X=18.58 $Y=1.075 $X2=0
+ $Y2=0
cc_856 N_A_2501_543#_M1032_g N_Q_N_c_1685_n 0.00555907f $X=18.58 $Y=2.77 $X2=0
+ $Y2=0
cc_857 N_A_2501_543#_c_1244_n N_VGND_c_1729_n 0.00270203f $X=16.035 $Y=1.745
+ $X2=0 $Y2=0
cc_858 N_A_2501_543#_c_1248_n N_VGND_c_1729_n 0.010531f $X=15.215 $Y=1.91 $X2=0
+ $Y2=0
cc_859 N_A_2501_543#_c_1308_n N_VGND_c_1729_n 0.00688253f $X=15.38 $Y=1.57 $X2=0
+ $Y2=0
cc_860 N_A_2501_543#_c_1238_n N_VGND_c_1731_n 0.0586104f $X=16.285 $Y=1.395
+ $X2=0 $Y2=0
cc_861 N_A_2501_543#_M1026_g N_VGND_c_1731_n 0.0596742f $X=17.18 $Y=0.91 $X2=0
+ $Y2=0
cc_862 N_A_2501_543#_c_1242_n N_VGND_c_1731_n 0.00909434f $X=17.48 $Y=1.845
+ $X2=0 $Y2=0
cc_863 N_A_2501_543#_M1034_g N_VGND_c_1733_n 0.0476742f $X=18.58 $Y=1.075 $X2=0
+ $Y2=0
cc_864 N_A_2501_543#_c_1238_n N_VGND_c_1735_n 0.00672879f $X=16.285 $Y=1.395
+ $X2=0 $Y2=0
cc_865 N_A_2501_543#_M1026_g N_VGND_c_1735_n 0.0139641f $X=17.18 $Y=0.91 $X2=0
+ $Y2=0
cc_866 N_A_2501_543#_M1034_g N_VGND_c_1735_n 0.00672879f $X=18.58 $Y=1.075 $X2=0
+ $Y2=0
cc_867 N_A_2501_543#_c_1246_n N_VGND_c_1735_n 0.0352103f $X=13.585 $Y=0.7 $X2=0
+ $Y2=0
cc_868 N_A_2501_543#_c_1249_n N_VGND_c_1735_n 0.0228422f $X=12.82 $Y=0.7 $X2=0
+ $Y2=0
cc_869 N_A_2501_543#_c_1247_n A_2715_173# 0.00170567f $X=13.67 $Y=1.825 $X2=0
+ $Y2=0
cc_870 N_A_3609_173#_c_1383_n N_VPWR_c_1440_n 0.0629871f $X=18.19 $Y=2.52 $X2=0
+ $Y2=0
cc_871 N_A_3609_173#_c_1398_n N_VPWR_c_1440_n 0.019212f $X=19.41 $Y=1.67 $X2=0
+ $Y2=0
cc_872 N_A_3609_173#_M1003_g N_VPWR_c_1440_n 0.0613135f $X=19.475 $Y=0.91 $X2=0
+ $Y2=0
cc_873 N_A_3609_173#_c_1383_n N_VPWR_c_1443_n 0.0170977f $X=18.19 $Y=2.52 $X2=0
+ $Y2=0
cc_874 N_A_3609_173#_M1003_g N_VPWR_c_1443_n 0.0145323f $X=19.475 $Y=0.91 $X2=0
+ $Y2=0
cc_875 N_A_3609_173#_c_1378_n N_Q_N_c_1685_n 0.0449641f $X=18.19 $Y=1.075 $X2=0
+ $Y2=0
cc_876 N_A_3609_173#_c_1383_n N_Q_N_c_1685_n 0.0962874f $X=18.19 $Y=2.52 $X2=0
+ $Y2=0
cc_877 N_A_3609_173#_c_1380_n N_Q_N_c_1685_n 0.0112061f $X=18.19 $Y=1.59 $X2=0
+ $Y2=0
cc_878 N_A_3609_173#_c_1398_n Q 0.0416943f $X=19.41 $Y=1.67 $X2=0 $Y2=0
cc_879 N_A_3609_173#_M1003_g Q 0.0356954f $X=19.475 $Y=0.91 $X2=0 $Y2=0
cc_880 N_A_3609_173#_M1003_g Q 0.0176721f $X=19.475 $Y=0.91 $X2=0 $Y2=0
cc_881 N_A_3609_173#_M1003_g N_Q_c_1704_n 0.0143814f $X=19.475 $Y=0.91 $X2=0
+ $Y2=0
cc_882 N_A_3609_173#_M1003_g Q 0.00506627f $X=19.475 $Y=0.91 $X2=0 $Y2=0
cc_883 N_A_3609_173#_c_1378_n N_VGND_c_1733_n 0.0379441f $X=18.19 $Y=1.075 $X2=0
+ $Y2=0
cc_884 N_A_3609_173#_c_1379_n N_VGND_c_1733_n 0.0548452f $X=19.245 $Y=1.59 $X2=0
+ $Y2=0
cc_885 N_A_3609_173#_c_1398_n N_VGND_c_1733_n 0.0192928f $X=19.41 $Y=1.67 $X2=0
+ $Y2=0
cc_886 N_A_3609_173#_M1003_g N_VGND_c_1733_n 0.0500693f $X=19.475 $Y=0.91 $X2=0
+ $Y2=0
cc_887 N_A_3609_173#_c_1378_n N_VGND_c_1735_n 0.0181496f $X=18.19 $Y=1.075 $X2=0
+ $Y2=0
cc_888 N_A_3609_173#_M1003_g N_VGND_c_1735_n 0.0136923f $X=19.475 $Y=0.91 $X2=0
+ $Y2=0
cc_889 N_VPWR_c_1443_n N_A_485_569#_c_1583_n 0.0195412f $X=19.37 $Y=3.59
+ $X2=19.92 $Y2=4.07
cc_890 N_VPWR_c_1422_n N_A_485_569#_c_1544_n 0.00461347f $X=4.22 $Y=2.97 $X2=0
+ $Y2=0
cc_891 N_VPWR_c_1422_n N_A_485_569#_c_1546_n 0.0677529f $X=4.22 $Y=2.97 $X2=0
+ $Y2=0
cc_892 N_VPWR_c_1422_n N_A_485_569#_c_1606_n 0.0321966f $X=4.22 $Y=2.97 $X2=0
+ $Y2=0
cc_893 N_VPWR_c_1443_n N_A_485_569#_c_1606_n 0.0199629f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_894 N_VPWR_c_1425_n N_A_485_569#_c_1547_n 0.00479486f $X=5.78 $Y=2.565 $X2=0
+ $Y2=0
cc_895 N_VPWR_c_1443_n N_A_485_569#_c_1547_n 0.033543f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_896 N_VPWR_c_1422_n N_A_485_569#_c_1550_n 0.00461913f $X=4.22 $Y=2.97 $X2=0
+ $Y2=0
cc_897 N_VPWR_c_1443_n N_A_485_569#_c_1550_n 0.00754921f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_898 N_VPWR_c_1425_n N_A_485_569#_c_1553_n 0.0871892f $X=5.78 $Y=2.565 $X2=0
+ $Y2=0
cc_899 N_VPWR_c_1443_n N_A_485_569#_c_1553_n 0.0214561f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_900 N_VPWR_c_1425_n N_A_485_569#_c_1554_n 0.0136256f $X=5.78 $Y=2.565 $X2=0
+ $Y2=0
cc_901 N_VPWR_c_1425_n N_A_485_569#_c_1556_n 0.0408796f $X=5.78 $Y=2.565 $X2=0
+ $Y2=0
cc_902 N_VPWR_c_1443_n N_A_485_569#_c_1557_n 0.0767071f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_903 N_VPWR_c_1425_n N_A_485_569#_c_1560_n 0.0123381f $X=5.78 $Y=2.565 $X2=0
+ $Y2=0
cc_904 N_VPWR_c_1443_n N_A_485_569#_c_1560_n 0.010882f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_905 N_VPWR_c_1443_n N_A_485_569#_c_1565_n 0.0182755f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_906 N_VPWR_c_1428_n A_1710_556# 0.00448957f $X=9.4 $Y=3.06 $X2=0 $Y2=3.985
cc_907 N_VPWR_c_1431_n A_2359_543# 0.00538136f $X=11.79 $Y=3.59 $X2=0 $Y2=3.985
cc_908 N_VPWR_c_1443_n A_2359_543# 9.79604e-19 $X=19.37 $Y=3.59 $X2=0 $Y2=3.985
cc_909 N_VPWR_c_1434_n A_2687_543# 0.00482885f $X=14.285 $Y=2.985 $X2=0
+ $Y2=3.985
cc_910 N_VPWR_c_1437_n N_Q_N_c_1685_n 0.097785f $X=16.84 $Y=2.36 $X2=10.08
+ $Y2=4.07
cc_911 N_VPWR_c_1443_n N_Q_N_c_1685_n 0.0499636f $X=19.37 $Y=3.59 $X2=10.08
+ $Y2=4.07
cc_912 N_VPWR_c_1443_n Q 0.015253f $X=19.37 $Y=3.59 $X2=0.24 $Y2=4.07
cc_913 N_VPWR_c_1440_n Q 0.0711583f $X=19.085 $Y=2.52 $X2=0 $Y2=0
cc_914 N_A_485_569#_c_1537_n N_VGND_c_1721_n 0.0021618f $X=3.135 $Y=0.83 $X2=0
+ $Y2=0
cc_915 N_A_485_569#_M1007_s N_VGND_c_1735_n 0.00225203f $X=6.78 $Y=0.6 $X2=0
+ $Y2=0
cc_916 N_A_485_569#_c_1537_n N_VGND_c_1735_n 0.0191245f $X=3.135 $Y=0.83 $X2=0
+ $Y2=0
cc_917 N_A_485_569#_c_1539_n N_VGND_c_1735_n 0.0112819f $X=6.925 $Y=0.835 $X2=0
+ $Y2=0
cc_918 N_A_485_569#_c_1540_n N_VGND_c_1735_n 0.0303718f $X=2.59 $Y=0.745 $X2=0
+ $Y2=0
cc_919 N_A_485_569#_c_1537_n A_646_107# 0.00213576f $X=3.135 $Y=0.83 $X2=0 $Y2=0
cc_920 N_A_485_569#_c_1538_n A_646_107# 3.29858e-19 $X=3.22 $Y=2.455 $X2=0 $Y2=0
cc_921 N_Q_N_c_1685_n N_VGND_c_1731_n 0.053125f $X=17.57 $Y=0.66 $X2=0 $Y2=0
cc_922 N_Q_N_c_1685_n N_VGND_c_1735_n 0.0390307f $X=17.57 $Y=0.66 $X2=0 $Y2=0
cc_923 N_Q_c_1704_n N_VGND_c_1733_n 0.0526655f $X=19.865 $Y=0.66 $X2=0 $Y2=0
cc_924 N_Q_c_1704_n N_VGND_c_1735_n 0.0338855f $X=19.865 $Y=0.66 $X2=0 $Y2=0
cc_925 N_VGND_c_1735_n A_348_107# 0.00261802f $X=19.37 $Y=0.48 $X2=0 $Y2=0
cc_926 N_VGND_c_1735_n A_646_107# 0.00624885f $X=19.37 $Y=0.48 $X2=0 $Y2=0
cc_927 N_VGND_c_1725_n A_1669_120# 0.00491355f $X=8.525 $Y=0.48 $X2=0 $Y2=0
cc_928 N_VGND_c_1735_n A_1669_120# 0.00275248f $X=19.37 $Y=0.48 $X2=0 $Y2=0
cc_929 N_VGND_c_1735_n A_2077_107# 0.00224881f $X=19.37 $Y=0.48 $X2=0 $Y2=0
cc_930 N_VGND_c_1735_n A_2394_107# 0.00297013f $X=19.37 $Y=0.48 $X2=0 $Y2=0
cc_931 N_VGND_c_1729_n A_2857_173# 0.0042905f $X=14.465 $Y=0.48 $X2=0 $Y2=0
