# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__dlxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dlxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.795000 3.100000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.700000 0.515000 8.050000 3.755000 ;
    END
  END Q
  PIN GATE
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.540000 1.175000 0.870000 1.725000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 8.160000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 8.160000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 8.160000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 8.160000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.985000 8.160000 4.155000 ;
      RECT 0.110000  0.495000 0.665000 0.995000 ;
      RECT 0.110000  0.995000 0.360000 1.905000 ;
      RECT 0.110000  1.905000 1.795000 2.015000 ;
      RECT 0.110000  2.015000 1.780000 2.075000 ;
      RECT 0.110000  2.075000 0.360000 2.985000 ;
      RECT 0.540000  2.255000 1.430000 3.705000 ;
      RECT 0.845000  0.365000 1.795000 0.995000 ;
      RECT 1.540000  1.345000 1.795000 1.905000 ;
      RECT 1.610000  2.075000 1.780000 2.645000 ;
      RECT 1.610000  2.645000 3.190000 2.815000 ;
      RECT 1.890000  2.995000 2.840000 3.705000 ;
      RECT 1.960000  2.195000 2.290000 2.465000 ;
      RECT 1.975000  0.515000 2.225000 1.445000 ;
      RECT 1.975000  1.445000 3.880000 1.615000 ;
      RECT 1.975000  1.615000 2.290000 2.195000 ;
      RECT 2.405000  0.365000 2.995000 0.975000 ;
      RECT 3.020000  2.815000 3.190000 3.635000 ;
      RECT 3.020000  3.635000 4.050000 3.805000 ;
      RECT 3.225000  0.495000 3.555000 0.995000 ;
      RECT 3.370000  2.165000 4.230000 2.335000 ;
      RECT 3.370000  2.335000 3.540000 2.895000 ;
      RECT 3.370000  2.895000 3.700000 3.455000 ;
      RECT 3.385000  0.995000 3.555000 1.095000 ;
      RECT 3.385000  1.095000 4.230000 1.265000 ;
      RECT 3.550000  1.615000 3.880000 1.985000 ;
      RECT 3.720000  2.515000 4.740000 2.715000 ;
      RECT 3.880000  2.715000 4.050000 3.635000 ;
      RECT 4.005000  0.495000 4.335000 0.745000 ;
      RECT 4.005000  0.745000 5.090000 0.915000 ;
      RECT 4.060000  1.265000 4.230000 2.165000 ;
      RECT 4.230000  2.895000 5.090000 3.065000 ;
      RECT 4.230000  3.065000 4.480000 3.725000 ;
      RECT 4.410000  1.095000 4.740000 2.515000 ;
      RECT 4.920000  0.915000 5.090000 1.835000 ;
      RECT 4.920000  1.835000 6.680000 2.005000 ;
      RECT 4.920000  2.005000 5.090000 2.895000 ;
      RECT 5.270000  0.365000 5.860000 0.895000 ;
      RECT 5.270000  2.895000 6.220000 3.705000 ;
      RECT 5.430000  1.075000 5.760000 1.425000 ;
      RECT 5.430000  1.425000 7.030000 1.595000 ;
      RECT 5.430000  1.595000 5.760000 1.655000 ;
      RECT 6.025000  2.185000 7.030000 2.355000 ;
      RECT 6.025000  2.355000 6.355000 2.675000 ;
      RECT 6.045000  0.845000 6.375000 1.425000 ;
      RECT 6.350000  1.775000 6.680000 1.835000 ;
      RECT 6.535000  2.535000 7.485000 3.755000 ;
      RECT 6.555000  0.365000 7.505000 1.245000 ;
      RECT 6.860000  1.595000 7.030000 2.185000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.540000  3.505000 0.710000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.875000  0.395000 1.045000 0.565000 ;
      RECT 0.900000  3.505000 1.070000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.235000  0.395000 1.405000 0.565000 ;
      RECT 1.260000  3.505000 1.430000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  0.395000 1.765000 0.565000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.920000  3.505000 2.090000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.280000  3.505000 2.450000 3.675000 ;
      RECT 2.435000  0.395000 2.605000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.640000  3.505000 2.810000 3.675000 ;
      RECT 2.795000  0.395000 2.965000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 5.300000  0.395000 5.470000 0.565000 ;
      RECT 5.300000  3.505000 5.470000 3.675000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.985000 5.605000 4.155000 ;
      RECT 5.660000  0.395000 5.830000 0.565000 ;
      RECT 5.660000  3.505000 5.830000 3.675000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.985000 6.085000 4.155000 ;
      RECT 6.020000  3.505000 6.190000 3.675000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.985000 6.565000 4.155000 ;
      RECT 6.565000  3.505000 6.735000 3.675000 ;
      RECT 6.585000  0.395000 6.755000 0.565000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.985000 7.045000 4.155000 ;
      RECT 6.925000  3.505000 7.095000 3.675000 ;
      RECT 6.945000  0.395000 7.115000 0.565000 ;
      RECT 7.285000  3.505000 7.455000 3.675000 ;
      RECT 7.305000  0.395000 7.475000 0.565000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
  END
END sky130_fd_sc_hvl__dlxtp_1
END LIBRARY
