* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__nand3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 VGND C a_243_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_385_107# A Y VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_243_107# B a_385_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends
