* File: sky130_fd_sc_hvl__buf_1.pex.spice
* Created: Wed Sep  2 09:03:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__BUF_1%VNB 5 7 11 25
r17 7 25 5.20833e-05 $w=2.4e-06 $l=1e-09 $layer=MET1_cond $X=1.2 $Y=0.057
+ $X2=1.2 $Y2=0.058
r18 7 11 0.00296875 $w=2.4e-06 $l=5.7e-08 $layer=MET1_cond $X=1.2 $Y=0.057
+ $X2=1.2 $Y2=0
r19 5 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r20 5 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_1%VPB 4 6 14 21
r18 10 21 0.00296875 $w=2.4e-06 $l=5.7e-08 $layer=MET1_cond $X=1.2 $Y=4.07
+ $X2=1.2 $Y2=4.013
r19 10 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=4.07
+ $X2=2.16 $Y2=4.07
r20 9 14 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=2.16 $Y2=4.07
r21 9 10 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r22 6 21 5.20833e-05 $w=2.4e-06 $l=1e-09 $layer=MET1_cond $X=1.2 $Y=4.012
+ $X2=1.2 $Y2=4.013
r23 4 14 72.8 $w=1.7e-07 $l=2.20209e-06 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=2.16 $Y2=4.07
r24 4 9 72.8 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_1%A_84_81# 1 2 9 12 16 17 19 20 23 27 29 31
r47 25 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=1.285 $X2=2.1
+ $Y2=1.2
r48 25 27 48.6331 $w=2.48e-07 $l=1.055e-06 $layer=LI1_cond $X=2.1 $Y=1.285
+ $X2=2.1 $Y2=2.34
r49 21 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=1.115 $X2=2.1
+ $Y2=1.2
r50 21 23 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.1 $Y=1.115 $X2=2.1
+ $Y2=0.745
r51 19 29 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.975 $Y=1.2 $X2=2.1
+ $Y2=1.2
r52 19 20 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.975 $Y=1.2
+ $X2=1.005 $Y2=1.2
r53 17 32 29.6268 $w=6.05e-07 $l=3.15e-07 $layer=POLY_cond $X=0.722 $Y=1.58
+ $X2=0.722 $Y2=1.895
r54 17 31 18.1303 $w=6.05e-07 $l=1.85e-07 $layer=POLY_cond $X=0.722 $Y=1.58
+ $X2=0.722 $Y2=1.395
r55 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.84
+ $Y=1.58 $X2=0.84 $Y2=1.58
r56 14 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.84 $Y=1.285
+ $X2=1.005 $Y2=1.2
r57 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.84 $Y=1.285
+ $X2=0.84 $Y2=1.58
r58 12 32 114.496 $w=5e-07 $l=1.07e-06 $layer=POLY_cond $X=0.775 $Y=2.965
+ $X2=0.775 $Y2=1.895
r59 9 31 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.67 $Y=0.91 $X2=0.67
+ $Y2=1.395
r60 2 27 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=2.215 $X2=2.06 $Y2=2.34
r61 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.535 $X2=2.06 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_1%A 1 2 3 4 5 12 16 18
r21 15 18 111.286 $w=5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.67 $Y=1.55 $X2=1.67
+ $Y2=2.59
r22 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.63
+ $Y=1.55 $X2=1.63 $Y2=1.55
r23 12 15 86.1397 $w=5e-07 $l=8.05e-07 $layer=POLY_cond $X=1.67 $Y=0.745
+ $X2=1.67 $Y2=1.55
r24 4 5 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=2.775 $X2=1.63
+ $Y2=3.145
r25 3 4 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=2.405 $X2=1.63
+ $Y2=2.775
r26 2 3 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=2.035 $X2=1.63
+ $Y2=2.405
r27 1 2 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=1.665 $X2=1.63
+ $Y2=2.035
r28 1 16 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.63 $Y=1.665
+ $X2=1.63 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_1%X 1 2 7 8 9 10 11 12 13 24 36 46
r18 46 47 6.43827 $w=4.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.332 $Y=2.34
+ $X2=0.332 $Y2=2.175
r19 34 36 0.344408 $w=4.33e-07 $l=1.3e-08 $layer=LI1_cond $X=0.332 $Y=2.392
+ $X2=0.332 $Y2=2.405
r20 13 43 11.7894 $w=4.33e-07 $l=4.45e-07 $layer=LI1_cond $X=0.332 $Y=3.145
+ $X2=0.332 $Y2=3.59
r21 12 13 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.332 $Y=2.775
+ $X2=0.332 $Y2=3.145
r22 11 34 0.953746 $w=4.33e-07 $l=3.6e-08 $layer=LI1_cond $X=0.332 $Y=2.356
+ $X2=0.332 $Y2=2.392
r23 11 46 0.423887 $w=4.33e-07 $l=1.6e-08 $layer=LI1_cond $X=0.332 $Y=2.356
+ $X2=0.332 $Y2=2.34
r24 11 12 8.84864 $w=4.33e-07 $l=3.34e-07 $layer=LI1_cond $X=0.332 $Y=2.441
+ $X2=0.332 $Y2=2.775
r25 11 36 0.953746 $w=4.33e-07 $l=3.6e-08 $layer=LI1_cond $X=0.332 $Y=2.441
+ $X2=0.332 $Y2=2.405
r26 10 47 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.175
r27 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=2.035
r28 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295 $X2=0.24
+ $Y2=1.665
r29 7 8 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925 $X2=0.24
+ $Y2=1.295
r30 7 24 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=0.68
r31 2 46 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.24
+ $Y=2.215 $X2=0.385 $Y2=2.34
r32 2 43 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.24
+ $Y=2.215 $X2=0.385 $Y2=3.59
r33 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.535 $X2=0.28 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_1%VPWR 1 4 7
r16 7 10 26.9387 $w=5.53e-07 $l=1.25e-06 $layer=LI1_cond $X=1.007 $Y=2.34
+ $X2=1.007 $Y2=3.59
r17 4 10 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.185 $Y=3.59
+ $X2=1.185 $Y2=3.59
r18 1 10 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.025
+ $Y=2.215 $X2=1.165 $Y2=3.59
r19 1 7 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.025
+ $Y=2.215 $X2=1.165 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_1%VGND 1 4 7
r21 7 13 2.684 $w=1.248e-06 $l=2.75e-07 $layer=LI1_cond $X=1.17 $Y=0.48 $X2=1.17
+ $Y2=0.755
r22 7 8 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.71 $Y=0.48 $X2=1.71
+ $Y2=0.48
r23 7 8 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.63 $Y=0.48 $X2=0.63
+ $Y2=0.48
r24 4 8 0.00208333 $w=2.4e-06 $l=4e-08 $layer=MET1_cond $X=1.2 $Y=0.44 $X2=1.2
+ $Y2=0.48
r25 1 13 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=0.92
+ $Y=0.535 $X2=1.06 $Y2=0.755
.ends

