* File: sky130_fd_sc_hvl__buf_4.pex.spice
* Created: Wed Sep  2 09:04:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__BUF_4%VNB 5 7 11 25
r32 7 25 2.60417e-05 $w=4.8e-06 $l=1e-09 $layer=MET1_cond $X=2.4 $Y=0.057
+ $X2=2.4 $Y2=0.058
r33 7 11 0.00148437 $w=4.8e-06 $l=5.7e-08 $layer=MET1_cond $X=2.4 $Y=0.057
+ $X2=2.4 $Y2=0
r34 5 11 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r35 5 11 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_4%VPB 4 6 14 21
r38 10 21 0.00148437 $w=4.8e-06 $l=5.7e-08 $layer=MET1_cond $X=2.4 $Y=4.07
+ $X2=2.4 $Y2=4.013
r39 10 14 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.56 $Y=4.07
+ $X2=4.56 $Y2=4.07
r40 9 14 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=4.56
+ $Y2=4.07
r41 9 10 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r42 6 21 2.60417e-05 $w=4.8e-06 $l=1e-09 $layer=MET1_cond $X=2.4 $Y=4.012
+ $X2=2.4 $Y2=4.013
r43 4 14 36.4 $w=1.7e-07 $l=4.6023e-06 $layer=licon1_NTAP_notbjt $count=5 $X=0
+ $Y=3.985 $X2=4.56 $Y2=4.07
r44 4 9 36.4 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=5 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_4%A_149_81# 1 2 9 13 17 21 25 29 33 37 39 44 48
+ 52 56 60 62
r103 67 68 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.555 $Y=1.665
+ $X2=3.335 $Y2=1.665
r104 66 67 83.4646 $w=5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.775 $Y=1.665
+ $X2=2.555 $Y2=1.665
r105 60 68 10.7006 $w=5e-07 $l=1e-07 $layer=POLY_cond $X=3.435 $Y=1.665
+ $X2=3.335 $Y2=1.665
r106 59 60 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.435
+ $Y=1.64 $X2=3.435 $Y2=1.64
r107 56 59 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.515 $Y=1.51
+ $X2=3.515 $Y2=1.64
r108 52 54 57.6222 $w=2.48e-07 $l=1.25e-06 $layer=LI1_cond $X=4.545 $Y=2.34
+ $X2=4.545 $Y2=3.59
r109 50 62 3.24686 $w=2.9e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.545 $Y=1.595
+ $X2=4.505 $Y2=1.51
r110 50 52 34.3428 $w=2.48e-07 $l=7.45e-07 $layer=LI1_cond $X=4.545 $Y=1.595
+ $X2=4.545 $Y2=2.34
r111 46 62 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.505 $Y=1.425
+ $X2=4.505 $Y2=1.51
r112 46 48 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=4.505 $Y=1.425
+ $X2=4.505 $Y2=0.66
r113 45 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=1.51
+ $X2=3.515 $Y2=1.51
r114 44 62 3.3199 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.34 $Y=1.51
+ $X2=4.505 $Y2=1.51
r115 44 45 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.34 $Y=1.51
+ $X2=3.6 $Y2=1.51
r116 42 66 4.28024 $w=5e-07 $l=4e-08 $layer=POLY_cond $X=1.735 $Y=1.665
+ $X2=1.775 $Y2=1.665
r117 42 63 79.1844 $w=5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.735 $Y=1.665
+ $X2=0.995 $Y2=1.665
r118 41 42 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=1.735
+ $Y=1.64 $X2=1.735 $Y2=1.64
r119 39 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=1.64
+ $X2=3.515 $Y2=1.64
r120 39 41 110.583 $w=1.68e-07 $l=1.695e-06 $layer=LI1_cond $X=3.43 $Y=1.64
+ $X2=1.735 $Y2=1.64
r121 35 68 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.335 $Y=1.915
+ $X2=3.335 $Y2=1.665
r122 35 37 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=3.335 $Y=1.915
+ $X2=3.335 $Y2=2.965
r123 31 68 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.335 $Y=1.415
+ $X2=3.335 $Y2=1.665
r124 31 33 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.335 $Y=1.415
+ $X2=3.335 $Y2=0.91
r125 27 67 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.555 $Y=1.915
+ $X2=2.555 $Y2=1.665
r126 27 29 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.555 $Y=1.915
+ $X2=2.555 $Y2=2.965
r127 23 67 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.555 $Y=1.415
+ $X2=2.555 $Y2=1.665
r128 23 25 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.555 $Y=1.415
+ $X2=2.555 $Y2=0.91
r129 19 66 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.775 $Y=1.915
+ $X2=1.775 $Y2=1.665
r130 19 21 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=1.775 $Y=1.915
+ $X2=1.775 $Y2=2.965
r131 15 66 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.775 $Y=1.415
+ $X2=1.775 $Y2=1.665
r132 15 17 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.775 $Y=1.415
+ $X2=1.775 $Y2=0.91
r133 11 63 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.995 $Y=1.915
+ $X2=0.995 $Y2=1.665
r134 11 13 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=0.995 $Y=1.915
+ $X2=0.995 $Y2=2.965
r135 7 63 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.995 $Y=1.415
+ $X2=0.995 $Y2=1.665
r136 7 9 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.995 $Y=1.415
+ $X2=0.995 $Y2=0.91
r137 2 54 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=4.365
+ $Y=2.215 $X2=4.505 $Y2=3.59
r138 2 52 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.365
+ $Y=2.215 $X2=4.505 $Y2=2.34
r139 1 48 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.365
+ $Y=0.535 $X2=4.505 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_4%A 1 4 8 10
r22 7 10 115.031 $w=5e-07 $l=1.075e-06 $layer=POLY_cond $X=4.115 $Y=1.89
+ $X2=4.115 $Y2=2.965
r23 7 8 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05 $Y=1.89
+ $X2=4.05 $Y2=1.89
r24 4 7 104.866 $w=5e-07 $l=9.8e-07 $layer=POLY_cond $X=4.115 $Y=0.91 $X2=4.115
+ $Y2=1.89
r25 1 8 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=4.05 $Y=2.035
+ $X2=4.05 $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_4%VPWR 1 2 3 10 13 23 33 40
r41 37 40 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.405 $Y=3.63
+ $X2=4.125 $Y2=3.63
r42 36 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.125 $Y=3.59
+ $X2=4.125 $Y2=3.59
r43 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.405 $Y=3.59
+ $X2=3.405 $Y2=3.59
r44 33 36 15.4747 $w=9.48e-07 $l=1.205e-06 $layer=LI1_cond $X=3.765 $Y=2.385
+ $X2=3.765 $Y2=3.59
r45 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.765 $Y=3.59
+ $X2=1.765 $Y2=3.59
r46 23 26 16.0526 $w=9.48e-07 $l=1.25e-06 $layer=LI1_cond $X=2.125 $Y=2.34
+ $X2=2.125 $Y2=3.59
r47 20 27 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=0.925 $Y=3.63
+ $X2=1.765 $Y2=3.63
r48 17 20 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.205 $Y=3.63
+ $X2=0.925 $Y2=3.63
r49 16 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.925 $Y=3.59
+ $X2=0.925 $Y2=3.59
r50 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.205 $Y=3.59
+ $X2=0.205 $Y2=3.59
r51 13 16 16.0526 $w=9.48e-07 $l=1.25e-06 $layer=LI1_cond $X=0.565 $Y=2.34
+ $X2=0.565 $Y2=3.59
r52 10 37 0.385825 $w=3.7e-07 $l=1.005e-06 $layer=MET1_cond $X=2.4 $Y=3.63
+ $X2=3.405 $Y2=3.63
r53 10 27 0.24378 $w=3.7e-07 $l=6.35e-07 $layer=MET1_cond $X=2.4 $Y=3.63
+ $X2=1.765 $Y2=3.63
r54 10 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.485 $Y=3.59
+ $X2=2.485 $Y2=3.59
r55 3 36 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=3.585
+ $Y=2.215 $X2=3.725 $Y2=3.59
r56 3 33 300 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=2 $X=3.585
+ $Y=2.215 $X2=3.725 $Y2=2.385
r57 2 26 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.025
+ $Y=2.215 $X2=2.165 $Y2=3.59
r58 2 23 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.025
+ $Y=2.215 $X2=2.165 $Y2=2.34
r59 1 16 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.46
+ $Y=2.215 $X2=0.605 $Y2=3.59
r60 1 13 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.46
+ $Y=2.215 $X2=0.605 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_4%X 1 2 3 4 15 18 19 21 25 27 31 35 39 41 43 44
r64 43 44 24.051 $w=2.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.72 $Y2=1.665
r65 41 44 25.0531 $w=2.28e-07 $l=5e-07 $layer=LI1_cond $X=1.22 $Y=1.665 $X2=0.72
+ $Y2=1.665
r66 41 42 20.3333 $w=1.95e-07 $l=3.25e-07 $layer=LI1_cond $X=1.345 $Y=1.665
+ $X2=1.345 $Y2=1.99
r67 35 37 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=2.945 $Y=2.34
+ $X2=2.945 $Y2=3.59
r68 33 35 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.945 $Y=2.075
+ $X2=2.945 $Y2=2.34
r69 29 31 25.1233 $w=2.48e-07 $l=5.45e-07 $layer=LI1_cond $X=2.905 $Y=1.205
+ $X2=2.905 $Y2=0.66
r70 28 42 1.54022 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.47 $Y=1.99
+ $X2=1.345 $Y2=1.99
r71 27 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.78 $Y=1.99
+ $X2=2.945 $Y2=2.075
r72 27 28 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=2.78 $Y=1.99
+ $X2=1.47 $Y2=1.99
r73 26 39 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.47 $Y=1.29
+ $X2=1.345 $Y2=1.29
r74 25 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.78 $Y=1.29
+ $X2=2.905 $Y2=1.205
r75 25 26 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=2.78 $Y=1.29
+ $X2=1.47 $Y2=1.29
r76 21 23 57.6222 $w=2.48e-07 $l=1.25e-06 $layer=LI1_cond $X=1.345 $Y=2.34
+ $X2=1.345 $Y2=3.59
r77 19 42 4.77136 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.345 $Y=2.075
+ $X2=1.345 $Y2=1.99
r78 19 21 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.345 $Y=2.075
+ $X2=1.345 $Y2=2.34
r79 18 41 7.42769 $w=1.95e-07 $l=1.3351e-07 $layer=LI1_cond $X=1.305 $Y=1.55
+ $X2=1.345 $Y2=1.665
r80 17 39 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.305 $Y=1.375
+ $X2=1.345 $Y2=1.29
r81 17 18 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.305 $Y=1.375
+ $X2=1.305 $Y2=1.55
r82 13 39 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.345 $Y=1.205
+ $X2=1.345 $Y2=1.29
r83 13 15 25.1233 $w=2.48e-07 $l=5.45e-07 $layer=LI1_cond $X=1.345 $Y=1.205
+ $X2=1.345 $Y2=0.66
r84 4 37 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.805
+ $Y=2.215 $X2=2.945 $Y2=3.59
r85 4 35 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.805
+ $Y=2.215 $X2=2.945 $Y2=2.34
r86 3 23 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.245
+ $Y=2.215 $X2=1.385 $Y2=3.59
r87 3 21 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.245
+ $Y=2.215 $X2=1.385 $Y2=2.34
r88 2 31 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.805
+ $Y=0.535 $X2=2.945 $Y2=0.66
r89 1 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.245
+ $Y=0.535 $X2=1.385 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__BUF_4%VGND 1 2 3 10 13 22 31 35
r40 32 35 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.325 $Y=0.44
+ $X2=4.045 $Y2=0.44
r41 31 37 2.31158 $w=9.48e-07 $l=1.8e-07 $layer=LI1_cond $X=3.685 $Y=0.48
+ $X2=3.685 $Y2=0.66
r42 31 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.045 $Y=0.48
+ $X2=4.045 $Y2=0.48
r43 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.325 $Y=0.48
+ $X2=3.325 $Y2=0.48
r44 22 28 4.10947 $w=9.48e-07 $l=3.2e-07 $layer=LI1_cond $X=2.125 $Y=0.48
+ $X2=2.125 $Y2=0.8
r45 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.765 $Y=0.48
+ $X2=1.765 $Y2=0.48
r46 17 23 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=0.925 $Y=0.44
+ $X2=1.765 $Y2=0.44
r47 14 17 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.205 $Y=0.44
+ $X2=0.925 $Y2=0.44
r48 13 19 2.31158 $w=9.48e-07 $l=1.8e-07 $layer=LI1_cond $X=0.565 $Y=0.48
+ $X2=0.565 $Y2=0.66
r49 13 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.925 $Y=0.48
+ $X2=0.925 $Y2=0.48
r50 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.205 $Y=0.48
+ $X2=0.205 $Y2=0.48
r51 10 32 0.355112 $w=3.7e-07 $l=9.25e-07 $layer=MET1_cond $X=2.4 $Y=0.44
+ $X2=3.325 $Y2=0.44
r52 10 23 0.24378 $w=3.7e-07 $l=6.35e-07 $layer=MET1_cond $X=2.4 $Y=0.44
+ $X2=1.765 $Y2=0.44
r53 10 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.485 $Y=0.48
+ $X2=2.485 $Y2=0.48
r54 3 37 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.585
+ $Y=0.535 $X2=3.725 $Y2=0.66
r55 2 28 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.535 $X2=2.165 $Y2=0.8
r56 1 19 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.46
+ $Y=0.535 $X2=0.605 $Y2=0.66
.ends

