* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__decap_8 VGND VNB VPB VPWR
M1000 VPWR VGND VPWR VPB phv w=1e+06u l=1e+06u
+  ad=8.4e+11p pd=7.68e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nhv w=750000u l=1e+06u
+  ad=6.225e+11p pd=6.16e+06u as=0p ps=0u
M1002 VPWR VGND VPWR VPB phv w=1e+06u l=1e+06u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND VPWR VGND VNB nhv w=750000u l=1e+06u
+  ad=0p pd=0u as=0p ps=0u
.ends
