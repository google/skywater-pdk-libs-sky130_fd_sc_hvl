# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__mux4_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__mux4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.48000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A0
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.770000 1.550000 7.100000 2.520000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.400000 2.300000 4.730000 3.260000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.525000 1.515000 2.150000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 2.300000 3.845000 2.915000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 2.330000 2.155000 2.500000 ;
        RECT 0.565000 2.500000 0.895000 2.915000 ;
        RECT 1.905000 2.305000 2.155000 2.330000 ;
        RECT 1.905000 2.500000 2.155000 3.635000 ;
        RECT 1.905000 3.635000 3.060000 3.805000 ;
        RECT 2.685000 1.445000 5.420000 1.770000 ;
        RECT 2.685000 1.770000 2.855000 2.800000 ;
        RECT 2.685000 2.800000 3.060000 2.970000 ;
        RECT 2.890000 2.970000 3.060000 3.635000 ;
        RECT 4.925000 0.810000 5.420000 1.445000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.810000 1.920000 8.220000 2.885000 ;
        RECT 7.810000 2.885000 9.290000 2.915000 ;
        RECT 8.050000 2.915000 9.290000 3.055000 ;
        RECT 9.120000 1.315000 9.370000 1.985000 ;
        RECT 9.120000 1.985000 9.290000 2.885000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.120000 0.605000 12.370000 3.735000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.620000 0.365000  1.570000 0.995000 ;
        RECT  3.250000 0.365000  4.200000 0.915000 ;
        RECT  7.120000 0.365000  7.650000 0.995000 ;
        RECT 11.050000 0.365000 11.940000 1.415000 ;
      LAYER mcon ;
        RECT  0.650000 0.395000  0.820000 0.565000 ;
        RECT  1.010000 0.395000  1.180000 0.565000 ;
        RECT  1.370000 0.395000  1.540000 0.565000 ;
        RECT  3.280000 0.395000  3.450000 0.565000 ;
        RECT  3.640000 0.395000  3.810000 0.565000 ;
        RECT  4.000000 0.395000  4.170000 0.565000 ;
        RECT  7.120000 0.395000  7.290000 0.565000 ;
        RECT  7.480000 0.395000  7.650000 0.565000 ;
        RECT 11.050000 0.395000 11.220000 0.565000 ;
        RECT 11.410000 0.395000 11.580000 0.565000 ;
        RECT 11.770000 0.395000 11.940000 0.565000 ;
      LAYER met1 ;
        RECT 0.000000 0.255000 12.480000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 12.480000 0.085000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.115000 12.480000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 12.480000 4.155000 ;
      LAYER mcon ;
        RECT  0.155000 3.985000  0.325000 4.155000 ;
        RECT  0.635000 3.985000  0.805000 4.155000 ;
        RECT  1.115000 3.985000  1.285000 4.155000 ;
        RECT  1.595000 3.985000  1.765000 4.155000 ;
        RECT  2.075000 3.985000  2.245000 4.155000 ;
        RECT  2.555000 3.985000  2.725000 4.155000 ;
        RECT  3.035000 3.985000  3.205000 4.155000 ;
        RECT  3.515000 3.985000  3.685000 4.155000 ;
        RECT  3.995000 3.985000  4.165000 4.155000 ;
        RECT  4.475000 3.985000  4.645000 4.155000 ;
        RECT  4.955000 3.985000  5.125000 4.155000 ;
        RECT  5.435000 3.985000  5.605000 4.155000 ;
        RECT  5.915000 3.985000  6.085000 4.155000 ;
        RECT  6.395000 3.985000  6.565000 4.155000 ;
        RECT  6.875000 3.985000  7.045000 4.155000 ;
        RECT  7.355000 3.985000  7.525000 4.155000 ;
        RECT  7.835000 3.985000  8.005000 4.155000 ;
        RECT  8.315000 3.985000  8.485000 4.155000 ;
        RECT  8.795000 3.985000  8.965000 4.155000 ;
        RECT  9.275000 3.985000  9.445000 4.155000 ;
        RECT  9.755000 3.985000  9.925000 4.155000 ;
        RECT 10.235000 3.985000 10.405000 4.155000 ;
        RECT 10.715000 3.985000 10.885000 4.155000 ;
        RECT 11.195000 3.985000 11.365000 4.155000 ;
        RECT 11.675000 3.985000 11.845000 4.155000 ;
        RECT 12.155000 3.985000 12.325000 4.155000 ;
      LAYER met1 ;
        RECT 0.000000 3.955000 12.480000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.620000 3.095000  1.570000 3.705000 ;
        RECT  3.270000 3.095000  4.220000 3.705000 ;
        RECT  6.330000 3.095000  7.280000 3.705000 ;
        RECT 11.050000 2.175000 11.940000 3.755000 ;
      LAYER mcon ;
        RECT  0.650000 3.505000  0.820000 3.675000 ;
        RECT  1.010000 3.505000  1.180000 3.675000 ;
        RECT  1.370000 3.505000  1.540000 3.675000 ;
        RECT  3.300000 3.505000  3.470000 3.675000 ;
        RECT  3.660000 3.505000  3.830000 3.675000 ;
        RECT  4.020000 3.505000  4.190000 3.675000 ;
        RECT  6.360000 3.505000  6.530000 3.675000 ;
        RECT  6.720000 3.505000  6.890000 3.675000 ;
        RECT  7.080000 3.505000  7.250000 3.675000 ;
        RECT 11.050000 3.505000 11.220000 3.675000 ;
        RECT 11.410000 3.505000 11.580000 3.675000 ;
        RECT 11.770000 3.505000 11.940000 3.675000 ;
      LAYER met1 ;
        RECT 0.000000 3.445000 12.480000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.110000 0.515000  0.440000 1.175000 ;
      RECT  0.110000 1.175000  2.155000 1.345000 ;
      RECT  0.110000 1.345000  0.280000 3.115000 ;
      RECT  0.110000 3.115000  0.440000 3.575000 ;
      RECT  1.905000 1.345000  2.155000 2.035000 ;
      RECT  2.335000 0.495000  2.710000 1.095000 ;
      RECT  2.335000 1.095000  4.550000 1.265000 ;
      RECT  2.335000 1.265000  2.505000 3.175000 ;
      RECT  2.335000 3.175000  2.710000 3.455000 ;
      RECT  3.035000 1.950000  6.240000 2.120000 ;
      RECT  3.035000 2.120000  3.285000 2.620000 ;
      RECT  4.380000 0.265000  6.940000 0.435000 ;
      RECT  4.380000 0.435000  4.550000 1.095000 ;
      RECT  5.005000 2.120000  5.335000 2.915000 ;
      RECT  5.460000 3.095000  5.790000 3.595000 ;
      RECT  5.600000 0.615000  6.590000 0.915000 ;
      RECT  5.620000 2.745000  7.630000 2.915000 ;
      RECT  5.620000 2.915000  5.790000 3.095000 ;
      RECT  5.910000 1.095000  6.240000 1.950000 ;
      RECT  6.420000 0.915000  6.590000 2.745000 ;
      RECT  6.770000 0.435000  6.940000 1.175000 ;
      RECT  6.770000 1.175000  8.000000 1.345000 ;
      RECT  7.460000 1.570000  8.350000 1.740000 ;
      RECT  7.460000 1.740000  7.630000 2.745000 ;
      RECT  7.460000 2.915000  7.630000 3.115000 ;
      RECT  7.460000 3.115000  7.870000 3.535000 ;
      RECT  7.830000 0.265000  8.700000 0.435000 ;
      RECT  7.830000 0.435000  8.000000 1.175000 ;
      RECT  8.180000 0.615000  8.350000 1.570000 ;
      RECT  8.320000 3.235000  8.650000 3.635000 ;
      RECT  8.320000 3.635000 10.870000 3.805000 ;
      RECT  8.530000 0.435000  8.700000 0.965000 ;
      RECT  8.530000 0.965000  9.990000 1.035000 ;
      RECT  8.530000 1.035000  9.720000 1.135000 ;
      RECT  8.880000 0.265000 10.870000 0.435000 ;
      RECT  8.880000 0.435000  9.210000 0.785000 ;
      RECT  9.470000 3.115000  9.800000 3.455000 ;
      RECT  9.550000 0.615000  9.990000 0.965000 ;
      RECT  9.550000 1.135000  9.720000 3.115000 ;
      RECT  9.900000 2.115000 10.520000 2.655000 ;
      RECT  9.900000 2.655000 10.150000 2.915000 ;
      RECT 10.270000 0.915000 10.520000 2.115000 ;
      RECT 10.700000 0.435000 10.870000 1.595000 ;
      RECT 10.700000 1.595000 11.915000 1.925000 ;
      RECT 10.700000 1.925000 10.870000 3.635000 ;
  END
END sky130_fd_sc_hvl__mux4_1
