# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__or3_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__or3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.915000 1.080000 2.450000 1.390000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.910000 1.535000 3.260000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 1.080000 1.315000 1.390000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.460000 0.495000 3.715000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.530000 0.365000 1.385000 0.910000 ;
        RECT 2.620000 0.365000 3.290000 1.325000 ;
      LAYER mcon ;
        RECT 0.580000 0.395000 0.750000 0.565000 ;
        RECT 1.165000 0.395000 1.335000 0.565000 ;
        RECT 2.690000 0.395000 2.860000 0.565000 ;
        RECT 3.050000 0.395000 3.220000 0.565000 ;
      LAYER met1 ;
        RECT 0.000000 0.255000 3.840000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.840000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 3.840000 4.155000 ;
      LAYER mcon ;
        RECT 0.155000 3.985000 0.325000 4.155000 ;
        RECT 0.635000 3.985000 0.805000 4.155000 ;
        RECT 1.115000 3.985000 1.285000 4.155000 ;
        RECT 1.595000 3.985000 1.765000 4.155000 ;
        RECT 2.075000 3.985000 2.245000 4.155000 ;
        RECT 2.555000 3.985000 2.725000 4.155000 ;
        RECT 3.035000 3.985000 3.205000 4.155000 ;
        RECT 3.515000 3.985000 3.685000 4.155000 ;
      LAYER met1 ;
        RECT 0.000000 3.955000 3.840000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.620000 3.430000 3.280000 3.755000 ;
        RECT 1.705000 2.175000 3.280000 3.430000 ;
      LAYER mcon ;
        RECT 1.670000 3.505000 1.840000 3.675000 ;
        RECT 2.030000 3.505000 2.200000 3.675000 ;
        RECT 2.390000 3.505000 2.560000 3.675000 ;
        RECT 2.750000 3.505000 2.920000 3.675000 ;
        RECT 3.110000 3.505000 3.280000 3.675000 ;
      LAYER met1 ;
        RECT 0.000000 3.445000 3.840000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.145000 0.495000 0.360000 1.560000 ;
      RECT 0.145000 1.560000 3.255000 1.730000 ;
      RECT 0.145000 1.730000 0.395000 2.780000 ;
      RECT 1.565000 0.495000 1.965000 0.910000 ;
      RECT 1.565000 0.910000 1.735000 1.560000 ;
      RECT 2.925000 1.730000 3.255000 1.935000 ;
  END
END sky130_fd_sc_hvl__or3_1
