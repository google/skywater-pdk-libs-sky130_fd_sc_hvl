# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__dfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__dfrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.36000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.415000 0.810000 3.745000 2.105000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.611250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.900000 0.665000 15.235000 3.735000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  2.695000 1.620000  3.235000 2.490000 ;
        RECT  3.065000 0.460000  6.010000 0.630000 ;
        RECT  3.065000 0.630000  3.235000 1.620000 ;
        RECT  5.840000 0.630000  6.010000 1.125000 ;
        RECT  5.840000 1.125000  8.460000 1.295000 ;
        RECT  6.605000 1.825000  8.460000 1.995000 ;
        RECT  8.290000 0.265000 10.950000 0.435000 ;
        RECT  8.290000 0.435000  8.460000 1.125000 ;
        RECT  8.290000 1.295000  8.460000 1.825000 ;
        RECT 10.780000 0.435000 10.950000 1.095000 ;
        RECT 10.780000 1.095000 11.785000 1.265000 ;
        RECT 11.455000 1.265000 11.785000 1.655000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.175000 0.890000 2.150000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.560000 0.365000  1.510000 0.995000 ;
        RECT  2.200000 0.365000  2.790000 1.245000 ;
        RECT  7.160000 0.365000  8.110000 0.945000 ;
        RECT 11.130000 0.365000 12.080000 0.915000 ;
        RECT 13.735000 0.365000 14.685000 1.495000 ;
      LAYER mcon ;
        RECT  0.590000 0.395000  0.760000 0.565000 ;
        RECT  0.950000 0.395000  1.120000 0.565000 ;
        RECT  1.310000 0.395000  1.480000 0.565000 ;
        RECT  2.230000 0.395000  2.400000 0.565000 ;
        RECT  2.590000 0.395000  2.760000 0.565000 ;
        RECT  7.190000 0.395000  7.360000 0.565000 ;
        RECT  7.550000 0.395000  7.720000 0.565000 ;
        RECT  7.910000 0.395000  8.080000 0.565000 ;
        RECT 11.160000 0.395000 11.330000 0.565000 ;
        RECT 11.520000 0.395000 11.690000 0.565000 ;
        RECT 11.880000 0.395000 12.050000 0.565000 ;
        RECT 13.765000 0.395000 13.935000 0.565000 ;
        RECT 14.125000 0.395000 14.295000 0.565000 ;
        RECT 14.485000 0.395000 14.655000 0.565000 ;
      LAYER met1 ;
        RECT 0.000000 0.255000 15.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 15.360000 0.085000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.115000 15.360000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 15.360000 4.155000 ;
      LAYER mcon ;
        RECT  0.155000 3.985000  0.325000 4.155000 ;
        RECT  0.635000 3.985000  0.805000 4.155000 ;
        RECT  1.115000 3.985000  1.285000 4.155000 ;
        RECT  1.595000 3.985000  1.765000 4.155000 ;
        RECT  2.075000 3.985000  2.245000 4.155000 ;
        RECT  2.555000 3.985000  2.725000 4.155000 ;
        RECT  3.035000 3.985000  3.205000 4.155000 ;
        RECT  3.515000 3.985000  3.685000 4.155000 ;
        RECT  3.995000 3.985000  4.165000 4.155000 ;
        RECT  4.475000 3.985000  4.645000 4.155000 ;
        RECT  4.955000 3.985000  5.125000 4.155000 ;
        RECT  5.435000 3.985000  5.605000 4.155000 ;
        RECT  5.915000 3.985000  6.085000 4.155000 ;
        RECT  6.395000 3.985000  6.565000 4.155000 ;
        RECT  6.875000 3.985000  7.045000 4.155000 ;
        RECT  7.355000 3.985000  7.525000 4.155000 ;
        RECT  7.835000 3.985000  8.005000 4.155000 ;
        RECT  8.315000 3.985000  8.485000 4.155000 ;
        RECT  8.795000 3.985000  8.965000 4.155000 ;
        RECT  9.275000 3.985000  9.445000 4.155000 ;
        RECT  9.755000 3.985000  9.925000 4.155000 ;
        RECT 10.235000 3.985000 10.405000 4.155000 ;
        RECT 10.715000 3.985000 10.885000 4.155000 ;
        RECT 11.195000 3.985000 11.365000 4.155000 ;
        RECT 11.675000 3.985000 11.845000 4.155000 ;
        RECT 12.155000 3.985000 12.325000 4.155000 ;
        RECT 12.635000 3.985000 12.805000 4.155000 ;
        RECT 13.115000 3.985000 13.285000 4.155000 ;
        RECT 13.595000 3.985000 13.765000 4.155000 ;
        RECT 14.075000 3.985000 14.245000 4.155000 ;
        RECT 14.555000 3.985000 14.725000 4.155000 ;
        RECT 15.035000 3.985000 15.205000 4.155000 ;
      LAYER met1 ;
        RECT 0.000000 3.955000 15.360000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.630000 2.725000  1.220000 3.705000 ;
        RECT  3.020000 3.370000  3.350000 3.705000 ;
        RECT  5.450000 3.225000  6.400000 3.705000 ;
        RECT  7.790000 3.455000  8.740000 3.755000 ;
        RECT 10.485000 2.675000 11.435000 3.705000 ;
        RECT 12.270000 2.885000 13.165000 3.705000 ;
        RECT 13.775000 2.195000 14.720000 3.735000 ;
      LAYER mcon ;
        RECT  0.660000 3.505000  0.830000 3.675000 ;
        RECT  1.020000 3.505000  1.190000 3.675000 ;
        RECT  3.050000 3.505000  3.220000 3.675000 ;
        RECT  5.480000 3.505000  5.650000 3.675000 ;
        RECT  5.840000 3.505000  6.010000 3.675000 ;
        RECT  6.200000 3.505000  6.370000 3.675000 ;
        RECT  7.820000 3.505000  7.990000 3.675000 ;
        RECT  8.180000 3.505000  8.350000 3.675000 ;
        RECT  8.540000 3.505000  8.710000 3.675000 ;
        RECT 10.515000 3.505000 10.685000 3.675000 ;
        RECT 10.875000 3.505000 11.045000 3.675000 ;
        RECT 11.235000 3.505000 11.405000 3.675000 ;
        RECT 12.270000 3.505000 12.440000 3.675000 ;
        RECT 12.630000 3.505000 12.800000 3.675000 ;
        RECT 12.990000 3.505000 13.160000 3.675000 ;
        RECT 13.800000 3.505000 13.970000 3.675000 ;
        RECT 14.160000 3.505000 14.330000 3.675000 ;
        RECT 14.520000 3.505000 14.690000 3.675000 ;
      LAYER met1 ;
        RECT 0.000000 3.445000 15.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.110000 0.495000  0.380000 2.355000 ;
      RECT  0.110000 2.355000  1.570000 2.525000 ;
      RECT  0.110000 2.525000  0.440000 3.455000 ;
      RECT  1.240000 1.855000  1.570000 2.355000 ;
      RECT  1.400000 2.525000  1.570000 3.635000 ;
      RECT  1.400000 3.635000  2.840000 3.805000 ;
      RECT  1.690000 0.495000  2.020000 0.995000 ;
      RECT  1.750000 0.995000  2.020000 1.920000 ;
      RECT  1.750000 1.920000  2.275000 2.150000 ;
      RECT  1.750000 2.150000  2.000000 3.455000 ;
      RECT  2.240000 2.670000  4.050000 2.840000 ;
      RECT  2.240000 2.840000  2.490000 3.455000 ;
      RECT  2.670000 3.020000  3.700000 3.190000 ;
      RECT  2.670000 3.190000  2.840000 3.635000 ;
      RECT  3.530000 3.190000  3.700000 3.635000 ;
      RECT  3.530000 3.635000  5.270000 3.805000 ;
      RECT  3.880000 2.320000  4.100000 2.490000 ;
      RECT  3.880000 2.490000  4.050000 2.670000 ;
      RECT  3.880000 2.840000  4.050000 3.455000 ;
      RECT  3.930000 0.825000  4.200000 1.325000 ;
      RECT  3.930000 1.325000  4.100000 2.320000 ;
      RECT  4.230000 2.670000  4.450000 3.000000 ;
      RECT  4.280000 1.920000  5.305000 2.150000 ;
      RECT  4.280000 2.150000  4.450000 2.670000 ;
      RECT  4.580000 3.200000  4.910000 3.455000 ;
      RECT  4.630000 2.330000  5.660000 2.500000 ;
      RECT  4.630000 2.500000  4.800000 3.200000 ;
      RECT  4.650000 0.825000  4.980000 1.075000 ;
      RECT  4.650000 1.075000  5.660000 1.245000 ;
      RECT  4.975000 1.425000  5.305000 1.920000 ;
      RECT  4.980000 2.680000  5.310000 2.875000 ;
      RECT  4.980000 2.875000  6.750000 3.000000 ;
      RECT  5.100000 3.000000  6.750000 3.045000 ;
      RECT  5.100000 3.045000  5.270000 3.635000 ;
      RECT  5.490000 1.245000  5.660000 1.475000 ;
      RECT  5.490000 1.475000  8.110000 1.645000 ;
      RECT  5.490000 1.645000  5.660000 2.330000 ;
      RECT  5.490000 2.500000  5.660000 2.525000 ;
      RECT  5.490000 2.525000  7.260000 2.695000 ;
      RECT  5.840000 1.825000  6.170000 2.175000 ;
      RECT  5.840000 2.175000  8.900000 2.345000 ;
      RECT  6.580000 3.045000  6.750000 3.635000 ;
      RECT  6.580000 3.635000  7.610000 3.805000 ;
      RECT  6.930000 2.695000  7.260000 3.455000 ;
      RECT  7.440000 3.105000  9.250000 3.275000 ;
      RECT  7.440000 3.275000  7.610000 3.635000 ;
      RECT  8.570000 2.345000  8.900000 2.925000 ;
      RECT  8.640000 0.615000  8.970000 1.325000 ;
      RECT  8.640000 1.325000  8.900000 2.175000 ;
      RECT  9.080000 1.585000 10.250000 1.755000 ;
      RECT  9.080000 1.755000  9.250000 3.105000 ;
      RECT  9.430000 0.615000 10.600000 0.785000 ;
      RECT  9.430000 0.785000  9.760000 1.325000 ;
      RECT  9.430000 2.675000 10.305000 2.845000 ;
      RECT  9.430000 2.845000  9.680000 3.755000 ;
      RECT  9.625000 1.935000  9.955000 2.435000 ;
      RECT  9.965000 1.085000 10.250000 1.585000 ;
      RECT 10.135000 2.185000 12.495000 2.355000 ;
      RECT 10.135000 2.355000 10.305000 2.675000 ;
      RECT 10.430000 0.785000 10.600000 2.185000 ;
      RECT 10.805000 1.445000 11.135000 1.835000 ;
      RECT 10.805000 1.835000 12.845000 2.005000 ;
      RECT 11.840000 2.535000 12.845000 2.705000 ;
      RECT 11.840000 2.705000 12.090000 3.175000 ;
      RECT 12.620000 0.495000 12.950000 0.995000 ;
      RECT 12.620000 0.995000 12.845000 1.835000 ;
      RECT 12.675000 2.005000 12.845000 2.535000 ;
      RECT 13.225000 0.995000 13.555000 1.495000 ;
      RECT 13.345000 1.495000 13.555000 1.675000 ;
      RECT 13.345000 1.675000 14.720000 2.005000 ;
      RECT 13.345000 2.005000 13.595000 3.005000 ;
    LAYER mcon ;
      RECT 2.075000 1.950000 2.245000 2.120000 ;
      RECT 4.475000 1.950000 4.645000 2.120000 ;
      RECT 9.755000 1.950000 9.925000 2.120000 ;
    LAYER met1 ;
      RECT 2.015000 1.920000 2.305000 1.965000 ;
      RECT 2.015000 1.965000 9.985000 2.105000 ;
      RECT 2.015000 2.105000 2.305000 2.150000 ;
      RECT 4.415000 1.920000 4.705000 1.965000 ;
      RECT 4.415000 2.105000 4.705000 2.150000 ;
      RECT 9.695000 1.920000 9.985000 1.965000 ;
      RECT 9.695000 2.105000 9.985000 2.150000 ;
  END
END sky130_fd_sc_hvl__dfrtp_1
