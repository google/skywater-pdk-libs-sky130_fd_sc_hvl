# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
SITE unithvdbl
    SYMMETRY y  ;
    CLASS CORE  ;
    SIZE  0.480 BY 8.140 ;
END unithvdbl
MACRO sky130_fd_sc_hvl__a22o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.505000 4.645000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.825000 1.505000 5.155000 1.750000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 0.810000 3.205000 1.750000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.775000 2.320000 3.260000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.495000 0.380000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 5.280000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 5.280000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 5.280000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 5.280000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.985000 5.280000 4.155000 ;
      RECT 0.550000  0.365000 2.260000 1.245000 ;
      RECT 0.560000  2.175000 1.460000 3.755000 ;
      RECT 0.585000  1.425000 2.855000 1.595000 ;
      RECT 0.585000  1.595000 0.915000 1.755000 ;
      RECT 1.640000  2.175000 1.810000 3.635000 ;
      RECT 1.640000  3.635000 3.530000 3.805000 ;
      RECT 2.500000  1.595000 2.830000 3.455000 ;
      RECT 2.685000  0.460000 3.635000 0.630000 ;
      RECT 2.685000  0.630000 2.855000 1.425000 ;
      RECT 3.280000  1.930000 5.170000 2.100000 ;
      RECT 3.280000  2.100000 3.530000 3.635000 ;
      RECT 3.385000  0.630000 3.635000 1.325000 ;
      RECT 3.710000  2.280000 4.660000 3.755000 ;
      RECT 3.815000  0.365000 5.125000 1.325000 ;
      RECT 4.840000  2.100000 5.170000 3.735000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.565000  3.505000 0.735000 3.675000 ;
      RECT 0.600000  0.395000 0.770000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.925000  3.505000 1.095000 3.675000 ;
      RECT 0.960000  0.395000 1.130000 0.565000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.285000  3.505000 1.455000 3.675000 ;
      RECT 1.320000  0.395000 1.490000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.680000  0.395000 1.850000 0.565000 ;
      RECT 2.040000  0.395000 2.210000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.740000  3.505000 3.910000 3.675000 ;
      RECT 3.845000  0.395000 4.015000 0.565000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.100000  3.505000 4.270000 3.675000 ;
      RECT 4.205000  0.395000 4.375000 0.565000 ;
      RECT 4.460000  3.505000 4.630000 3.675000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.565000  0.395000 4.735000 0.565000 ;
      RECT 4.925000  0.395000 5.095000 0.565000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
  END
END sky130_fd_sc_hvl__a22o_1
