* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 a_2310_107# a_938_107# a_2123_543# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.344e+11p ps=1.48e+06u
M1001 VGND a_2352_81# a_2310_107# VNB nhv w=420000u l=500000u
+  ad=1.05015e+12p pd=1.074e+07u as=0p ps=0u
M1002 a_2352_81# a_2123_543# VGND VNB nhv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
M1003 VPWR SCE a_30_593# VPB phv w=420000u l=500000u
+  ad=1.6012e+12p pd=1.475e+07u as=1.197e+11p ps=1.41e+06u
M1004 VPWR a_2352_81# a_2302_543# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=1.05e+11p ps=1.34e+06u
M1005 a_2352_81# a_2123_543# VPWR VPB phv w=1e+06u l=500000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1006 a_641_593# a_30_593# a_484_107# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=2.289e+11p ps=2.77e+06u
M1007 VPWR SCD a_641_593# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_938_107# CLK VGND VNB nhv w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1009 a_938_107# CLK VPWR VPB phv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
M1010 VPWR a_2352_81# Q VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=3.975e+11p ps=3.53e+06u
M1011 VGND SCE a_30_593# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1012 VGND a_2352_81# Q VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u
M1013 a_1688_81# a_1490_107# VGND VNB nhv w=750000u l=500000u
+  ad=2.5995e+11p pd=2.29e+06u as=0p ps=0u
M1014 a_343_593# SCE VPWR VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1015 a_640_107# SCE a_484_107# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=2.709e+11p ps=2.97e+06u
M1016 a_484_107# D a_343_593# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1688_81# a_1490_107# VPWR VPB phv w=1e+06u l=500000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1018 VGND SCD a_640_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1204_107# a_938_107# VGND VNB nhv w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1020 a_1204_107# a_938_107# VPWR VPB phv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
M1021 a_1646_107# a_1204_107# a_1490_107# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1022 VGND a_1688_81# a_1646_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_2302_543# a_1204_107# a_2123_543# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=3.312e+11p ps=2.79e+06u
M1024 a_1646_543# a_938_107# a_1490_107# VPB phv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1025 a_342_107# D VGND VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1026 VPWR a_1688_81# a_1646_543# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_484_107# a_30_593# a_342_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1490_107# a_938_107# a_484_107# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_2123_543# a_1204_107# a_1688_81# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1490_107# a_1204_107# a_484_107# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_2123_543# a_938_107# a_1688_81# VPB phv w=1e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
