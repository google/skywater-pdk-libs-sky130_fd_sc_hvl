* File: sky130_fd_sc_hvl__mux2_1.pxi.spice
* Created: Fri Aug 28 09:37:42 2020
* 
x_PM_SKY130_FD_SC_HVL__MUX2_1%VNB N_VNB_M1009_b VNB N_VNB_c_5_p VNB
+ PM_SKY130_FD_SC_HVL__MUX2_1%VNB
x_PM_SKY130_FD_SC_HVL__MUX2_1%VPB N_VPB_M1002_b VPB N_VPB_c_43_p VPB
+ PM_SKY130_FD_SC_HVL__MUX2_1%VPB
x_PM_SKY130_FD_SC_HVL__MUX2_1%A_94_81# N_A_94_81#_M1006_d N_A_94_81#_M1007_d
+ N_A_94_81#_c_72_n N_A_94_81#_c_73_n N_A_94_81#_c_103_p N_A_94_81#_c_90_p
+ N_A_94_81#_c_80_n N_A_94_81#_c_97_p N_A_94_81#_c_88_p N_A_94_81#_c_74_n
+ N_A_94_81#_c_75_n N_A_94_81#_c_81_n N_A_94_81#_M1009_g N_A_94_81#_M1002_g
+ PM_SKY130_FD_SC_HVL__MUX2_1%A_94_81#
x_PM_SKY130_FD_SC_HVL__MUX2_1%S N_S_c_152_n N_S_c_153_n N_S_c_154_n N_S_c_155_n
+ N_S_c_156_n N_S_c_176_p S S N_S_M1001_g N_S_M1004_g N_S_M1008_g N_S_M1010_g
+ PM_SKY130_FD_SC_HVL__MUX2_1%S
x_PM_SKY130_FD_SC_HVL__MUX2_1%A0 N_A0_M1007_g N_A0_c_222_n N_A0_c_223_n
+ N_A0_c_229_n N_A0_c_224_n A0 A0 N_A0_M1011_g N_A0_c_230_n
+ PM_SKY130_FD_SC_HVL__MUX2_1%A0
x_PM_SKY130_FD_SC_HVL__MUX2_1%A1 N_A1_c_283_n N_A1_M1006_g N_A1_c_286_n A1
+ N_A1_c_288_n N_A1_M1000_g PM_SKY130_FD_SC_HVL__MUX2_1%A1
x_PM_SKY130_FD_SC_HVL__MUX2_1%A_713_81# N_A_713_81#_M1008_d N_A_713_81#_M1010_d
+ N_A_713_81#_M1003_g N_A_713_81#_c_338_n N_A_713_81#_M1005_g
+ N_A_713_81#_c_339_n N_A_713_81#_c_340_n N_A_713_81#_c_342_n
+ N_A_713_81#_c_360_n N_A_713_81#_c_343_n PM_SKY130_FD_SC_HVL__MUX2_1%A_713_81#
x_PM_SKY130_FD_SC_HVL__MUX2_1%X N_X_M1009_s N_X_M1002_s X X X X X X X
+ N_X_c_383_n X PM_SKY130_FD_SC_HVL__MUX2_1%X
x_PM_SKY130_FD_SC_HVL__MUX2_1%VPWR N_VPWR_M1002_d N_VPWR_M1005_d VPWR
+ N_VPWR_c_397_n N_VPWR_c_400_n N_VPWR_c_403_n PM_SKY130_FD_SC_HVL__MUX2_1%VPWR
x_PM_SKY130_FD_SC_HVL__MUX2_1%VGND N_VGND_M1009_d N_VGND_M1003_d VGND
+ N_VGND_c_431_n N_VGND_c_433_n N_VGND_c_435_n PM_SKY130_FD_SC_HVL__MUX2_1%VGND
cc_1 N_VNB_M1009_b N_A_94_81#_c_72_n 0.0158688f $X=-0.33 $Y=-0.265 $X2=1.945
+ $Y2=1.44
cc_2 N_VNB_M1009_b N_A_94_81#_c_73_n 0.00549993f $X=-0.33 $Y=-0.265 $X2=2.03
+ $Y2=2.415
cc_3 N_VNB_M1009_b N_A_94_81#_c_74_n 0.00124242f $X=-0.33 $Y=-0.265 $X2=2.03
+ $Y2=1.44
cc_4 N_VNB_M1009_b N_A_94_81#_c_75_n 0.0148882f $X=-0.33 $Y=-0.265 $X2=2.715
+ $Y2=0.745
cc_5 N_VNB_c_5_p N_A_94_81#_c_75_n 0.00157394f $X=0.24 $Y=0 $X2=2.715 $Y2=0.745
cc_6 N_VNB_M1009_b N_A_94_81#_M1009_g 0.092832f $X=-0.33 $Y=-0.265 $X2=0.72
+ $Y2=0.91
cc_7 N_VNB_c_5_p N_A_94_81#_M1009_g 5.86481e-19 $X=0.24 $Y=0 $X2=0.72 $Y2=0.91
cc_8 N_VNB_M1009_b N_S_M1001_g 0.110438f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_M1009_b N_S_M1008_g 0.120198f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_10 N_VNB_c_5_p N_S_M1008_g 5.81826e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_11 N_VNB_M1009_b N_A0_c_222_n 0.00487441f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_12 N_VNB_M1009_b N_A0_c_223_n 0.004174f $X=-0.33 $Y=-0.265 $X2=1.945 $Y2=1.44
cc_13 N_VNB_M1009_b N_A0_c_224_n 0.00286374f $X=-0.33 $Y=-0.265 $X2=2.03
+ $Y2=2.415
cc_14 N_VNB_M1009_b A0 0.00381372f $X=-0.33 $Y=-0.265 $X2=2.115 $Y2=1.44
cc_15 N_VNB_M1009_b N_A0_M1011_g 0.0744716f $X=-0.33 $Y=-0.265 $X2=2.47
+ $Y2=1.355
cc_16 N_VNB_c_5_p N_A0_M1011_g 9.54195e-19 $X=0.24 $Y=0 $X2=2.47 $Y2=1.355
cc_17 N_VNB_M1009_b N_A1_c_283_n 0.0679619f $X=-0.33 $Y=-0.265 $X2=2.575
+ $Y2=0.535
cc_18 N_VNB_M1009_b N_A1_M1006_g 0.0445944f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_19 N_VNB_c_5_p N_A1_M1006_g 0.00172686f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_20 N_VNB_M1009_b N_A1_c_286_n 0.0325204f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_21 N_VNB_M1009_b A1 0.00392158f $X=-0.33 $Y=-0.265 $X2=2.03 $Y2=1.525
cc_22 N_VNB_M1009_b N_A1_c_288_n 0.0118122f $X=-0.33 $Y=-0.265 $X2=2.115
+ $Y2=1.44
cc_23 N_VNB_M1009_b N_A_713_81#_M1003_g 0.038243f $X=-0.33 $Y=-0.265 $X2=2.03
+ $Y2=1.525
cc_24 N_VNB_M1009_b N_A_713_81#_c_338_n 0.0769514f $X=-0.33 $Y=-0.265 $X2=2.385
+ $Y2=1.44
cc_25 N_VNB_M1009_b N_A_713_81#_c_339_n 0.0117525f $X=-0.33 $Y=-0.265 $X2=0.785
+ $Y2=1.44
cc_26 N_VNB_M1009_b N_A_713_81#_c_340_n 0.0305191f $X=-0.33 $Y=-0.265 $X2=0.785
+ $Y2=1.58
cc_27 N_VNB_c_5_p N_A_713_81#_c_340_n 5.81195e-19 $X=0.24 $Y=0 $X2=0.785
+ $Y2=1.58
cc_28 N_VNB_M1009_b N_A_713_81#_c_342_n 0.0314483f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_29 N_VNB_M1009_b N_A_713_81#_c_343_n 0.00770964f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_30 N_VNB_M1009_b N_X_c_383_n 0.0703834f $X=-0.33 $Y=-0.265 $X2=2.47 $Y2=0.705
cc_31 N_VNB_c_5_p N_X_c_383_n 6.74937e-19 $X=0.24 $Y=0 $X2=2.47 $Y2=0.705
cc_32 N_VNB_M1009_b N_VGND_c_431_n 0.0823021f $X=-0.33 $Y=-0.265 $X2=2.03
+ $Y2=2.415
cc_33 N_VNB_c_5_p N_VGND_c_431_n 0.00456362f $X=0.24 $Y=0 $X2=2.03 $Y2=2.415
cc_34 N_VNB_M1009_b N_VGND_c_433_n 0.0810147f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_35 N_VNB_c_5_p N_VGND_c_433_n 0.00472015f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_36 N_VNB_M1009_b N_VGND_c_435_n 0.0896289f $X=-0.33 $Y=-0.265 $X2=2.715
+ $Y2=0.705
cc_37 N_VNB_c_5_p N_VGND_c_435_n 0.564575f $X=0.24 $Y=0 $X2=2.715 $Y2=0.705
cc_38 N_VPB_M1002_b N_A_94_81#_c_73_n 0.00387885f $X=-0.33 $Y=1.885 $X2=2.03
+ $Y2=2.415
cc_39 N_VPB_M1002_b N_A_94_81#_c_80_n 2.35532e-19 $X=-0.33 $Y=1.885 $X2=2.115
+ $Y2=2.5
cc_40 N_VPB_M1002_b N_A_94_81#_c_81_n 0.00536064f $X=-0.33 $Y=1.885 $X2=2.715
+ $Y2=2.5
cc_41 N_VPB_M1002_b N_A_94_81#_M1009_g 0.063533f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=0.91
cc_42 VPB N_A_94_81#_M1009_g 0.00970178f $X=0 $Y=3.955 $X2=0.72 $Y2=0.91
cc_43 N_VPB_c_43_p N_A_94_81#_M1009_g 0.0158814f $X=5.04 $Y=4.07 $X2=0.72
+ $Y2=0.91
cc_44 N_VPB_M1002_b N_S_c_152_n 0.00396206f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_45 N_VPB_M1002_b N_S_c_153_n 0.0397993f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_46 N_VPB_M1002_b N_S_c_154_n 0.00656678f $X=-0.33 $Y=1.885 $X2=1.945 $Y2=1.44
cc_47 N_VPB_M1002_b N_S_c_155_n 0.00389099f $X=-0.33 $Y=1.885 $X2=2.03 $Y2=1.525
cc_48 N_VPB_M1002_b N_S_c_156_n 0.0153477f $X=-0.33 $Y=1.885 $X2=2.03 $Y2=2.415
cc_49 N_VPB_M1002_b N_S_M1001_g 0.0808021f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_50 N_VPB_M1002_b N_S_M1008_g 0.0837942f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_51 N_VPB_M1002_b N_A0_c_223_n 0.00381078f $X=-0.33 $Y=1.885 $X2=1.945
+ $Y2=1.44
cc_52 N_VPB_M1002_b N_A0_c_229_n 0.0423288f $X=-0.33 $Y=1.885 $X2=0.95 $Y2=1.44
cc_53 N_VPB_M1002_b N_A0_c_230_n 0.0327f $X=-0.33 $Y=1.885 $X2=2.47 $Y2=0.705
cc_54 N_VPB_M1002_b A1 0.00199489f $X=-0.33 $Y=1.885 $X2=2.03 $Y2=1.525
cc_55 N_VPB_M1002_b N_A1_c_288_n 0.0753104f $X=-0.33 $Y=1.885 $X2=2.115 $Y2=1.44
cc_56 N_VPB_M1002_b N_A_713_81#_c_338_n 0.0384082f $X=-0.33 $Y=1.885 $X2=2.385
+ $Y2=1.44
cc_57 N_VPB_M1002_b N_A_713_81#_M1005_g 0.0357236f $X=-0.33 $Y=1.885 $X2=2.55
+ $Y2=2.5
cc_58 N_VPB_M1002_b N_A_713_81#_c_342_n 0.0520845f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_59 N_VPB_M1002_b X 0.0704487f $X=-0.33 $Y=1.885 $X2=2.03 $Y2=2.415
cc_60 VPB X 0.00116953f $X=0 $Y=3.955 $X2=2.03 $Y2=2.415
cc_61 N_VPB_c_43_p X 0.019351f $X=5.04 $Y=4.07 $X2=2.03 $Y2=2.415
cc_62 N_VPB_M1002_b N_X_c_383_n 0.00204542f $X=-0.33 $Y=1.885 $X2=2.47 $Y2=0.705
cc_63 N_VPB_M1002_b N_VPWR_c_397_n 0.00718665f $X=-0.33 $Y=1.885 $X2=2.03
+ $Y2=2.415
cc_64 VPB N_VPWR_c_397_n 0.00228138f $X=0 $Y=3.955 $X2=2.03 $Y2=2.415
cc_65 N_VPB_c_43_p N_VPWR_c_397_n 0.0293794f $X=5.04 $Y=4.07 $X2=2.03 $Y2=2.415
cc_66 N_VPB_M1002_b N_VPWR_c_400_n 0.0672796f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_400_n 0.0037122f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_68 N_VPB_c_43_p N_VPWR_c_400_n 0.0565652f $X=5.04 $Y=4.07 $X2=0 $Y2=0
cc_69 N_VPB_M1002_b N_VPWR_c_403_n 0.110804f $X=-0.33 $Y=1.885 $X2=2.47
+ $Y2=0.705
cc_70 VPB N_VPWR_c_403_n 0.563986f $X=0 $Y=3.955 $X2=2.47 $Y2=0.705
cc_71 N_VPB_c_43_p N_VPWR_c_403_n 0.0313483f $X=5.04 $Y=4.07 $X2=2.47 $Y2=0.705
cc_72 N_A_94_81#_c_72_n N_S_c_152_n 0.0238596f $X=1.945 $Y=1.44 $X2=0 $Y2=0
cc_73 N_A_94_81#_c_73_n N_S_c_152_n 0.0510684f $X=2.03 $Y=2.415 $X2=0 $Y2=0
cc_74 N_A_94_81#_c_80_n N_S_c_152_n 0.0133752f $X=2.115 $Y=2.5 $X2=0 $Y2=0
cc_75 N_A_94_81#_c_88_p N_S_c_152_n 0.00127882f $X=0.785 $Y=1.44 $X2=0 $Y2=0
cc_76 N_A_94_81#_M1009_g N_S_c_152_n 0.0029706f $X=0.72 $Y=0.91 $X2=0 $Y2=0
cc_77 N_A_94_81#_c_90_p N_S_c_153_n 0.0135765f $X=2.55 $Y=2.5 $X2=0 $Y2=0
cc_78 N_A_94_81#_c_80_n N_S_c_153_n 0.00510433f $X=2.115 $Y=2.5 $X2=0 $Y2=0
cc_79 N_A_94_81#_c_81_n N_S_c_153_n 0.0247177f $X=2.715 $Y=2.5 $X2=0 $Y2=0
cc_80 N_A_94_81#_c_81_n N_S_c_155_n 0.0341066f $X=2.715 $Y=2.5 $X2=0 $Y2=0
cc_81 N_A_94_81#_c_72_n N_S_M1001_g 0.0312875f $X=1.945 $Y=1.44 $X2=0 $Y2=0
cc_82 N_A_94_81#_c_73_n N_S_M1001_g 0.0134098f $X=2.03 $Y=2.415 $X2=0 $Y2=0
cc_83 N_A_94_81#_c_80_n N_S_M1001_g 0.00132298f $X=2.115 $Y=2.5 $X2=0 $Y2=0
cc_84 N_A_94_81#_c_97_p N_S_M1001_g 8.46355e-19 $X=2.47 $Y=1.355 $X2=0 $Y2=0
cc_85 N_A_94_81#_c_88_p N_S_M1001_g 0.00144981f $X=0.785 $Y=1.44 $X2=0 $Y2=0
cc_86 N_A_94_81#_c_75_n N_S_M1001_g 2.38138e-19 $X=2.715 $Y=0.745 $X2=0 $Y2=0
cc_87 N_A_94_81#_c_81_n N_S_M1001_g 0.00101042f $X=2.715 $Y=2.5 $X2=0 $Y2=0
cc_88 N_A_94_81#_M1009_g N_S_M1001_g 0.060098f $X=0.72 $Y=0.91 $X2=0 $Y2=0
cc_89 N_A_94_81#_c_73_n N_A0_c_222_n 0.00701237f $X=2.03 $Y=2.415 $X2=-0.33
+ $Y2=-0.265
cc_90 N_A_94_81#_c_103_p N_A0_c_222_n 0.0102924f $X=2.385 $Y=1.44 $X2=-0.33
+ $Y2=-0.265
cc_91 N_A_94_81#_c_73_n N_A0_c_223_n 0.032938f $X=2.03 $Y=2.415 $X2=0 $Y2=0
cc_92 N_A_94_81#_c_103_p N_A0_c_223_n 0.0155862f $X=2.385 $Y=1.44 $X2=0 $Y2=0
cc_93 N_A_94_81#_c_90_p N_A0_c_223_n 0.0179247f $X=2.55 $Y=2.5 $X2=0 $Y2=0
cc_94 N_A_94_81#_c_81_n N_A0_c_223_n 0.0167977f $X=2.715 $Y=2.5 $X2=0 $Y2=0
cc_95 N_A_94_81#_c_73_n N_A0_c_229_n 0.0123274f $X=2.03 $Y=2.415 $X2=0 $Y2=0
cc_96 N_A_94_81#_c_103_p N_A0_c_229_n 0.00104005f $X=2.385 $Y=1.44 $X2=0 $Y2=0
cc_97 N_A_94_81#_c_81_n N_A0_c_229_n 0.00197681f $X=2.715 $Y=2.5 $X2=0 $Y2=0
cc_98 N_A_94_81#_c_103_p N_A0_c_224_n 0.00298742f $X=2.385 $Y=1.44 $X2=0.24
+ $Y2=0
cc_99 N_A_94_81#_c_97_p N_A0_c_224_n 0.0200622f $X=2.47 $Y=1.355 $X2=0.24 $Y2=0
cc_100 N_A_94_81#_c_75_n N_A0_c_224_n 0.00922606f $X=2.715 $Y=0.745 $X2=0.24
+ $Y2=0
cc_101 N_A_94_81#_c_97_p N_A0_M1011_g 0.00138629f $X=2.47 $Y=1.355 $X2=5.04
+ $Y2=0
cc_102 N_A_94_81#_c_75_n N_A0_M1011_g 0.0072915f $X=2.715 $Y=0.745 $X2=5.04
+ $Y2=0
cc_103 N_A_94_81#_c_73_n N_A0_c_230_n 0.00341817f $X=2.03 $Y=2.415 $X2=2.64
+ $Y2=0.058
cc_104 N_A_94_81#_c_90_p N_A0_c_230_n 0.0239874f $X=2.55 $Y=2.5 $X2=2.64
+ $Y2=0.058
cc_105 N_A_94_81#_c_80_n N_A0_c_230_n 0.00237364f $X=2.115 $Y=2.5 $X2=2.64
+ $Y2=0.058
cc_106 N_A_94_81#_c_81_n N_A0_c_230_n 0.0107391f $X=2.715 $Y=2.5 $X2=2.64
+ $Y2=0.058
cc_107 N_A_94_81#_c_73_n N_A1_c_283_n 0.00554675f $X=2.03 $Y=2.415 $X2=0 $Y2=0
cc_108 N_A_94_81#_c_103_p N_A1_c_283_n 0.0232881f $X=2.385 $Y=1.44 $X2=0 $Y2=0
cc_109 N_A_94_81#_c_90_p N_A1_c_283_n 6.38456e-19 $X=2.55 $Y=2.5 $X2=0 $Y2=0
cc_110 N_A_94_81#_c_97_p N_A1_c_283_n 0.0103414f $X=2.47 $Y=1.355 $X2=0 $Y2=0
cc_111 N_A_94_81#_c_74_n N_A1_c_283_n 0.00278928f $X=2.03 $Y=1.44 $X2=0 $Y2=0
cc_112 N_A_94_81#_c_97_p N_A1_M1006_g 0.00818287f $X=2.47 $Y=1.355 $X2=0 $Y2=0
cc_113 N_A_94_81#_c_75_n N_A1_M1006_g 0.0161843f $X=2.715 $Y=0.745 $X2=0 $Y2=0
cc_114 N_A_94_81#_c_75_n N_A1_c_286_n 0.0027566f $X=2.715 $Y=0.745 $X2=-0.33
+ $Y2=-0.265
cc_115 N_A_94_81#_c_81_n N_A1_c_286_n 8.33971e-19 $X=2.715 $Y=2.5 $X2=-0.33
+ $Y2=-0.265
cc_116 N_A_94_81#_c_81_n N_A1_c_288_n 0.0102496f $X=2.715 $Y=2.5 $X2=0 $Y2=0
cc_117 N_A_94_81#_M1009_g X 0.0461046f $X=0.72 $Y=0.91 $X2=0.24 $Y2=0
cc_118 N_A_94_81#_c_88_p N_X_c_383_n 0.0265469f $X=0.785 $Y=1.44 $X2=2.64
+ $Y2=0.058
cc_119 N_A_94_81#_M1009_g N_X_c_383_n 0.0268613f $X=0.72 $Y=0.91 $X2=2.64
+ $Y2=0.058
cc_120 N_A_94_81#_c_72_n N_VPWR_c_397_n 0.00988032f $X=1.945 $Y=1.44 $X2=0.24
+ $Y2=0
cc_121 N_A_94_81#_c_88_p N_VPWR_c_397_n 0.0104143f $X=0.785 $Y=1.44 $X2=0.24
+ $Y2=0
cc_122 N_A_94_81#_M1009_g N_VPWR_c_397_n 0.0759589f $X=0.72 $Y=0.91 $X2=0.24
+ $Y2=0
cc_123 N_A_94_81#_M1009_g N_VPWR_c_403_n 0.0111903f $X=0.72 $Y=0.91 $X2=2.64
+ $Y2=0.058
cc_124 N_A_94_81#_c_80_n A_373_491# 0.00251327f $X=2.115 $Y=2.5 $X2=0 $Y2=0
cc_125 N_A_94_81#_c_72_n N_VGND_c_431_n 0.0733115f $X=1.945 $Y=1.44 $X2=0.24
+ $Y2=0
cc_126 N_A_94_81#_c_103_p N_VGND_c_431_n 0.00644157f $X=2.385 $Y=1.44 $X2=0.24
+ $Y2=0
cc_127 N_A_94_81#_c_97_p N_VGND_c_431_n 0.0187564f $X=2.47 $Y=1.355 $X2=0.24
+ $Y2=0
cc_128 N_A_94_81#_c_88_p N_VGND_c_431_n 0.0254318f $X=0.785 $Y=1.44 $X2=0.24
+ $Y2=0
cc_129 N_A_94_81#_c_74_n N_VGND_c_431_n 0.0149264f $X=2.03 $Y=1.44 $X2=0.24
+ $Y2=0
cc_130 N_A_94_81#_c_75_n N_VGND_c_431_n 0.0306875f $X=2.715 $Y=0.745 $X2=0.24
+ $Y2=0
cc_131 N_A_94_81#_M1009_g N_VGND_c_431_n 0.0488456f $X=0.72 $Y=0.91 $X2=0.24
+ $Y2=0
cc_132 N_A_94_81#_c_75_n N_VGND_c_433_n 0.0308395f $X=2.715 $Y=0.745 $X2=2.64
+ $Y2=0.058
cc_133 N_A_94_81#_c_97_p N_VGND_c_435_n 5.40886e-19 $X=2.47 $Y=1.355 $X2=0 $Y2=0
cc_134 N_A_94_81#_c_75_n N_VGND_c_435_n 0.0302781f $X=2.715 $Y=0.745 $X2=0 $Y2=0
cc_135 N_A_94_81#_M1009_g N_VGND_c_435_n 0.00874126f $X=0.72 $Y=0.91 $X2=0 $Y2=0
cc_136 N_S_c_176_p N_A0_c_223_n 0.00373087f $X=3.23 $Y=2.22 $X2=0 $Y2=0
cc_137 N_S_c_152_n N_A0_c_229_n 5.1915e-19 $X=1.6 $Y=1.79 $X2=0 $Y2=0
cc_138 N_S_c_176_p N_A0_c_229_n 6.22052e-19 $X=3.23 $Y=2.22 $X2=0 $Y2=0
cc_139 N_S_M1001_g N_A0_c_229_n 0.0696267f $X=1.615 $Y=0.745 $X2=0 $Y2=0
cc_140 N_S_c_152_n N_A0_c_230_n 0.00248043f $X=1.6 $Y=1.79 $X2=2.64 $Y2=0.058
cc_141 N_S_c_153_n N_A0_c_230_n 0.0164452f $X=3.06 $Y=3.18 $X2=2.64 $Y2=0.058
cc_142 N_S_c_155_n N_A0_c_230_n 9.37231e-19 $X=3.145 $Y=3.095 $X2=2.64 $Y2=0.058
cc_143 N_S_M1001_g N_A1_c_283_n 0.00759058f $X=1.615 $Y=0.745 $X2=0 $Y2=0
cc_144 N_S_M1001_g N_A1_M1006_g 0.0800556f $X=1.615 $Y=0.745 $X2=0 $Y2=0
cc_145 N_S_c_156_n A1 0.03308f $X=4.365 $Y=2.22 $X2=0 $Y2=0
cc_146 N_S_c_176_p A1 0.0111776f $X=3.23 $Y=2.22 $X2=0 $Y2=0
cc_147 N_S_M1008_g A1 6.36654e-19 $X=4.595 $Y=0.745 $X2=0 $Y2=0
cc_148 N_S_c_153_n N_A1_c_288_n 0.00887434f $X=3.06 $Y=3.18 $X2=0 $Y2=0
cc_149 N_S_c_155_n N_A1_c_288_n 0.0309744f $X=3.145 $Y=3.095 $X2=0 $Y2=0
cc_150 N_S_c_156_n N_A1_c_288_n 0.0107274f $X=4.365 $Y=2.22 $X2=0 $Y2=0
cc_151 N_S_c_176_p N_A1_c_288_n 0.00889969f $X=3.23 $Y=2.22 $X2=0 $Y2=0
cc_152 N_S_M1008_g N_A_713_81#_M1003_g 0.0154157f $X=4.595 $Y=0.745 $X2=0 $Y2=0
cc_153 N_S_c_155_n N_A_713_81#_c_338_n 0.00107088f $X=3.145 $Y=3.095 $X2=0.24
+ $Y2=0
cc_154 N_S_c_156_n N_A_713_81#_c_338_n 0.034719f $X=4.365 $Y=2.22 $X2=0.24 $Y2=0
cc_155 S N_A_713_81#_c_338_n 0.00336448f $X=4.475 $Y=1.58 $X2=0.24 $Y2=0
cc_156 N_S_M1008_g N_A_713_81#_c_338_n 0.0793996f $X=4.595 $Y=0.745 $X2=0.24
+ $Y2=0
cc_157 N_S_c_155_n N_A_713_81#_M1005_g 3.98484e-19 $X=3.145 $Y=3.095 $X2=0 $Y2=0
cc_158 N_S_M1008_g N_A_713_81#_M1005_g 0.0154157f $X=4.595 $Y=0.745 $X2=0 $Y2=0
cc_159 S N_A_713_81#_c_339_n 0.0159465f $X=4.475 $Y=1.58 $X2=5.04 $Y2=0
cc_160 N_S_M1008_g N_A_713_81#_c_339_n 0.0348893f $X=4.595 $Y=0.745 $X2=5.04
+ $Y2=0
cc_161 N_S_M1008_g N_A_713_81#_c_340_n 0.00860936f $X=4.595 $Y=0.745 $X2=2.64
+ $Y2=0
cc_162 N_S_c_156_n N_A_713_81#_c_342_n 0.0113057f $X=4.365 $Y=2.22 $X2=2.64
+ $Y2=0.058
cc_163 S N_A_713_81#_c_342_n 0.0365203f $X=4.475 $Y=1.58 $X2=2.64 $Y2=0.058
cc_164 N_S_M1008_g N_A_713_81#_c_342_n 0.0436763f $X=4.595 $Y=0.745 $X2=2.64
+ $Y2=0.058
cc_165 N_S_c_156_n N_A_713_81#_c_360_n 0.0103788f $X=4.365 $Y=2.22 $X2=0 $Y2=0
cc_166 S N_A_713_81#_c_360_n 0.0120899f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_167 N_S_M1008_g N_A_713_81#_c_360_n 0.00278011f $X=4.595 $Y=0.745 $X2=0 $Y2=0
cc_168 N_S_c_152_n N_VPWR_c_397_n 0.0718349f $X=1.6 $Y=1.79 $X2=0.24 $Y2=0
cc_169 N_S_c_154_n N_VPWR_c_397_n 0.0147522f $X=1.765 $Y=3.18 $X2=0.24 $Y2=0
cc_170 N_S_M1001_g N_VPWR_c_397_n 0.00840955f $X=1.615 $Y=0.745 $X2=0.24 $Y2=0
cc_171 N_S_c_153_n N_VPWR_c_400_n 0.0152318f $X=3.06 $Y=3.18 $X2=0 $Y2=0
cc_172 N_S_c_155_n N_VPWR_c_400_n 0.0294963f $X=3.145 $Y=3.095 $X2=0 $Y2=0
cc_173 N_S_c_156_n N_VPWR_c_400_n 0.0859615f $X=4.365 $Y=2.22 $X2=0 $Y2=0
cc_174 N_S_M1008_g N_VPWR_c_400_n 0.043583f $X=4.595 $Y=0.745 $X2=0 $Y2=0
cc_175 N_S_c_153_n N_VPWR_c_403_n 0.0737737f $X=3.06 $Y=3.18 $X2=2.64 $Y2=0.058
cc_176 N_S_c_154_n N_VPWR_c_403_n 0.0187303f $X=1.765 $Y=3.18 $X2=2.64 $Y2=0.058
cc_177 N_S_M1001_g N_VPWR_c_403_n 0.00191289f $X=1.615 $Y=0.745 $X2=2.64
+ $Y2=0.058
cc_178 N_S_M1008_g N_VPWR_c_403_n 0.00338982f $X=4.595 $Y=0.745 $X2=2.64
+ $Y2=0.058
cc_179 N_S_M1001_g N_VGND_c_431_n 0.0700333f $X=1.615 $Y=0.745 $X2=0.24 $Y2=0
cc_180 N_S_M1008_g N_VGND_c_433_n 0.0357772f $X=4.595 $Y=0.745 $X2=2.64
+ $Y2=0.058
cc_181 N_S_M1008_g N_VGND_c_435_n 0.00504702f $X=4.595 $Y=0.745 $X2=0 $Y2=0
cc_182 N_A0_c_222_n N_A1_c_283_n 0.00596893f $X=2.82 $Y=1.785 $X2=0 $Y2=0
cc_183 N_A0_c_223_n N_A1_c_283_n 0.00883921f $X=2.46 $Y=2.13 $X2=0 $Y2=0
cc_184 N_A0_c_229_n N_A1_c_283_n 0.0377405f $X=2.46 $Y=2.13 $X2=0 $Y2=0
cc_185 N_A0_c_224_n N_A1_c_283_n 0.00231902f $X=2.905 $Y=1.242 $X2=0 $Y2=0
cc_186 N_A0_M1011_g N_A1_c_283_n 0.016933f $X=3.105 $Y=0.745 $X2=0 $Y2=0
cc_187 N_A0_M1011_g N_A1_M1006_g 0.014941f $X=3.105 $Y=0.745 $X2=0 $Y2=0
cc_188 N_A0_c_222_n N_A1_c_286_n 0.0135855f $X=2.82 $Y=1.785 $X2=-0.33
+ $Y2=-0.265
cc_189 A0 N_A1_c_286_n 0.00167535f $X=3.515 $Y=1.21 $X2=-0.33 $Y2=-0.265
cc_190 N_A0_M1011_g N_A1_c_286_n 0.0349758f $X=3.105 $Y=0.745 $X2=-0.33
+ $Y2=-0.265
cc_191 N_A0_c_222_n A1 0.0155817f $X=2.82 $Y=1.785 $X2=0 $Y2=0
cc_192 N_A0_c_223_n A1 0.0134167f $X=2.46 $Y=2.13 $X2=0 $Y2=0
cc_193 A0 A1 0.0460436f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A0_M1011_g A1 0.00172967f $X=3.105 $Y=0.745 $X2=0 $Y2=0
cc_195 N_A0_c_222_n N_A1_c_288_n 9.79366e-19 $X=2.82 $Y=1.785 $X2=0 $Y2=0
cc_196 N_A0_c_223_n N_A1_c_288_n 0.0110653f $X=2.46 $Y=2.13 $X2=0 $Y2=0
cc_197 N_A0_c_229_n N_A1_c_288_n 0.0275095f $X=2.46 $Y=2.13 $X2=0 $Y2=0
cc_198 N_A0_c_230_n N_A1_c_288_n 0.013887f $X=2.36 $Y=2.345 $X2=0 $Y2=0
cc_199 N_A0_M1011_g N_A_713_81#_M1003_g 0.0670903f $X=3.105 $Y=0.745 $X2=0 $Y2=0
cc_200 N_A0_c_222_n N_A_713_81#_c_338_n 0.00444148f $X=2.82 $Y=1.785 $X2=0.24
+ $Y2=0
cc_201 A0 N_A_713_81#_c_338_n 0.0137458f $X=3.515 $Y=1.21 $X2=0.24 $Y2=0
cc_202 A0 N_A_713_81#_c_360_n 0.0222228f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_203 N_A0_M1011_g N_VGND_c_431_n 5.95043e-19 $X=3.105 $Y=0.745 $X2=0.24 $Y2=0
cc_204 A0 N_VGND_c_433_n 0.0408688f $X=3.515 $Y=1.21 $X2=2.64 $Y2=0.058
cc_205 N_A0_M1011_g N_VGND_c_433_n 0.0343767f $X=3.105 $Y=0.745 $X2=2.64
+ $Y2=0.058
cc_206 N_A0_c_224_n N_VGND_c_435_n 0.00153694f $X=2.905 $Y=1.242 $X2=0 $Y2=0
cc_207 A0 N_VGND_c_435_n 0.00744178f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_208 N_A0_M1011_g N_VGND_c_435_n 0.00527908f $X=3.105 $Y=0.745 $X2=0 $Y2=0
cc_209 N_A1_c_286_n N_A_713_81#_c_338_n 0.0473498f $X=2.855 $Y=1.68 $X2=0.24
+ $Y2=0
cc_210 A1 N_A_713_81#_c_338_n 0.0188359f $X=3.515 $Y=1.58 $X2=0.24 $Y2=0
cc_211 N_A1_c_288_n N_A_713_81#_M1005_g 0.0473498f $X=3.17 $Y=1.79 $X2=0 $Y2=0
cc_212 A1 N_A_713_81#_c_360_n 0.0150897f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_213 N_A1_c_288_n N_VPWR_c_400_n 0.00270923f $X=3.17 $Y=1.79 $X2=0 $Y2=0
cc_214 N_A1_c_288_n N_VPWR_c_403_n 0.00339257f $X=3.17 $Y=1.79 $X2=2.64
+ $Y2=0.058
cc_215 N_A1_c_283_n N_VGND_c_431_n 0.00515068f $X=2.325 $Y=1.085 $X2=0.24 $Y2=0
cc_216 N_A1_M1006_g N_VGND_c_431_n 0.0260486f $X=2.325 $Y=0.745 $X2=0.24 $Y2=0
cc_217 N_A1_M1006_g N_VGND_c_433_n 8.23157e-19 $X=2.325 $Y=0.745 $X2=2.64
+ $Y2=0.058
cc_218 N_A1_M1006_g N_VGND_c_435_n 0.0126453f $X=2.325 $Y=0.745 $X2=0 $Y2=0
cc_219 N_A_713_81#_M1005_g N_VPWR_c_400_n 0.0481996f $X=3.815 $Y=2.665 $X2=0
+ $Y2=0
cc_220 N_A_713_81#_c_342_n N_VPWR_c_400_n 0.0183139f $X=4.985 $Y=2.665 $X2=0
+ $Y2=0
cc_221 N_A_713_81#_c_342_n N_VPWR_c_403_n 0.0100913f $X=4.985 $Y=2.665 $X2=2.64
+ $Y2=0.058
cc_222 N_A_713_81#_M1003_g N_VGND_c_433_n 0.0515995f $X=3.815 $Y=0.745 $X2=2.64
+ $Y2=0.058
cc_223 N_A_713_81#_c_338_n N_VGND_c_433_n 0.00172996f $X=3.815 $Y=2.325 $X2=2.64
+ $Y2=0.058
cc_224 N_A_713_81#_c_339_n N_VGND_c_433_n 0.0380785f $X=4.9 $Y=1.19 $X2=2.64
+ $Y2=0.058
cc_225 N_A_713_81#_c_340_n N_VGND_c_433_n 0.0185197f $X=4.985 $Y=0.745 $X2=2.64
+ $Y2=0.058
cc_226 N_A_713_81#_c_360_n N_VGND_c_433_n 0.0160761f $X=3.95 $Y=1.27 $X2=2.64
+ $Y2=0.058
cc_227 N_A_713_81#_M1008_d N_VGND_c_435_n 6.6843e-19 $X=4.845 $Y=0.535 $X2=0
+ $Y2=0
cc_228 N_A_713_81#_c_339_n N_VGND_c_435_n 0.00801952f $X=4.9 $Y=1.19 $X2=0 $Y2=0
cc_229 N_A_713_81#_c_340_n N_VGND_c_435_n 0.0263695f $X=4.985 $Y=0.745 $X2=0
+ $Y2=0
cc_230 N_A_713_81#_c_360_n N_VGND_c_435_n 0.00105268f $X=3.95 $Y=1.27 $X2=0
+ $Y2=0
cc_231 X N_VPWR_c_397_n 0.114975f $X=0.155 $Y=1.95 $X2=0.24 $Y2=0
cc_232 X N_VPWR_c_403_n 0.0468685f $X=0.155 $Y=1.95 $X2=2.64 $Y2=0.058
cc_233 N_X_c_383_n N_VGND_c_431_n 0.0288929f $X=0.33 $Y=0.66 $X2=0.24 $Y2=0
cc_234 N_X_M1009_s N_VGND_c_435_n 0.00221032f $X=0.185 $Y=0.535 $X2=0 $Y2=0
cc_235 N_X_c_383_n N_VGND_c_435_n 0.0298505f $X=0.33 $Y=0.66 $X2=0 $Y2=0
cc_236 N_VPWR_c_400_n A_671_491# 0.00111679f $X=4.205 $Y=2.665 $X2=0 $Y2=3.985
cc_237 N_VGND_c_433_n A_671_107# 0.00108638f $X=4.61 $Y=0.48 $X2=0 $Y2=0
