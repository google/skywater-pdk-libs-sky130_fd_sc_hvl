# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
SITE unithvdbl
    SYMMETRY y  ;
    CLASS CORE  ;
    SIZE  0.480 BY 8.140 ;
END unithvdbl
MACRO sky130_fd_sc_hvl__lsbufhv2hv_lh_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  8.140000 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    ANTENNAGATEAREA  0.750000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.495000 1.530000 2.805000 2.200000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.120000 4.405000 10.450000 7.625000 ;
    END
  END X
  PIN LOWHVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 3.590000 3.355000 4.780000 4.025000 ;
        RECT 3.740000 2.325000 4.330000 3.355000 ;
    END
    PORT
      LAYER mcon ;
        RECT 3.770000 3.050000 3.940000 3.220000 ;
        RECT 4.130000 3.050000 4.300000 3.220000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 10.490000 3.305000 ;
    END
  END LOWHVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 3.300000 6.085000 3.890000 7.715000 ;
        RECT 3.300000 7.715000 7.010000 7.885000 ;
        RECT 4.860000 6.165000 5.450000 7.715000 ;
        RECT 6.420000 6.165000 7.010000 7.715000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.740000 0.255000 9.540000 0.425000 ;
        RECT 3.740000 0.425000 4.330000 1.475000 ;
        RECT 5.830000 0.425000 6.420000 1.975000 ;
        RECT 7.390000 0.425000 7.980000 1.975000 ;
        RECT 8.950000 0.425000 9.540000 1.975000 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.210000 6.835000 9.800000 7.745000 ;
    END
    PORT
      LAYER mcon ;
        RECT 3.330000 7.545000 3.500000 7.715000 ;
        RECT 3.690000 7.545000 3.860000 7.715000 ;
        RECT 3.770000 0.425000 3.940000 0.595000 ;
        RECT 4.130000 0.425000 4.300000 0.595000 ;
        RECT 4.890000 7.545000 5.060000 7.715000 ;
        RECT 5.250000 7.545000 5.420000 7.715000 ;
        RECT 5.860000 0.425000 6.030000 0.595000 ;
        RECT 6.220000 0.425000 6.390000 0.595000 ;
        RECT 6.450000 7.545000 6.620000 7.715000 ;
        RECT 6.810000 7.545000 6.980000 7.715000 ;
        RECT 7.420000 0.425000 7.590000 0.595000 ;
        RECT 7.780000 0.425000 7.950000 0.595000 ;
        RECT 8.980000 0.425000 9.150000 0.595000 ;
        RECT 9.240000 7.545000 9.410000 7.715000 ;
        RECT 9.340000 0.425000 9.510000 0.595000 ;
        RECT 9.600000 7.545000 9.770000 7.715000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 10.560000 0.625000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 10.560000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.560000 0.085000 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000000 8.055000 10.560000 8.225000 ;
    END
    PORT
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.155000  8.055000  0.325000 8.225000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  0.635000  8.055000  0.805000 8.225000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.115000  8.055000  1.285000 8.225000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  1.595000  8.055000  1.765000 8.225000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.075000  8.055000  2.245000 8.225000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  2.555000  8.055000  2.725000 8.225000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.035000  8.055000  3.205000 8.225000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.515000  8.055000  3.685000 8.225000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  3.995000  8.055000  4.165000 8.225000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.475000  8.055000  4.645000 8.225000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  4.955000  8.055000  5.125000 8.225000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.435000  8.055000  5.605000 8.225000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  5.915000  8.055000  6.085000 8.225000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.395000  8.055000  6.565000 8.225000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  6.875000  8.055000  7.045000 8.225000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.355000  8.055000  7.525000 8.225000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  7.835000  8.055000  8.005000 8.225000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.315000  8.055000  8.485000 8.225000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  8.795000  8.055000  8.965000 8.225000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.275000  8.055000  9.445000 8.225000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT  9.755000  8.055000  9.925000 8.225000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.235000  8.055000 10.405000 8.225000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 10.560000 0.115000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 10.560000 8.255000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 0.800000 4.155000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.715000 3.985000 10.560000 4.155000 ;
    END
    PORT
      LAYER mcon ;
        RECT  0.155000 3.985000  0.325000 4.155000 ;
        RECT  8.795000 3.985000  8.965000 4.155000 ;
        RECT  9.275000 3.985000  9.445000 4.155000 ;
        RECT  9.755000 3.985000  9.925000 4.155000 ;
        RECT 10.235000 3.985000 10.405000 4.155000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 10.560000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 8.790000 4.405000 9.800000 4.800000 ;
        RECT 9.210000 4.800000 9.800000 5.945000 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.940000 2.795000 9.530000 3.705000 ;
    END
    PORT
      LAYER mcon ;
        RECT 8.880000 4.495000 9.050000 4.665000 ;
        RECT 8.970000 3.475000 9.140000 3.645000 ;
        RECT 9.240000 4.495000 9.410000 4.665000 ;
        RECT 9.330000 3.475000 9.500000 3.645000 ;
        RECT 9.600000 4.495000 9.770000 4.665000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 10.560000 3.815000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 10.560000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 3.090000 0.685000 3.420000 1.745000 ;
      RECT 3.090000 1.745000 4.845000 1.995000 ;
      RECT 3.090000 1.995000 3.420000 5.165000 ;
      RECT 3.090000 5.165000 5.660000 5.495000 ;
      RECT 4.210000 5.665000 7.930000 5.995000 ;
      RECT 4.210000 5.995000 4.540000 7.545000 ;
      RECT 4.650000 0.685000 4.980000 1.145000 ;
      RECT 4.650000 1.145000 5.660000 1.475000 ;
      RECT 4.650000 2.165000 6.570000 2.475000 ;
      RECT 4.650000 2.475000 4.980000 3.115000 ;
      RECT 5.330000 1.475000 5.660000 2.145000 ;
      RECT 5.330000 2.145000 6.570000 2.165000 ;
      RECT 5.770000 5.995000 6.100000 7.545000 ;
      RECT 6.740000 0.595000 7.070000 2.145000 ;
      RECT 6.740000 2.145000 8.630000 2.475000 ;
      RECT 7.375000 3.605000 8.045000 3.935000 ;
      RECT 7.600000 2.795000 8.545000 3.125000 ;
      RECT 7.600000 3.125000 7.930000 3.435000 ;
      RECT 7.600000 3.935000 7.930000 5.665000 ;
      RECT 8.215000 2.475000 8.545000 2.795000 ;
      RECT 8.215000 3.125000 8.545000 5.205000 ;
      RECT 8.215000 5.205000 8.965000 5.535000 ;
      RECT 8.300000 0.595000 8.630000 2.145000 ;
      RECT 8.635000 5.535000 8.965000 6.555000 ;
  END
END sky130_fd_sc_hvl__lsbufhv2hv_lh_1
END LIBRARY
