* File: sky130_fd_sc_hvl__decap_4.pxi.spice
* Created: Wed Sep  2 09:04:42 2020
* 
x_PM_SKY130_FD_SC_HVL__DECAP_4%VNB N_VNB_M1000_b VNB N_VNB_c_4_p VNB
+ PM_SKY130_FD_SC_HVL__DECAP_4%VNB
x_PM_SKY130_FD_SC_HVL__DECAP_4%VPB N_VPB_M1001_b VPB N_VPB_c_13_p VPB
+ PM_SKY130_FD_SC_HVL__DECAP_4%VPB
x_PM_SKY130_FD_SC_HVL__DECAP_4%VGND N_VGND_M1000_s N_VGND_M1001_g N_VGND_c_23_n
+ N_VGND_c_24_n VGND N_VGND_c_27_n N_VGND_c_29_n
+ PM_SKY130_FD_SC_HVL__DECAP_4%VGND
x_PM_SKY130_FD_SC_HVL__DECAP_4%VPWR N_VPWR_M1001_s N_VPWR_c_49_n N_VPWR_M1000_g
+ N_VPWR_c_51_n N_VPWR_c_50_n VPWR N_VPWR_c_53_n N_VPWR_c_56_n
+ PM_SKY130_FD_SC_HVL__DECAP_4%VPWR
cc_1 N_VNB_M1000_b N_VGND_c_23_n 0.0107972f $X=-0.33 $Y=-0.265 $X2=0.64
+ $Y2=1.865
cc_2 N_VNB_M1000_b N_VGND_c_24_n 0.0225594f $X=-0.33 $Y=-0.265 $X2=0.64
+ $Y2=1.865
cc_3 N_VNB_M1000_b VGND 0.0587464f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0.255
cc_4 N_VNB_c_4_p VGND 0.205241f $X=0.24 $Y=0 $X2=0 $Y2=0.255
cc_5 N_VNB_M1000_b N_VGND_c_27_n 0.0460398f $X=-0.33 $Y=-0.265 $X2=0.805
+ $Y2=0.807
cc_6 N_VNB_c_4_p N_VGND_c_27_n 0.00180697f $X=0.24 $Y=0 $X2=0.805 $Y2=0.807
cc_7 N_VNB_M1000_b N_VGND_c_29_n 0.0782402f $X=-0.33 $Y=-0.265 $X2=1.615
+ $Y2=0.81
cc_8 N_VNB_c_4_p N_VGND_c_29_n 0.00276229f $X=0.24 $Y=0 $X2=1.615 $Y2=0.81
cc_9 N_VNB_M1000_b N_VPWR_c_49_n 0.107645f $X=-0.33 $Y=-0.265 $X2=0.64 $Y2=2.575
cc_10 N_VNB_M1000_b N_VPWR_c_50_n 0.0504004f $X=-0.33 $Y=-0.265 $X2=0.64
+ $Y2=1.865
cc_11 N_VPB_M1001_b N_VGND_M1001_g 0.0980196f $X=-0.33 $Y=1.885 $X2=0.975
+ $Y2=3.205
cc_12 VPB N_VGND_M1001_g 0.0192755f $X=0 $Y=3.955 $X2=0.975 $Y2=3.205
cc_13 N_VPB_c_13_p N_VGND_M1001_g 0.0270955f $X=1.68 $Y=4.07 $X2=0.975 $Y2=3.205
cc_14 N_VPB_M1001_b N_VGND_c_24_n 0.075174f $X=-0.33 $Y=1.885 $X2=0.64 $Y2=1.865
cc_15 N_VPB_M1001_b N_VPWR_c_51_n 0.0283976f $X=-0.33 $Y=1.885 $X2=0.64 $Y2=1.25
cc_16 N_VPB_M1001_b N_VPWR_c_50_n 0.0278937f $X=-0.33 $Y=1.885 $X2=0.64
+ $Y2=1.865
cc_17 N_VPB_M1001_b N_VPWR_c_53_n 0.0502013f $X=-0.33 $Y=1.885 $X2=0.3 $Y2=0.48
cc_18 VPB N_VPWR_c_53_n 0.20361f $X=0 $Y=3.955 $X2=0.3 $Y2=0.48
cc_19 N_VPB_c_13_p N_VPWR_c_53_n 0.00844f $X=1.68 $Y=4.07 $X2=0.3 $Y2=0.48
cc_20 N_VPB_M1001_b N_VPWR_c_56_n 0.023387f $X=-0.33 $Y=1.885 $X2=0.335
+ $Y2=0.807
cc_21 VPB N_VPWR_c_56_n 0.00617543f $X=0 $Y=3.955 $X2=0.335 $Y2=0.807
cc_22 N_VPB_c_13_p N_VPWR_c_56_n 0.0723308f $X=1.68 $Y=4.07 $X2=0.335 $Y2=0.807
cc_23 N_VGND_c_23_n N_VPWR_c_49_n 0.029299f $X=0.64 $Y=1.865 $X2=0 $Y2=0
cc_24 N_VGND_c_24_n N_VPWR_c_49_n 0.0198526f $X=0.64 $Y=1.865 $X2=0 $Y2=0
cc_25 N_VGND_c_27_n N_VPWR_c_49_n 0.0392278f $X=0.805 $Y=0.807 $X2=0 $Y2=0
cc_26 N_VGND_c_29_n N_VPWR_c_49_n 0.0917584f $X=1.615 $Y=0.81 $X2=0 $Y2=0
cc_27 N_VGND_M1001_g N_VPWR_c_51_n 0.0201449f $X=0.975 $Y=3.205 $X2=0 $Y2=0
cc_28 N_VGND_c_23_n N_VPWR_c_51_n 0.0209133f $X=0.64 $Y=1.865 $X2=0 $Y2=0
cc_29 N_VGND_c_24_n N_VPWR_c_51_n 0.0222329f $X=0.64 $Y=1.865 $X2=0 $Y2=0
cc_30 N_VGND_c_29_n N_VPWR_c_51_n 0.0125221f $X=1.615 $Y=0.81 $X2=0 $Y2=0
cc_31 N_VGND_M1001_g N_VPWR_c_50_n 0.0093132f $X=0.975 $Y=3.205 $X2=0 $Y2=0
cc_32 N_VGND_c_23_n N_VPWR_c_50_n 0.0102577f $X=0.64 $Y=1.865 $X2=0 $Y2=0
cc_33 N_VGND_c_24_n N_VPWR_c_50_n 0.0206283f $X=0.64 $Y=1.865 $X2=0 $Y2=0
cc_34 N_VGND_M1001_g N_VPWR_c_53_n 0.00398809f $X=0.975 $Y=3.205 $X2=0 $Y2=0
cc_35 N_VGND_M1001_g N_VPWR_c_56_n 0.130335f $X=0.975 $Y=3.205 $X2=0 $Y2=0
cc_36 N_VGND_c_23_n N_VPWR_c_56_n 0.00894257f $X=0.64 $Y=1.865 $X2=0 $Y2=0
