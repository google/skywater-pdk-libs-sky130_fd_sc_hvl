* File: sky130_fd_sc_hvl__dlclkp_1.pxi.spice
* Created: Fri Aug 28 09:34:56 2020
* 
x_PM_SKY130_FD_SC_HVL__DLCLKP_1%VNB N_VNB_M1002_b VNB N_VNB_c_3_p VNB
+ PM_SKY130_FD_SC_HVL__DLCLKP_1%VNB
x_PM_SKY130_FD_SC_HVL__DLCLKP_1%VPB N_VPB_M1000_b VPB N_VPB_c_97_p N_VPB_c_98_p
+ VPB PM_SKY130_FD_SC_HVL__DLCLKP_1%VPB
x_PM_SKY130_FD_SC_HVL__DLCLKP_1%GATE GATE GATE N_GATE_M1002_g N_GATE_c_181_p
+ N_GATE_M1000_g PM_SKY130_FD_SC_HVL__DLCLKP_1%GATE
x_PM_SKY130_FD_SC_HVL__DLCLKP_1%A_231_71# N_A_231_71#_M1005_d
+ N_A_231_71#_M1006_d N_A_231_71#_M1012_g N_A_231_71#_M1013_g
+ N_A_231_71#_c_192_n N_A_231_71#_c_194_n N_A_231_71#_c_196_n
+ N_A_231_71#_c_217_p N_A_231_71#_c_218_p N_A_231_71#_c_198_n
+ N_A_231_71#_c_199_n N_A_231_71#_c_200_n N_A_231_71#_c_207_n
+ N_A_231_71#_c_208_n N_A_231_71#_c_209_n N_A_231_71#_c_201_n
+ N_A_231_71#_c_219_p N_A_231_71#_c_202_n N_A_231_71#_M1017_g
+ N_A_231_71#_M1018_g N_A_231_71#_c_204_n
+ PM_SKY130_FD_SC_HVL__DLCLKP_1%A_231_71#
x_PM_SKY130_FD_SC_HVL__DLCLKP_1%A_239_419# N_A_239_419#_M1017_s
+ N_A_239_419#_M1018_s N_A_239_419#_M1007_g N_A_239_419#_M1004_g
+ N_A_239_419#_c_312_n N_A_239_419#_c_313_n N_A_239_419#_c_307_n
+ N_A_239_419#_c_315_n N_A_239_419#_c_316_n N_A_239_419#_c_317_n
+ N_A_239_419#_c_318_n N_A_239_419#_c_321_n N_A_239_419#_c_308_n
+ N_A_239_419#_c_325_n N_A_239_419#_c_326_n N_A_239_419#_c_309_n
+ N_A_239_419#_c_327_n N_A_239_419#_c_353_n N_A_239_419#_c_310_n
+ N_A_239_419#_c_355_n PM_SKY130_FD_SC_HVL__DLCLKP_1%A_239_419#
x_PM_SKY130_FD_SC_HVL__DLCLKP_1%A_1069_133# N_A_1069_133#_M1001_d
+ N_A_1069_133#_M1008_d N_A_1069_133#_M1009_g N_A_1069_133#_M1014_g
+ N_A_1069_133#_c_447_n N_A_1069_133#_c_429_n N_A_1069_133#_c_430_n
+ N_A_1069_133#_c_438_n N_A_1069_133#_c_431_n N_A_1069_133#_c_439_n
+ N_A_1069_133#_c_432_n N_A_1069_133#_c_433_n N_A_1069_133#_c_478_p
+ N_A_1069_133#_M1015_g N_A_1069_133#_M1003_g
+ PM_SKY130_FD_SC_HVL__DLCLKP_1%A_1069_133#
x_PM_SKY130_FD_SC_HVL__DLCLKP_1%A_303_311# N_A_303_311#_M1012_d
+ N_A_303_311#_M1004_s N_A_303_311#_M1007_d N_A_303_311#_M1013_s
+ N_A_303_311#_c_506_n N_A_303_311#_c_507_n N_A_303_311#_c_508_n
+ N_A_303_311#_c_510_n N_A_303_311#_c_512_n N_A_303_311#_c_514_n
+ N_A_303_311#_c_515_n N_A_303_311#_c_528_n N_A_303_311#_c_516_n
+ N_A_303_311#_c_517_n N_A_303_311#_c_533_n N_A_303_311#_c_518_n
+ N_A_303_311#_c_520_n N_A_303_311#_c_555_n N_A_303_311#_c_521_n
+ N_A_303_311#_c_592_n N_A_303_311#_c_522_n N_A_303_311#_c_524_n
+ N_A_303_311#_M1001_g N_A_303_311#_M1008_g
+ PM_SKY130_FD_SC_HVL__DLCLKP_1%A_303_311#
x_PM_SKY130_FD_SC_HVL__DLCLKP_1%CLK N_CLK_c_647_n N_CLK_M1006_g N_CLK_c_648_n
+ N_CLK_c_649_n N_CLK_c_650_n N_CLK_c_651_n N_CLK_c_654_n N_CLK_c_657_n
+ N_CLK_c_658_n N_CLK_c_659_n N_CLK_c_660_n N_CLK_c_661_n N_CLK_c_662_n
+ N_CLK_c_698_n CLK N_CLK_M1005_g N_CLK_M1011_g N_CLK_M1019_g
+ PM_SKY130_FD_SC_HVL__DLCLKP_1%CLK
x_PM_SKY130_FD_SC_HVL__DLCLKP_1%A_1438_171# N_A_1438_171#_M1015_s
+ N_A_1438_171#_M1003_d N_A_1438_171#_M1010_g N_A_1438_171#_M1016_g
+ N_A_1438_171#_c_748_n N_A_1438_171#_c_749_n N_A_1438_171#_c_750_n
+ N_A_1438_171#_c_751_n N_A_1438_171#_c_752_n N_A_1438_171#_c_753_n
+ N_A_1438_171#_c_754_n N_A_1438_171#_c_755_n
+ PM_SKY130_FD_SC_HVL__DLCLKP_1%A_1438_171#
x_PM_SKY130_FD_SC_HVL__DLCLKP_1%VPWR N_VPWR_M1000_s N_VPWR_M1018_d
+ N_VPWR_M1014_d N_VPWR_M1003_s N_VPWR_M1019_d N_VPWR_c_806_n N_VPWR_c_807_n
+ N_VPWR_c_808_n N_VPWR_c_811_n N_VPWR_c_812_n N_VPWR_c_815_n N_VPWR_c_816_n
+ N_VPWR_c_817_n N_VPWR_c_820_n N_VPWR_c_823_n N_VPWR_c_826_n VPWR
+ N_VPWR_c_827_n N_VPWR_c_830_n N_VPWR_c_831_n N_VPWR_c_832_n N_VPWR_c_833_n
+ N_VPWR_c_834_n N_VPWR_c_835_n VPWR PM_SKY130_FD_SC_HVL__DLCLKP_1%VPWR
x_PM_SKY130_FD_SC_HVL__DLCLKP_1%GCLK N_GCLK_M1010_d N_GCLK_M1016_d
+ N_GCLK_c_918_n GCLK GCLK GCLK GCLK GCLK PM_SKY130_FD_SC_HVL__DLCLKP_1%GCLK
x_PM_SKY130_FD_SC_HVL__DLCLKP_1%VGND N_VGND_M1002_s N_VGND_M1017_d
+ N_VGND_M1009_d N_VGND_M1011_d N_VGND_c_939_n N_VGND_c_940_n N_VGND_c_942_n
+ N_VGND_c_943_n N_VGND_c_944_n VGND N_VGND_c_946_n N_VGND_c_948_n
+ N_VGND_c_950_n N_VGND_c_952_n N_VGND_c_954_n N_VGND_c_955_n VGND
+ PM_SKY130_FD_SC_HVL__DLCLKP_1%VGND
cc_1 N_VNB_M1002_b N_GATE_M1002_g 0.126162f $X=-0.33 $Y=-0.265 $X2=0.695
+ $Y2=1.005
cc_2 N_VNB_M1002_b N_A_231_71#_c_192_n 0.0634507f $X=-0.33 $Y=-0.265 $X2=0.775
+ $Y2=1.55
cc_3 N_VNB_c_3_p N_A_231_71#_c_192_n 0.00550194f $X=9.84 $Y=0 $X2=0.775 $Y2=1.55
cc_4 N_VNB_M1002_b N_A_231_71#_c_194_n 0.0743713f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_5 N_VNB_c_3_p N_A_231_71#_c_194_n 0.00328416f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_6 N_VNB_M1002_b N_A_231_71#_c_196_n 0.0152894f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_7 N_VNB_c_3_p N_A_231_71#_c_196_n 4.82472e-19 $X=9.84 $Y=0 $X2=0 $Y2=0
cc_8 N_VNB_M1002_b N_A_231_71#_c_198_n 0.0126815f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_M1002_b N_A_231_71#_c_199_n 0.00277336f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_10 N_VNB_M1002_b N_A_231_71#_c_200_n 0.0129133f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_11 N_VNB_M1002_b N_A_231_71#_c_201_n 0.00224896f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1002_b N_A_231_71#_c_202_n 0.00367317f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1002_b N_A_231_71#_M1017_g 0.0908702f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_M1002_b N_A_231_71#_c_204_n 0.0421391f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_15 N_VNB_M1002_b N_A_239_419#_M1004_g 0.0604877f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_16 N_VNB_M1002_b N_A_239_419#_c_307_n 0.0151404f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_17 N_VNB_M1002_b N_A_239_419#_c_308_n 0.00363766f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_18 N_VNB_M1002_b N_A_239_419#_c_309_n 0.00564967f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_19 N_VNB_M1002_b N_A_239_419#_c_310_n 0.0335596f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_20 N_VNB_M1002_b N_A_1069_133#_M1009_g 0.0338f $X=-0.33 $Y=-0.265 $X2=0.775
+ $Y2=1.55
cc_21 N_VNB_M1002_b N_A_1069_133#_c_429_n 0.0397895f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_22 N_VNB_M1002_b N_A_1069_133#_c_430_n 0.00536223f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_23 N_VNB_M1002_b N_A_1069_133#_c_431_n 0.0148799f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_24 N_VNB_M1002_b N_A_1069_133#_c_432_n 0.0265939f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_25 N_VNB_M1002_b N_A_1069_133#_c_433_n 0.00508451f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_26 N_VNB_M1002_b N_A_1069_133#_M1015_g 0.0909271f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_27 N_VNB_M1002_b N_A_303_311#_c_506_n 0.069934f $X=-0.33 $Y=-0.265 $X2=0.775
+ $Y2=1.55
cc_28 N_VNB_M1002_b N_A_303_311#_c_507_n 0.105057f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_29 N_VNB_M1002_b N_A_303_311#_c_508_n 0.0663755f $X=-0.33 $Y=-0.265 $X2=0.775
+ $Y2=1.665
cc_30 N_VNB_c_3_p N_A_303_311#_c_508_n 0.0316377f $X=9.84 $Y=0 $X2=0.775
+ $Y2=1.665
cc_31 N_VNB_M1002_b N_A_303_311#_c_510_n 0.119956f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_32 N_VNB_c_3_p N_A_303_311#_c_510_n 0.00150618f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_33 N_VNB_M1002_b N_A_303_311#_c_512_n 0.0516893f $X=-0.33 $Y=-0.265 $X2=0.775
+ $Y2=2.035
cc_34 N_VNB_c_3_p N_A_303_311#_c_512_n 0.00276103f $X=9.84 $Y=0 $X2=0.775
+ $Y2=2.035
cc_35 N_VNB_M1002_b N_A_303_311#_c_514_n 0.053714f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_36 N_VNB_M1002_b N_A_303_311#_c_515_n 0.0142313f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_37 N_VNB_M1002_b N_A_303_311#_c_516_n 0.0045155f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_38 N_VNB_M1002_b N_A_303_311#_c_517_n 0.0125159f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_39 N_VNB_M1002_b N_A_303_311#_c_518_n 0.0406009f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_c_3_p N_A_303_311#_c_518_n 0.00229126f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_41 N_VNB_M1002_b N_A_303_311#_c_520_n 0.00549533f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_42 N_VNB_M1002_b N_A_303_311#_c_521_n 0.0106611f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_43 N_VNB_M1002_b N_A_303_311#_c_522_n 0.026646f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_44 N_VNB_c_3_p N_A_303_311#_c_522_n 0.00261574f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_45 N_VNB_M1002_b N_A_303_311#_c_524_n 0.0938162f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_c_3_p N_A_303_311#_c_524_n 0.00309187f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_47 N_VNB_M1002_b N_A_303_311#_M1001_g 0.0767951f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_M1002_b N_CLK_M1005_g 0.0947429f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_49 N_VNB_M1002_b N_CLK_M1011_g 0.0787159f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_50 N_VNB_M1002_b N_A_1438_171#_M1016_g 0.0159007f $X=-0.33 $Y=-0.265
+ $X2=0.695 $Y2=2.6
cc_51 N_VNB_M1002_b N_A_1438_171#_c_748_n 0.00402158f $X=-0.33 $Y=-0.265
+ $X2=0.775 $Y2=1.55
cc_52 N_VNB_M1002_b N_A_1438_171#_c_749_n 0.0020232f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_53 N_VNB_M1002_b N_A_1438_171#_c_750_n 0.00617865f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_54 N_VNB_M1002_b N_A_1438_171#_c_751_n 5.41891e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_55 N_VNB_M1002_b N_A_1438_171#_c_752_n 0.00315839f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_56 N_VNB_M1002_b N_A_1438_171#_c_753_n 0.0468203f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_57 N_VNB_M1002_b N_A_1438_171#_c_754_n 0.0106063f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_58 N_VNB_M1002_b N_A_1438_171#_c_755_n 0.0450387f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_59 N_VNB_c_3_p N_A_1438_171#_c_755_n 5.3528e-19 $X=9.84 $Y=0 $X2=0 $Y2=0
cc_60 N_VNB_M1002_b N_GCLK_c_918_n 0.0321523f $X=-0.33 $Y=-0.265 $X2=0.775
+ $Y2=1.55
cc_61 N_VNB_c_3_p N_GCLK_c_918_n 8.26786e-19 $X=9.84 $Y=0 $X2=0.775 $Y2=1.55
cc_62 N_VNB_M1002_b GCLK 0.00790378f $X=-0.33 $Y=-0.265 $X2=0.695 $Y2=2.6
cc_63 N_VNB_M1002_b GCLK 0.0350821f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_64 N_VNB_M1002_b N_VGND_c_939_n 0.0221748f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_65 N_VNB_M1002_b N_VGND_c_940_n 0.0254446f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_66 N_VNB_c_3_p N_VGND_c_940_n 0.00111205f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_67 N_VNB_M1002_b N_VGND_c_942_n 0.00145347f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_68 N_VNB_M1002_b N_VGND_c_943_n 0.00532348f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_69 N_VNB_M1002_b N_VGND_c_944_n 0.0214543f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_70 N_VNB_c_3_p N_VGND_c_944_n 9.36563e-19 $X=9.84 $Y=0 $X2=0 $Y2=0
cc_71 N_VNB_M1002_b N_VGND_c_946_n 0.0214342f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_72 N_VNB_c_3_p N_VGND_c_946_n 8.48483e-19 $X=9.84 $Y=0 $X2=0 $Y2=0
cc_73 N_VNB_M1002_b N_VGND_c_948_n 0.0824567f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_74 N_VNB_c_3_p N_VGND_c_948_n 0.00335859f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_75 N_VNB_M1002_b N_VGND_c_950_n 0.212407f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_76 N_VNB_c_3_p N_VGND_c_950_n 0.00807515f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_77 N_VNB_M1002_b N_VGND_c_952_n 0.0662157f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_78 N_VNB_c_3_p N_VGND_c_952_n 0.00440274f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_79 N_VNB_M1002_b N_VGND_c_954_n 0.00571477f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_80 N_VNB_M1002_b N_VGND_c_955_n 0.187875f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_81 N_VNB_c_3_p N_VGND_c_955_n 1.06653f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_82 N_VPB_M1000_b N_GATE_M1002_g 0.0761689f $X=-0.33 $Y=1.885 $X2=0.695
+ $Y2=1.005
cc_83 N_VPB_M1000_b N_A_231_71#_M1013_g 0.0453476f $X=-0.33 $Y=1.885 $X2=0.695
+ $Y2=2.6
cc_84 N_VPB_M1000_b N_A_231_71#_c_200_n 0.00414357f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_85 N_VPB_M1000_b N_A_231_71#_c_207_n 0.00350272f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_86 N_VPB_M1000_b N_A_231_71#_c_208_n 0.0108959f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_87 N_VPB_M1000_b N_A_231_71#_c_209_n 0.0525353f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_88 N_VPB_M1000_b N_A_231_71#_M1017_g 0.0651597f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_89 N_VPB_M1000_b N_A_239_419#_M1007_g 0.0512017f $X=-0.33 $Y=1.885 $X2=0.775
+ $Y2=1.55
cc_90 N_VPB_M1000_b N_A_239_419#_c_312_n 0.0313488f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_91 N_VPB_M1000_b N_A_239_419#_c_313_n 0.0733867f $X=-0.33 $Y=1.885 $X2=0.775
+ $Y2=2.035
cc_92 N_VPB_M1000_b N_A_239_419#_c_307_n 0.00581433f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_93 N_VPB_M1000_b N_A_239_419#_c_315_n 0.00390726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_94 N_VPB_M1000_b N_A_239_419#_c_316_n 0.0106153f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_95 N_VPB_M1000_b N_A_239_419#_c_317_n 0.00475575f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_96 N_VPB_M1000_b N_A_239_419#_c_318_n 0.0222215f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_97 N_VPB_c_97_p N_A_239_419#_c_318_n 0.0422653f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_98 N_VPB_c_98_p N_A_239_419#_c_318_n 0.00639071f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_99 N_VPB_M1000_b N_A_239_419#_c_321_n 0.00328996f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_100 N_VPB_c_97_p N_A_239_419#_c_321_n 0.00449732f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_101 N_VPB_c_98_p N_A_239_419#_c_321_n 3.87253e-19 $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_102 N_VPB_M1000_b N_A_239_419#_c_308_n 3.93115e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_103 N_VPB_M1000_b N_A_239_419#_c_325_n 0.00797682f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_104 N_VPB_M1000_b N_A_239_419#_c_326_n 0.0128132f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_105 N_VPB_M1000_b N_A_239_419#_c_327_n 0.00263821f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_106 N_VPB_M1000_b N_A_239_419#_c_310_n 0.0197316f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_107 N_VPB_M1000_b N_A_1069_133#_M1014_g 0.0440333f $X=-0.33 $Y=1.885
+ $X2=0.775 $Y2=1.55
cc_108 N_VPB_M1000_b N_A_1069_133#_c_429_n 0.0197618f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_109 N_VPB_M1000_b N_A_1069_133#_c_430_n 0.004738f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_110 N_VPB_M1000_b N_A_1069_133#_c_438_n 0.00181811f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_111 N_VPB_M1000_b N_A_1069_133#_c_439_n 0.00952042f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_112 N_VPB_M1000_b N_A_1069_133#_c_433_n 0.00335443f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_113 N_VPB_M1000_b N_A_1069_133#_M1015_g 0.0561259f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_114 N_VPB_M1000_b N_A_303_311#_c_514_n 0.0216226f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_115 N_VPB_M1000_b N_A_303_311#_c_528_n 0.0213768f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_116 N_VPB_M1000_b N_A_303_311#_c_521_n 0.00994003f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_117 N_VPB_M1000_b N_A_303_311#_M1001_g 0.0643781f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_118 N_VPB_M1000_b N_CLK_c_647_n 0.0336146f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.58
cc_119 N_VPB_M1000_b N_CLK_c_648_n 0.0373698f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_120 N_VPB_M1000_b N_CLK_c_649_n 0.0756043f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_121 N_VPB_M1000_b N_CLK_c_650_n 0.0678298f $X=-0.33 $Y=1.885 $X2=0.695
+ $Y2=1.55
cc_122 N_VPB_M1000_b N_CLK_c_651_n 0.012325f $X=-0.33 $Y=1.885 $X2=0.775
+ $Y2=1.55
cc_123 N_VPB_c_97_p N_CLK_c_651_n 0.0187586f $X=9.84 $Y=4.07 $X2=0.775 $Y2=1.55
cc_124 N_VPB_c_98_p N_CLK_c_651_n 0.00608604f $X=9.84 $Y=4.07 $X2=0.775 $Y2=1.55
cc_125 N_VPB_M1000_b N_CLK_c_654_n 0.215131f $X=-0.33 $Y=1.885 $X2=0.775
+ $Y2=1.55
cc_126 N_VPB_c_97_p N_CLK_c_654_n 0.00977733f $X=9.84 $Y=4.07 $X2=0.775 $Y2=1.55
cc_127 N_VPB_c_98_p N_CLK_c_654_n 6.81527e-19 $X=9.84 $Y=4.07 $X2=0.775 $Y2=1.55
cc_128 N_VPB_M1000_b N_CLK_c_657_n 0.0105354f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_129 N_VPB_M1000_b N_CLK_c_658_n 0.0261719f $X=-0.33 $Y=1.885 $X2=0.775
+ $Y2=1.55
cc_130 N_VPB_M1000_b N_CLK_c_659_n 0.0179002f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_131 N_VPB_M1000_b N_CLK_c_660_n 0.00241086f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_132 N_VPB_M1000_b N_CLK_c_661_n 0.0221264f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_133 N_VPB_M1000_b N_CLK_c_662_n 2.06605e-19 $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_134 N_VPB_M1000_b N_CLK_M1005_g 0.0168621f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_135 N_VPB_M1000_b N_CLK_M1011_g 0.0312102f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_136 N_VPB_M1000_b N_A_1438_171#_M1016_g 0.0617617f $X=-0.33 $Y=1.885
+ $X2=0.695 $Y2=2.6
cc_137 N_VPB_c_97_p N_A_1438_171#_M1016_g 0.0148572f $X=9.84 $Y=4.07 $X2=0.695
+ $Y2=2.6
cc_138 N_VPB_c_98_p N_A_1438_171#_M1016_g 0.00970178f $X=9.84 $Y=4.07 $X2=0.695
+ $Y2=2.6
cc_139 N_VPB_M1000_b N_A_1438_171#_c_750_n 0.00690622f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_140 N_VPB_M1000_b N_VPWR_c_806_n 0.0809155f $X=-0.33 $Y=1.885 $X2=0.775
+ $Y2=2.035
cc_141 N_VPB_M1000_b N_VPWR_c_807_n 0.00939912f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_142 N_VPB_M1000_b N_VPWR_c_808_n 0.00835239f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_143 N_VPB_c_97_p N_VPWR_c_808_n 0.0332587f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_144 N_VPB_c_98_p N_VPWR_c_808_n 0.00157083f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_145 N_VPB_M1000_b N_VPWR_c_811_n 0.0233586f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_146 N_VPB_M1000_b N_VPWR_c_812_n 0.0100233f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_147 N_VPB_c_97_p N_VPWR_c_812_n 0.0705217f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_148 N_VPB_c_98_p N_VPWR_c_812_n 0.00339185f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_149 N_VPB_M1000_b N_VPWR_c_815_n 0.0336273f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_150 N_VPB_M1000_b N_VPWR_c_816_n 0.00800311f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_151 N_VPB_M1000_b N_VPWR_c_817_n 0.010434f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_152 N_VPB_c_97_p N_VPWR_c_817_n 0.0236698f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_153 N_VPB_c_98_p N_VPWR_c_817_n 0.00111205f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_154 N_VPB_M1000_b N_VPWR_c_820_n 0.0033245f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_155 N_VPB_c_97_p N_VPWR_c_820_n 0.0236698f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_156 N_VPB_c_98_p N_VPWR_c_820_n 0.00111205f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_157 N_VPB_M1000_b N_VPWR_c_823_n 0.00399863f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_158 N_VPB_c_97_p N_VPWR_c_823_n 0.137938f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_159 N_VPB_c_98_p N_VPWR_c_823_n 0.00719674f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_160 N_VPB_M1000_b N_VPWR_c_826_n 0.00393018f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_161 N_VPB_M1000_b N_VPWR_c_827_n 0.0118572f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_162 N_VPB_c_97_p N_VPWR_c_827_n 0.203327f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_163 N_VPB_c_98_p N_VPWR_c_827_n 0.00982734f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_164 N_VPB_M1000_b N_VPWR_c_830_n 0.00690303f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_165 N_VPB_M1000_b N_VPWR_c_831_n 0.0284576f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_166 N_VPB_M1000_b N_VPWR_c_832_n 0.0208331f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_167 N_VPB_M1000_b N_VPWR_c_833_n 0.0113673f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_168 N_VPB_M1000_b N_VPWR_c_834_n 0.00408898f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_169 N_VPB_M1000_b N_VPWR_c_835_n 0.111465f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_170 N_VPB_c_97_p N_VPWR_c_835_n 0.0364227f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_171 N_VPB_c_98_p N_VPWR_c_835_n 1.06867f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_172 N_VPB_M1000_b GCLK 0.0816296f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_173 N_VPB_c_97_p GCLK 0.0176346f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_174 N_VPB_c_98_p GCLK 0.00107864f $X=9.84 $Y=4.07 $X2=0 $Y2=0
cc_175 N_VPB_M1000_b GCLK 5.03744e-19 $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_176 N_GATE_M1002_g N_A_231_71#_c_194_n 0.00154721f $X=0.695 $Y=1.005 $X2=9.84
+ $Y2=0
cc_177 N_GATE_M1002_g N_A_231_71#_c_204_n 0.0445345f $X=0.695 $Y=1.005 $X2=0
+ $Y2=0
cc_178 N_GATE_M1002_g N_A_239_419#_M1007_g 0.0674163f $X=0.695 $Y=1.005 $X2=0
+ $Y2=0
cc_179 N_GATE_c_181_p N_A_239_419#_M1007_g 7.51674e-19 $X=0.775 $Y=1.55 $X2=0
+ $Y2=0
cc_180 N_GATE_M1002_g N_A_303_311#_c_514_n 0.00673523f $X=0.695 $Y=1.005 $X2=0
+ $Y2=0
cc_181 N_GATE_c_181_p N_A_303_311#_c_514_n 0.00162143f $X=0.775 $Y=1.55 $X2=0
+ $Y2=0
cc_182 N_GATE_M1002_g N_A_303_311#_c_533_n 0.0013419f $X=0.695 $Y=1.005 $X2=0
+ $Y2=0
cc_183 N_GATE_c_181_p N_A_303_311#_c_533_n 0.00827961f $X=0.775 $Y=1.55 $X2=0
+ $Y2=0
cc_184 N_GATE_M1002_g N_VPWR_c_806_n 0.00969653f $X=0.695 $Y=1.005 $X2=0 $Y2=0
cc_185 N_GATE_M1002_g N_VPWR_c_827_n 0.0156399f $X=0.695 $Y=1.005 $X2=0 $Y2=0
cc_186 N_GATE_M1002_g N_VPWR_c_835_n 0.0142618f $X=0.695 $Y=1.005 $X2=0 $Y2=0
cc_187 N_GATE_M1002_g N_VGND_c_939_n 0.0277882f $X=0.695 $Y=1.005 $X2=0 $Y2=0
cc_188 N_GATE_M1002_g N_VGND_c_946_n 0.0135337f $X=0.695 $Y=1.005 $X2=0 $Y2=0
cc_189 N_GATE_M1002_g N_VGND_c_955_n 0.0161918f $X=0.695 $Y=1.005 $X2=0 $Y2=0
cc_190 N_A_231_71#_c_199_n N_A_239_419#_M1004_g 0.00105329f $X=3.945 $Y=0.87
+ $X2=0 $Y2=0
cc_191 N_A_231_71#_c_200_n N_A_239_419#_M1004_g 0.00212952f $X=3.945 $Y=2.43
+ $X2=0 $Y2=0
cc_192 N_A_231_71#_c_202_n N_A_239_419#_M1004_g 6.26088e-19 $X=3.945 $Y=1.21
+ $X2=0 $Y2=0
cc_193 N_A_231_71#_M1017_g N_A_239_419#_c_313_n 3.73446e-19 $X=2.775 $Y=0.87
+ $X2=0 $Y2=0
cc_194 N_A_231_71#_c_217_p N_A_239_419#_c_307_n 0.0158903f $X=2.725 $Y=1.125
+ $X2=0.24 $Y2=0
cc_195 N_A_231_71#_c_218_p N_A_239_419#_c_307_n 0.0508419f $X=2.805 $Y=1.46
+ $X2=0.24 $Y2=0
cc_196 N_A_231_71#_c_219_p N_A_239_419#_c_307_n 0.0137194f $X=2.805 $Y=1.21
+ $X2=0.24 $Y2=0
cc_197 N_A_231_71#_M1017_g N_A_239_419#_c_307_n 0.0180957f $X=2.775 $Y=0.87
+ $X2=0.24 $Y2=0
cc_198 N_A_231_71#_M1017_g N_A_239_419#_c_315_n 0.0057721f $X=2.775 $Y=0.87
+ $X2=5.04 $Y2=0
cc_199 N_A_231_71#_c_218_p N_A_239_419#_c_316_n 0.0238596f $X=2.805 $Y=1.46
+ $X2=9.84 $Y2=0
cc_200 N_A_231_71#_c_200_n N_A_239_419#_c_316_n 0.0122925f $X=3.945 $Y=2.43
+ $X2=9.84 $Y2=0
cc_201 N_A_231_71#_M1017_g N_A_239_419#_c_316_n 0.046123f $X=2.775 $Y=0.87
+ $X2=9.84 $Y2=0
cc_202 N_A_231_71#_c_207_n N_A_239_419#_c_317_n 0.0156852f $X=4.07 $Y=3.11 $X2=0
+ $Y2=0
cc_203 N_A_231_71#_M1017_g N_A_239_419#_c_317_n 7.58866e-19 $X=2.775 $Y=0.87
+ $X2=0 $Y2=0
cc_204 N_A_231_71#_c_207_n N_A_239_419#_c_318_n 0.0160487f $X=4.07 $Y=3.11 $X2=0
+ $Y2=0
cc_205 N_A_231_71#_c_208_n N_A_239_419#_c_318_n 0.0741877f $X=5.01 $Y=3.13 $X2=0
+ $Y2=0
cc_206 N_A_231_71#_c_209_n N_A_239_419#_c_318_n 0.00450736f $X=5.01 $Y=3.13
+ $X2=0 $Y2=0
cc_207 N_A_231_71#_M1013_g N_A_239_419#_c_325_n 0.00250036f $X=4.885 $Y=2.495
+ $X2=0 $Y2=0
cc_208 N_A_231_71#_M1013_g N_A_239_419#_c_326_n 0.00670468f $X=4.885 $Y=2.495
+ $X2=0 $Y2=0
cc_209 N_A_231_71#_c_208_n N_A_239_419#_c_326_n 0.0166225f $X=5.01 $Y=3.13 $X2=0
+ $Y2=0
cc_210 N_A_231_71#_c_209_n N_A_239_419#_c_326_n 0.00646424f $X=5.01 $Y=3.13
+ $X2=0 $Y2=0
cc_211 N_A_231_71#_c_196_n N_A_239_419#_c_309_n 0.0173878f $X=2.64 $Y=0.45 $X2=0
+ $Y2=0
cc_212 N_A_231_71#_M1013_g N_A_239_419#_c_353_n 0.00322555f $X=4.885 $Y=2.495
+ $X2=0 $Y2=0
cc_213 N_A_231_71#_M1013_g N_A_239_419#_c_310_n 0.0385198f $X=4.885 $Y=2.495
+ $X2=0 $Y2=0
cc_214 N_A_231_71#_M1013_g N_A_239_419#_c_355_n 0.00234262f $X=4.885 $Y=2.495
+ $X2=0 $Y2=0
cc_215 N_A_231_71#_M1013_g N_A_1069_133#_M1014_g 0.0450374f $X=4.885 $Y=2.495
+ $X2=0 $Y2=0
cc_216 N_A_231_71#_c_194_n N_A_303_311#_c_506_n 0.0216006f $X=1.66 $Y=0.52 $X2=0
+ $Y2=0
cc_217 N_A_231_71#_c_196_n N_A_303_311#_c_506_n 0.0126221f $X=2.64 $Y=0.45 $X2=0
+ $Y2=0
cc_218 N_A_231_71#_c_217_p N_A_303_311#_c_506_n 0.00111324f $X=2.725 $Y=1.125
+ $X2=0 $Y2=0
cc_219 N_A_231_71#_c_201_n N_A_303_311#_c_506_n 0.00282797f $X=1.865 $Y=0.517
+ $X2=0 $Y2=0
cc_220 N_A_231_71#_M1017_g N_A_303_311#_c_506_n 0.0358705f $X=2.775 $Y=0.87
+ $X2=0 $Y2=0
cc_221 N_A_231_71#_c_204_n N_A_303_311#_c_506_n 0.0150583f $X=1.49 $Y=0.685
+ $X2=0 $Y2=0
cc_222 N_A_231_71#_c_196_n N_A_303_311#_c_507_n 0.00716755f $X=2.64 $Y=0.45
+ $X2=0 $Y2=0
cc_223 N_A_231_71#_c_199_n N_A_303_311#_c_507_n 0.00167765f $X=3.945 $Y=0.87
+ $X2=0 $Y2=0
cc_224 N_A_231_71#_M1017_g N_A_303_311#_c_507_n 0.0341663f $X=2.775 $Y=0.87
+ $X2=0 $Y2=0
cc_225 N_A_231_71#_c_204_n N_A_303_311#_c_514_n 0.0133095f $X=1.49 $Y=0.685
+ $X2=0 $Y2=0
cc_226 N_A_231_71#_c_192_n N_A_303_311#_c_515_n 0.0124004f $X=1.713 $Y=0.517
+ $X2=0 $Y2=0
cc_227 N_A_231_71#_c_194_n N_A_303_311#_c_515_n 0.00290424f $X=1.66 $Y=0.52
+ $X2=0 $Y2=0
cc_228 N_A_231_71#_c_196_n N_A_303_311#_c_515_n 0.00516417f $X=2.64 $Y=0.45
+ $X2=0 $Y2=0
cc_229 N_A_231_71#_c_204_n N_A_303_311#_c_515_n 0.0259809f $X=1.49 $Y=0.685
+ $X2=0 $Y2=0
cc_230 N_A_231_71#_M1017_g N_A_303_311#_c_528_n 0.00120708f $X=2.775 $Y=0.87
+ $X2=9.84 $Y2=0
cc_231 N_A_231_71#_c_199_n N_A_303_311#_c_516_n 0.0214295f $X=3.945 $Y=0.87
+ $X2=0 $Y2=0
cc_232 N_A_231_71#_c_202_n N_A_303_311#_c_516_n 0.0039395f $X=3.945 $Y=1.21
+ $X2=0 $Y2=0
cc_233 N_A_231_71#_c_204_n N_A_303_311#_c_533_n 5.99356e-19 $X=1.49 $Y=0.685
+ $X2=0 $Y2=0
cc_234 N_A_231_71#_c_200_n N_A_303_311#_c_520_n 0.00396656f $X=3.945 $Y=2.43
+ $X2=0 $Y2=0
cc_235 N_A_231_71#_c_202_n N_A_303_311#_c_520_n 0.00618616f $X=3.945 $Y=1.21
+ $X2=0 $Y2=0
cc_236 N_A_231_71#_M1013_g N_A_303_311#_c_555_n 0.0089084f $X=4.885 $Y=2.495
+ $X2=0 $Y2=0
cc_237 N_A_231_71#_c_208_n N_A_303_311#_c_555_n 0.0119223f $X=5.01 $Y=3.13 $X2=0
+ $Y2=0
cc_238 N_A_231_71#_c_209_n N_A_303_311#_c_555_n 0.0025817f $X=5.01 $Y=3.13 $X2=0
+ $Y2=0
cc_239 N_A_231_71#_M1013_g N_A_303_311#_c_521_n 0.00170117f $X=4.885 $Y=2.495
+ $X2=0 $Y2=0
cc_240 N_A_231_71#_c_200_n N_A_303_311#_c_521_n 0.0654634f $X=3.945 $Y=2.43
+ $X2=0 $Y2=0
cc_241 N_A_231_71#_c_200_n N_CLK_c_647_n 0.00115897f $X=3.945 $Y=2.43 $X2=0
+ $Y2=0
cc_242 N_A_231_71#_c_207_n N_CLK_c_647_n 0.00135212f $X=4.07 $Y=3.11 $X2=0 $Y2=0
cc_243 N_A_231_71#_M1013_g N_CLK_c_648_n 0.0213012f $X=4.885 $Y=2.495 $X2=0
+ $Y2=0
cc_244 N_A_231_71#_c_200_n N_CLK_c_648_n 0.0185005f $X=3.945 $Y=2.43 $X2=0 $Y2=0
cc_245 N_A_231_71#_c_200_n N_CLK_c_649_n 0.0128667f $X=3.945 $Y=2.43 $X2=0 $Y2=0
cc_246 N_A_231_71#_c_208_n N_CLK_c_649_n 0.0164123f $X=5.01 $Y=3.13 $X2=0 $Y2=0
cc_247 N_A_231_71#_c_209_n N_CLK_c_649_n 0.022375f $X=5.01 $Y=3.13 $X2=0 $Y2=0
cc_248 N_A_231_71#_c_208_n N_CLK_c_650_n 0.00123896f $X=5.01 $Y=3.13 $X2=0 $Y2=0
cc_249 N_A_231_71#_c_209_n N_CLK_c_650_n 0.0431406f $X=5.01 $Y=3.13 $X2=0 $Y2=0
cc_250 N_A_231_71#_c_218_p CLK 0.0192413f $X=2.805 $Y=1.46 $X2=0 $Y2=0
cc_251 N_A_231_71#_c_198_n CLK 0.0244185f $X=3.82 $Y=1.21 $X2=0 $Y2=0
cc_252 N_A_231_71#_c_200_n CLK 0.038989f $X=3.945 $Y=2.43 $X2=0 $Y2=0
cc_253 N_A_231_71#_M1017_g CLK 0.0020333f $X=2.775 $Y=0.87 $X2=0 $Y2=0
cc_254 N_A_231_71#_c_217_p N_CLK_M1005_g 7.08404e-19 $X=2.725 $Y=1.125 $X2=0
+ $Y2=0
cc_255 N_A_231_71#_c_218_p N_CLK_M1005_g 0.00305625f $X=2.805 $Y=1.46 $X2=0
+ $Y2=0
cc_256 N_A_231_71#_c_198_n N_CLK_M1005_g 0.0373744f $X=3.82 $Y=1.21 $X2=0 $Y2=0
cc_257 N_A_231_71#_c_199_n N_CLK_M1005_g 0.00254632f $X=3.945 $Y=0.87 $X2=0
+ $Y2=0
cc_258 N_A_231_71#_c_200_n N_CLK_M1005_g 0.0260173f $X=3.945 $Y=2.43 $X2=0 $Y2=0
cc_259 N_A_231_71#_M1017_g N_CLK_M1005_g 0.0783912f $X=2.775 $Y=0.87 $X2=0 $Y2=0
cc_260 N_A_231_71#_M1017_g N_VPWR_c_807_n 0.0191226f $X=2.775 $Y=0.87 $X2=0
+ $Y2=0
cc_261 N_A_231_71#_M1017_g N_VPWR_c_831_n 0.00260124f $X=2.775 $Y=0.87 $X2=0
+ $Y2=0
cc_262 N_A_231_71#_M1017_g N_VPWR_c_832_n 0.011461f $X=2.775 $Y=0.87 $X2=0 $Y2=0
cc_263 N_A_231_71#_c_207_n N_VPWR_c_835_n 0.00150099f $X=4.07 $Y=3.11 $X2=0
+ $Y2=0
cc_264 N_A_231_71#_c_208_n N_VPWR_c_835_n 0.00678346f $X=5.01 $Y=3.13 $X2=0
+ $Y2=0
cc_265 N_A_231_71#_M1017_g N_VPWR_c_835_n 0.0140641f $X=2.775 $Y=0.87 $X2=0
+ $Y2=0
cc_266 N_A_231_71#_c_194_n N_VGND_c_939_n 5.80438e-19 $X=1.66 $Y=0.52 $X2=0
+ $Y2=0
cc_267 N_A_231_71#_c_192_n N_VGND_c_946_n 0.00719691f $X=1.713 $Y=0.517 $X2=0
+ $Y2=0
cc_268 N_A_231_71#_c_194_n N_VGND_c_946_n 0.00133831f $X=1.66 $Y=0.52 $X2=0
+ $Y2=0
cc_269 N_A_231_71#_c_196_n N_VGND_c_952_n 0.0126369f $X=2.64 $Y=0.45 $X2=0 $Y2=0
cc_270 N_A_231_71#_c_217_p N_VGND_c_952_n 0.0296816f $X=2.725 $Y=1.125 $X2=0
+ $Y2=0
cc_271 N_A_231_71#_c_198_n N_VGND_c_952_n 0.029749f $X=3.82 $Y=1.21 $X2=0 $Y2=0
cc_272 N_A_231_71#_c_199_n N_VGND_c_952_n 0.00600645f $X=3.945 $Y=0.87 $X2=0
+ $Y2=0
cc_273 N_A_231_71#_M1017_g N_VGND_c_952_n 0.00987062f $X=2.775 $Y=0.87 $X2=0
+ $Y2=0
cc_274 N_A_231_71#_c_192_n N_VGND_c_955_n 0.0498777f $X=1.713 $Y=0.517 $X2=0
+ $Y2=0
cc_275 N_A_231_71#_c_194_n N_VGND_c_955_n 0.0110697f $X=1.66 $Y=0.52 $X2=0 $Y2=0
cc_276 N_A_231_71#_c_196_n N_VGND_c_955_n 0.0366193f $X=2.64 $Y=0.45 $X2=0 $Y2=0
cc_277 N_A_231_71#_c_217_p N_VGND_c_955_n 0.0145567f $X=2.725 $Y=1.125 $X2=0
+ $Y2=0
cc_278 N_A_231_71#_c_198_n N_VGND_c_955_n 0.00679347f $X=3.82 $Y=1.21 $X2=0
+ $Y2=0
cc_279 N_A_231_71#_c_199_n N_VGND_c_955_n 0.00978915f $X=3.945 $Y=0.87 $X2=0
+ $Y2=0
cc_280 N_A_231_71#_c_201_n N_VGND_c_955_n 0.0107132f $X=1.865 $Y=0.517 $X2=0
+ $Y2=0
cc_281 N_A_231_71#_c_219_p N_VGND_c_955_n 0.00545045f $X=2.805 $Y=1.21 $X2=0
+ $Y2=0
cc_282 N_A_231_71#_M1017_g N_VGND_c_955_n 0.00920703f $X=2.775 $Y=0.87 $X2=0
+ $Y2=0
cc_283 N_A_239_419#_M1004_g N_A_1069_133#_M1009_g 0.0497875f $X=4.885 $Y=1.005
+ $X2=0 $Y2=0
cc_284 N_A_239_419#_c_325_n N_A_1069_133#_M1014_g 0.0037708f $X=5.22 $Y=2.425
+ $X2=0 $Y2=0
cc_285 N_A_239_419#_c_326_n N_A_1069_133#_M1014_g 0.0152602f $X=5.43 $Y=3.385
+ $X2=0 $Y2=0
cc_286 N_A_239_419#_c_355_n N_A_1069_133#_M1014_g 0.0146326f $X=5.43 $Y=2.51
+ $X2=0 $Y2=0
cc_287 N_A_239_419#_M1004_g N_A_1069_133#_c_447_n 5.37106e-19 $X=4.885 $Y=1.005
+ $X2=0 $Y2=0
cc_288 N_A_239_419#_c_308_n N_A_1069_133#_c_447_n 0.0172818f $X=5.22 $Y=1.945
+ $X2=0 $Y2=0
cc_289 N_A_239_419#_c_310_n N_A_1069_133#_c_447_n 3.24891e-19 $X=5.14 $Y=1.78
+ $X2=0 $Y2=0
cc_290 N_A_239_419#_M1004_g N_A_1069_133#_c_429_n 0.0112001f $X=4.885 $Y=1.005
+ $X2=0 $Y2=0
cc_291 N_A_239_419#_c_308_n N_A_1069_133#_c_429_n 9.92402e-19 $X=5.22 $Y=1.945
+ $X2=0 $Y2=0
cc_292 N_A_239_419#_c_325_n N_A_1069_133#_c_429_n 0.00344043f $X=5.22 $Y=2.425
+ $X2=0 $Y2=0
cc_293 N_A_239_419#_c_310_n N_A_1069_133#_c_429_n 0.0209751f $X=5.14 $Y=1.78
+ $X2=0 $Y2=0
cc_294 N_A_239_419#_c_308_n N_A_1069_133#_c_438_n 0.00494204f $X=5.22 $Y=1.945
+ $X2=4.08 $Y2=0
cc_295 N_A_239_419#_c_325_n N_A_1069_133#_c_438_n 0.00950131f $X=5.22 $Y=2.425
+ $X2=4.08 $Y2=0
cc_296 N_A_239_419#_c_307_n N_A_303_311#_c_506_n 0.00721122f $X=2.372 $Y=2.145
+ $X2=0 $Y2=0
cc_297 N_A_239_419#_c_309_n N_A_303_311#_c_506_n 0.00587198f $X=2.385 $Y=0.87
+ $X2=0 $Y2=0
cc_298 N_A_239_419#_M1004_g N_A_303_311#_c_510_n 0.0339362f $X=4.885 $Y=1.005
+ $X2=9.84 $Y2=0
cc_299 N_A_239_419#_M1007_g N_A_303_311#_c_514_n 0.0133095f $X=1.445 $Y=2.6
+ $X2=0 $Y2=0
cc_300 N_A_239_419#_c_307_n N_A_303_311#_c_515_n 0.0271464f $X=2.372 $Y=2.145
+ $X2=0 $Y2=0
cc_301 N_A_239_419#_c_309_n N_A_303_311#_c_515_n 0.0163217f $X=2.385 $Y=0.87
+ $X2=0 $Y2=0
cc_302 N_A_239_419#_M1007_g N_A_303_311#_c_528_n 0.0472475f $X=1.445 $Y=2.6
+ $X2=9.84 $Y2=0
cc_303 N_A_239_419#_c_312_n N_A_303_311#_c_528_n 0.0260606f $X=2.275 $Y=3.275
+ $X2=9.84 $Y2=0
cc_304 N_A_239_419#_c_313_n N_A_303_311#_c_528_n 0.00410617f $X=1.7 $Y=3.3
+ $X2=9.84 $Y2=0
cc_305 N_A_239_419#_c_307_n N_A_303_311#_c_528_n 0.0148781f $X=2.372 $Y=2.145
+ $X2=9.84 $Y2=0
cc_306 N_A_239_419#_c_315_n N_A_303_311#_c_528_n 0.0382585f $X=2.385 $Y=2.43
+ $X2=9.84 $Y2=0
cc_307 N_A_239_419#_c_327_n N_A_303_311#_c_528_n 0.0106912f $X=2.385 $Y=2.23
+ $X2=9.84 $Y2=0
cc_308 N_A_239_419#_M1004_g N_A_303_311#_c_516_n 0.0155948f $X=4.885 $Y=1.005
+ $X2=0 $Y2=0
cc_309 N_A_239_419#_M1004_g N_A_303_311#_c_517_n 0.0295437f $X=4.885 $Y=1.005
+ $X2=0 $Y2=0
cc_310 N_A_239_419#_c_308_n N_A_303_311#_c_517_n 0.010157f $X=5.22 $Y=1.945
+ $X2=0 $Y2=0
cc_311 N_A_239_419#_c_353_n N_A_303_311#_c_517_n 0.0220125f $X=5.14 $Y=1.78
+ $X2=0 $Y2=0
cc_312 N_A_239_419#_c_310_n N_A_303_311#_c_517_n 0.00110502f $X=5.14 $Y=1.78
+ $X2=0 $Y2=0
cc_313 N_A_239_419#_M1007_g N_A_303_311#_c_533_n 5.99356e-19 $X=1.445 $Y=2.6
+ $X2=0 $Y2=0
cc_314 N_A_239_419#_c_307_n N_A_303_311#_c_533_n 0.0258793f $X=2.372 $Y=2.145
+ $X2=0 $Y2=0
cc_315 N_A_239_419#_M1004_g N_A_303_311#_c_520_n 0.004799f $X=4.885 $Y=1.005
+ $X2=0 $Y2=0
cc_316 N_A_239_419#_c_355_n N_A_303_311#_c_555_n 0.00548082f $X=5.43 $Y=2.51
+ $X2=0 $Y2=0
cc_317 N_A_239_419#_M1004_g N_A_303_311#_c_521_n 0.0180491f $X=4.885 $Y=1.005
+ $X2=0 $Y2=0
cc_318 N_A_239_419#_c_325_n N_A_303_311#_c_521_n 0.0105484f $X=5.22 $Y=2.425
+ $X2=0 $Y2=0
cc_319 N_A_239_419#_c_353_n N_A_303_311#_c_521_n 0.0259146f $X=5.14 $Y=1.78
+ $X2=0 $Y2=0
cc_320 N_A_239_419#_c_316_n N_CLK_c_647_n 0.0144999f $X=3.52 $Y=2.23 $X2=0 $Y2=0
cc_321 N_A_239_419#_c_317_n N_CLK_c_647_n 0.0357822f $X=3.605 $Y=3.385 $X2=0
+ $Y2=0
cc_322 N_A_239_419#_c_318_n N_CLK_c_647_n 0.00450678f $X=5.345 $Y=3.47 $X2=0
+ $Y2=0
cc_323 N_A_239_419#_c_317_n N_CLK_c_649_n 0.00479023f $X=3.605 $Y=3.385 $X2=0
+ $Y2=0
cc_324 N_A_239_419#_c_318_n N_CLK_c_649_n 0.00932609f $X=5.345 $Y=3.47 $X2=0
+ $Y2=0
cc_325 N_A_239_419#_c_318_n N_CLK_c_650_n 0.0215375f $X=5.345 $Y=3.47 $X2=0
+ $Y2=0
cc_326 N_A_239_419#_c_318_n N_CLK_c_651_n 0.00311696f $X=5.345 $Y=3.47 $X2=0
+ $Y2=0
cc_327 N_A_239_419#_c_316_n N_CLK_c_657_n 0.0111111f $X=3.52 $Y=2.23 $X2=0 $Y2=0
cc_328 N_A_239_419#_c_318_n N_CLK_c_658_n 0.00751504f $X=5.345 $Y=3.47 $X2=0
+ $Y2=0
cc_329 N_A_239_419#_c_326_n N_CLK_c_658_n 0.00582586f $X=5.43 $Y=3.385 $X2=0
+ $Y2=0
cc_330 N_A_239_419#_c_316_n CLK 0.0258168f $X=3.52 $Y=2.23 $X2=0 $Y2=0
cc_331 N_A_239_419#_c_316_n N_VPWR_M1018_d 0.00176461f $X=3.52 $Y=2.23 $X2=0
+ $Y2=0
cc_332 N_A_239_419#_c_312_n N_VPWR_c_807_n 0.00913655f $X=2.275 $Y=3.275 $X2=0
+ $Y2=0
cc_333 N_A_239_419#_c_315_n N_VPWR_c_807_n 0.0128292f $X=2.385 $Y=2.43 $X2=0
+ $Y2=0
cc_334 N_A_239_419#_c_316_n N_VPWR_c_807_n 0.0170777f $X=3.52 $Y=2.23 $X2=0
+ $Y2=0
cc_335 N_A_239_419#_c_317_n N_VPWR_c_807_n 0.0605163f $X=3.605 $Y=3.385 $X2=0
+ $Y2=0
cc_336 N_A_239_419#_c_321_n N_VPWR_c_807_n 0.004906f $X=3.69 $Y=3.47 $X2=0 $Y2=0
cc_337 N_A_239_419#_c_318_n N_VPWR_c_808_n 0.00771967f $X=5.345 $Y=3.47 $X2=4.08
+ $Y2=0.058
cc_338 N_A_239_419#_c_318_n N_VPWR_c_811_n 0.00297101f $X=5.345 $Y=3.47 $X2=9.84
+ $Y2=0
cc_339 N_A_239_419#_c_326_n N_VPWR_c_811_n 0.0391479f $X=5.43 $Y=3.385 $X2=9.84
+ $Y2=0
cc_340 N_A_239_419#_c_355_n N_VPWR_c_811_n 0.00800985f $X=5.43 $Y=2.51 $X2=9.84
+ $Y2=0
cc_341 N_A_239_419#_c_313_n N_VPWR_c_830_n 6.18412e-19 $X=1.7 $Y=3.3 $X2=0 $Y2=0
cc_342 N_A_239_419#_c_312_n N_VPWR_c_831_n 0.085387f $X=2.275 $Y=3.275 $X2=0
+ $Y2=0
cc_343 N_A_239_419#_c_313_n N_VPWR_c_831_n 0.0138098f $X=1.7 $Y=3.3 $X2=0 $Y2=0
cc_344 N_A_239_419#_c_321_n N_VPWR_c_832_n 0.00726573f $X=3.69 $Y=3.47 $X2=0
+ $Y2=0
cc_345 N_A_239_419#_c_312_n N_VPWR_c_835_n 0.0413643f $X=2.275 $Y=3.275 $X2=0
+ $Y2=0
cc_346 N_A_239_419#_c_313_n N_VPWR_c_835_n 0.0154534f $X=1.7 $Y=3.3 $X2=0 $Y2=0
cc_347 N_A_239_419#_c_318_n N_VPWR_c_835_n 0.0865538f $X=5.345 $Y=3.47 $X2=0
+ $Y2=0
cc_348 N_A_239_419#_c_321_n N_VPWR_c_835_n 0.0109394f $X=3.69 $Y=3.47 $X2=0
+ $Y2=0
cc_349 N_A_239_419#_c_325_n A_1027_457# 2.83863e-19 $X=5.22 $Y=2.425 $X2=0 $Y2=0
cc_350 N_A_239_419#_c_355_n A_1027_457# 0.00392031f $X=5.43 $Y=2.51 $X2=0 $Y2=0
cc_351 N_A_239_419#_M1004_g N_VGND_c_942_n 0.00109843f $X=4.885 $Y=1.005 $X2=0
+ $Y2=0
cc_352 N_A_239_419#_M1004_g N_VGND_c_948_n 0.0037848f $X=4.885 $Y=1.005 $X2=0
+ $Y2=0
cc_353 N_A_239_419#_M1004_g N_VGND_c_955_n 0.00881496f $X=4.885 $Y=1.005 $X2=0
+ $Y2=0
cc_354 N_A_239_419#_c_309_n N_VGND_c_955_n 0.00843397f $X=2.385 $Y=0.87 $X2=0
+ $Y2=0
cc_355 N_A_1069_133#_M1009_g N_A_303_311#_c_510_n 0.0324969f $X=5.595 $Y=1.005
+ $X2=9.84 $Y2=0
cc_356 N_A_1069_133#_M1009_g N_A_303_311#_c_516_n 0.00161875f $X=5.595 $Y=1.005
+ $X2=0 $Y2=0
cc_357 N_A_1069_133#_M1009_g N_A_303_311#_c_517_n 0.0242148f $X=5.595 $Y=1.005
+ $X2=0 $Y2=0
cc_358 N_A_1069_133#_c_447_n N_A_303_311#_c_517_n 0.0306372f $X=5.68 $Y=1.62
+ $X2=0 $Y2=0
cc_359 N_A_1069_133#_c_429_n N_A_303_311#_c_517_n 0.00714518f $X=5.68 $Y=1.62
+ $X2=0 $Y2=0
cc_360 N_A_1069_133#_c_430_n N_A_303_311#_c_517_n 0.0324239f $X=6.66 $Y=1.98
+ $X2=0 $Y2=0
cc_361 N_A_1069_133#_c_433_n N_A_303_311#_c_517_n 0.0236017f $X=6.795 $Y=1.72
+ $X2=0 $Y2=0
cc_362 N_A_1069_133#_M1014_g N_A_303_311#_c_555_n 3.32419e-19 $X=5.595 $Y=2.495
+ $X2=0 $Y2=0
cc_363 N_A_1069_133#_M1009_g N_A_303_311#_c_592_n 6.91395e-19 $X=5.595 $Y=1.005
+ $X2=0 $Y2=0
cc_364 N_A_1069_133#_c_431_n N_A_303_311#_c_592_n 0.0236017f $X=6.765 $Y=1.005
+ $X2=0 $Y2=0
cc_365 N_A_1069_133#_c_431_n N_A_303_311#_c_522_n 0.017839f $X=6.765 $Y=1.005
+ $X2=0 $Y2=0
cc_366 N_A_1069_133#_M1009_g N_A_303_311#_c_524_n 0.0357709f $X=5.595 $Y=1.005
+ $X2=0 $Y2=0
cc_367 N_A_1069_133#_c_431_n N_A_303_311#_c_524_n 0.00584031f $X=6.765 $Y=1.005
+ $X2=0 $Y2=0
cc_368 N_A_1069_133#_c_447_n N_A_303_311#_M1001_g 0.0020688f $X=5.68 $Y=1.62
+ $X2=0 $Y2=0
cc_369 N_A_1069_133#_c_429_n N_A_303_311#_M1001_g 0.0357709f $X=5.68 $Y=1.62
+ $X2=0 $Y2=0
cc_370 N_A_1069_133#_c_430_n N_A_303_311#_M1001_g 0.0491847f $X=6.66 $Y=1.98
+ $X2=0 $Y2=0
cc_371 N_A_1069_133#_c_431_n N_A_303_311#_M1001_g 0.0237744f $X=6.765 $Y=1.005
+ $X2=0 $Y2=0
cc_372 N_A_1069_133#_c_433_n N_A_303_311#_M1001_g 0.0122453f $X=6.795 $Y=1.72
+ $X2=0 $Y2=0
cc_373 N_A_1069_133#_c_439_n N_CLK_c_654_n 0.00643251f $X=6.765 $Y=2.495
+ $X2=0.24 $Y2=0
cc_374 N_A_1069_133#_M1015_g N_CLK_c_654_n 0.0344327f $X=7.705 $Y=1.065 $X2=0.24
+ $Y2=0
cc_375 N_A_1069_133#_M1014_g N_CLK_c_658_n 0.0129286f $X=5.595 $Y=2.495 $X2=0
+ $Y2=0
cc_376 N_A_1069_133#_M1015_g N_CLK_c_698_n 0.00112559f $X=7.705 $Y=1.065 $X2=0
+ $Y2=0
cc_377 N_A_1069_133#_c_478_p N_CLK_M1011_g 2.36295e-19 $X=7.62 $Y=1.55 $X2=0
+ $Y2=0
cc_378 N_A_1069_133#_M1015_g N_CLK_M1011_g 0.0754254f $X=7.705 $Y=1.065 $X2=0
+ $Y2=0
cc_379 N_A_1069_133#_c_431_n N_A_1438_171#_c_748_n 0.0238595f $X=6.765 $Y=1.005
+ $X2=0 $Y2=0
cc_380 N_A_1069_133#_c_432_n N_A_1438_171#_c_748_n 0.0119322f $X=7.455 $Y=1.72
+ $X2=0 $Y2=0
cc_381 N_A_1069_133#_c_478_p N_A_1438_171#_c_748_n 0.0261514f $X=7.62 $Y=1.55
+ $X2=0 $Y2=0
cc_382 N_A_1069_133#_M1015_g N_A_1438_171#_c_748_n 0.0366962f $X=7.705 $Y=1.065
+ $X2=0 $Y2=0
cc_383 N_A_1069_133#_M1015_g N_A_1438_171#_c_749_n 0.0034635f $X=7.705 $Y=1.065
+ $X2=0 $Y2=0
cc_384 N_A_1069_133#_c_478_p N_A_1438_171#_c_750_n 0.0383515f $X=7.62 $Y=1.55
+ $X2=0 $Y2=0
cc_385 N_A_1069_133#_M1015_g N_A_1438_171#_c_750_n 0.00955406f $X=7.705 $Y=1.065
+ $X2=0 $Y2=0
cc_386 N_A_1069_133#_c_478_p N_A_1438_171#_c_751_n 0.0135702f $X=7.62 $Y=1.55
+ $X2=9.84 $Y2=0
cc_387 N_A_1069_133#_M1015_g N_A_1438_171#_c_751_n 0.00179803f $X=7.705 $Y=1.065
+ $X2=9.84 $Y2=0
cc_388 N_A_1069_133#_M1014_g N_VPWR_c_808_n 0.00106781f $X=5.595 $Y=2.495
+ $X2=4.08 $Y2=0.058
cc_389 N_A_1069_133#_M1014_g N_VPWR_c_811_n 0.0133239f $X=5.595 $Y=2.495
+ $X2=9.84 $Y2=0
cc_390 N_A_1069_133#_c_430_n N_VPWR_c_811_n 0.0154662f $X=6.66 $Y=1.98 $X2=9.84
+ $Y2=0
cc_391 N_A_1069_133#_c_438_n N_VPWR_c_811_n 0.00145814f $X=5.845 $Y=1.98
+ $X2=9.84 $Y2=0
cc_392 N_A_1069_133#_c_439_n N_VPWR_c_815_n 0.0297913f $X=6.765 $Y=2.495 $X2=0
+ $Y2=0
cc_393 N_A_1069_133#_c_432_n N_VPWR_c_815_n 0.0125215f $X=7.455 $Y=1.72 $X2=0
+ $Y2=0
cc_394 N_A_1069_133#_c_478_p N_VPWR_c_815_n 0.00194478f $X=7.62 $Y=1.55 $X2=0
+ $Y2=0
cc_395 N_A_1069_133#_M1015_g N_VPWR_c_815_n 0.0286984f $X=7.705 $Y=1.065 $X2=0
+ $Y2=0
cc_396 N_A_1069_133#_M1015_g N_VPWR_c_823_n 0.00454598f $X=7.705 $Y=1.065 $X2=0
+ $Y2=0
cc_397 N_A_1069_133#_M1014_g N_VPWR_c_835_n 9.50176e-19 $X=5.595 $Y=2.495 $X2=0
+ $Y2=0
cc_398 N_A_1069_133#_M1015_g N_VPWR_c_835_n 0.00251212f $X=7.705 $Y=1.065 $X2=0
+ $Y2=0
cc_399 N_A_1069_133#_M1009_g N_VGND_c_942_n 0.0108286f $X=5.595 $Y=1.005 $X2=0
+ $Y2=0
cc_400 N_A_1069_133#_M1009_g N_VGND_c_948_n 0.00587618f $X=5.595 $Y=1.005 $X2=0
+ $Y2=0
cc_401 N_A_1069_133#_M1015_g N_VGND_c_950_n 0.0147248f $X=7.705 $Y=1.065 $X2=0
+ $Y2=0
cc_402 N_A_1069_133#_M1009_g N_VGND_c_955_n 0.00879005f $X=5.595 $Y=1.005 $X2=0
+ $Y2=0
cc_403 N_A_1069_133#_c_431_n N_VGND_c_955_n 0.00289736f $X=6.765 $Y=1.005 $X2=0
+ $Y2=0
cc_404 N_A_1069_133#_M1015_g N_VGND_c_955_n 0.016429f $X=7.705 $Y=1.065 $X2=0
+ $Y2=0
cc_405 N_A_303_311#_c_521_n N_CLK_c_648_n 0.00398333f $X=4.517 $Y=2.33 $X2=0
+ $Y2=0
cc_406 N_A_303_311#_c_555_n N_CLK_c_649_n 0.00398333f $X=4.495 $Y=2.495 $X2=0
+ $Y2=0
cc_407 N_A_303_311#_M1001_g N_CLK_c_654_n 0.0147455f $X=6.375 $Y=1.005 $X2=0.24
+ $Y2=0
cc_408 N_A_303_311#_c_507_n N_CLK_M1005_g 0.0324429f $X=4.095 $Y=0.245 $X2=0
+ $Y2=0
cc_409 N_A_303_311#_c_512_n N_CLK_M1005_g 0.00221725f $X=4.425 $Y=0.38 $X2=0
+ $Y2=0
cc_410 N_A_303_311#_c_516_n N_CLK_M1005_g 0.00389537f $X=4.495 $Y=1.005 $X2=0
+ $Y2=0
cc_411 N_A_303_311#_c_520_n N_CLK_M1005_g 6.43661e-19 $X=4.517 $Y=1.28 $X2=0
+ $Y2=0
cc_412 N_A_303_311#_M1001_g N_VPWR_c_811_n 0.0189496f $X=6.375 $Y=1.005 $X2=9.84
+ $Y2=0
cc_413 N_A_303_311#_M1001_g N_VPWR_c_812_n 0.00374542f $X=6.375 $Y=1.005 $X2=0
+ $Y2=0
cc_414 N_A_303_311#_M1001_g N_VPWR_c_815_n 0.0053996f $X=6.375 $Y=1.005 $X2=0
+ $Y2=0
cc_415 N_A_303_311#_M1001_g N_VPWR_c_835_n 0.00264801f $X=6.375 $Y=1.005 $X2=0
+ $Y2=0
cc_416 N_A_303_311#_c_517_n N_VGND_M1009_d 0.00173723f $X=6.125 $Y=1.28 $X2=0
+ $Y2=0
cc_417 N_A_303_311#_c_510_n N_VGND_c_940_n 0.015523f $X=6.125 $Y=0.38 $X2=9.84
+ $Y2=0
cc_418 N_A_303_311#_c_522_n N_VGND_c_940_n 0.017883f $X=6.745 $Y=0.52 $X2=9.84
+ $Y2=0
cc_419 N_A_303_311#_c_524_n N_VGND_c_940_n 0.00836226f $X=6.375 $Y=0.685
+ $X2=9.84 $Y2=0
cc_420 N_A_303_311#_c_517_n N_VGND_c_942_n 0.0167644f $X=6.125 $Y=1.28 $X2=0
+ $Y2=0
cc_421 N_A_303_311#_c_592_n N_VGND_c_942_n 0.02528f $X=6.307 $Y=1.195 $X2=0
+ $Y2=0
cc_422 N_A_303_311#_c_522_n N_VGND_c_942_n 0.00343497f $X=6.745 $Y=0.52 $X2=0
+ $Y2=0
cc_423 N_A_303_311#_c_524_n N_VGND_c_942_n 0.00197519f $X=6.375 $Y=0.685 $X2=0
+ $Y2=0
cc_424 N_A_303_311#_M1001_g N_VGND_c_942_n 0.00713723f $X=6.375 $Y=1.005 $X2=0
+ $Y2=0
cc_425 N_A_303_311#_c_510_n N_VGND_c_948_n 0.0384057f $X=6.125 $Y=0.38 $X2=0
+ $Y2=0
cc_426 N_A_303_311#_c_512_n N_VGND_c_948_n 6.41874e-19 $X=4.425 $Y=0.38 $X2=0
+ $Y2=0
cc_427 N_A_303_311#_c_516_n N_VGND_c_948_n 0.00650831f $X=4.495 $Y=1.005 $X2=0
+ $Y2=0
cc_428 N_A_303_311#_c_517_n N_VGND_c_948_n 0.0159246f $X=6.125 $Y=1.28 $X2=0
+ $Y2=0
cc_429 N_A_303_311#_c_518_n N_VGND_c_948_n 0.0194878f $X=4.517 $Y=0.395 $X2=0
+ $Y2=0
cc_430 N_A_303_311#_c_522_n N_VGND_c_950_n 0.0188956f $X=6.745 $Y=0.52 $X2=0
+ $Y2=0
cc_431 N_A_303_311#_c_524_n N_VGND_c_950_n 0.00183241f $X=6.375 $Y=0.685 $X2=0
+ $Y2=0
cc_432 N_A_303_311#_c_507_n N_VGND_c_952_n 0.0246623f $X=4.095 $Y=0.245 $X2=0
+ $Y2=0
cc_433 N_A_303_311#_c_512_n N_VGND_c_952_n 0.00176449f $X=4.425 $Y=0.38 $X2=0
+ $Y2=0
cc_434 N_A_303_311#_c_518_n N_VGND_c_952_n 0.0193397f $X=4.517 $Y=0.395 $X2=0
+ $Y2=0
cc_435 N_A_303_311#_c_506_n N_VGND_c_955_n 0.00917846f $X=2.11 $Y=1.555 $X2=0
+ $Y2=0
cc_436 N_A_303_311#_c_507_n N_VGND_c_955_n 0.0118444f $X=4.095 $Y=0.245 $X2=0
+ $Y2=0
cc_437 N_A_303_311#_c_508_n N_VGND_c_955_n 0.00156424f $X=2.185 $Y=0.245 $X2=0
+ $Y2=0
cc_438 N_A_303_311#_c_510_n N_VGND_c_955_n 0.00168196f $X=6.125 $Y=0.38 $X2=0
+ $Y2=0
cc_439 N_A_303_311#_c_512_n N_VGND_c_955_n 0.00702695f $X=4.425 $Y=0.38 $X2=0
+ $Y2=0
cc_440 N_A_303_311#_c_515_n N_VGND_c_955_n 0.00569458f $X=1.835 $Y=1.005 $X2=0
+ $Y2=0
cc_441 N_A_303_311#_c_516_n N_VGND_c_955_n 0.0221788f $X=4.495 $Y=1.005 $X2=0
+ $Y2=0
cc_442 N_A_303_311#_c_517_n N_VGND_c_955_n 0.0333443f $X=6.125 $Y=1.28 $X2=0
+ $Y2=0
cc_443 N_A_303_311#_c_518_n N_VGND_c_955_n 0.0276326f $X=4.517 $Y=0.395 $X2=0
+ $Y2=0
cc_444 N_A_303_311#_c_592_n N_VGND_c_955_n 0.00177927f $X=6.307 $Y=1.195 $X2=0
+ $Y2=0
cc_445 N_A_303_311#_c_522_n N_VGND_c_955_n 0.0401594f $X=6.745 $Y=0.52 $X2=0
+ $Y2=0
cc_446 N_A_303_311#_c_524_n N_VGND_c_955_n 0.0152583f $X=6.375 $Y=0.685 $X2=0
+ $Y2=0
cc_447 N_A_303_311#_c_517_n A_1027_159# 0.0017792f $X=6.125 $Y=1.28 $X2=0 $Y2=0
cc_448 N_CLK_c_662_n N_A_1438_171#_M1016_g 0.00119991f $X=8.417 $Y=3.125 $X2=0
+ $Y2=0
cc_449 N_CLK_c_698_n N_A_1438_171#_M1016_g 0.00186218f $X=8.515 $Y=1.89 $X2=0
+ $Y2=0
cc_450 N_CLK_M1011_g N_A_1438_171#_M1016_g 0.037824f $X=8.485 $Y=1.065 $X2=0
+ $Y2=0
cc_451 N_CLK_M1011_g N_A_1438_171#_c_749_n 0.00320621f $X=8.485 $Y=1.065 $X2=0
+ $Y2=0
cc_452 N_CLK_c_654_n N_A_1438_171#_c_750_n 0.00486018f $X=8.235 $Y=3.38 $X2=0
+ $Y2=0
cc_453 N_CLK_c_698_n N_A_1438_171#_c_750_n 0.0638256f $X=8.515 $Y=1.89 $X2=0
+ $Y2=0
cc_454 N_CLK_M1011_g N_A_1438_171#_c_750_n 0.0088703f $X=8.485 $Y=1.065 $X2=0
+ $Y2=0
cc_455 N_CLK_M1011_g N_A_1438_171#_c_752_n 0.00124571f $X=8.485 $Y=1.065 $X2=0
+ $Y2=0
cc_456 N_CLK_M1011_g N_A_1438_171#_c_753_n 0.0215344f $X=8.485 $Y=1.065 $X2=0
+ $Y2=0
cc_457 N_CLK_c_698_n N_A_1438_171#_c_754_n 0.0245959f $X=8.515 $Y=1.89 $X2=0
+ $Y2=0
cc_458 N_CLK_M1011_g N_A_1438_171#_c_754_n 0.0449828f $X=8.485 $Y=1.065 $X2=0
+ $Y2=0
cc_459 N_CLK_M1011_g N_A_1438_171#_c_755_n 0.0153138f $X=8.485 $Y=1.065 $X2=0
+ $Y2=0
cc_460 N_CLK_c_647_n N_VPWR_c_807_n 0.013978f $X=3.555 $Y=2.21 $X2=0 $Y2=0
cc_461 N_CLK_c_654_n N_VPWR_c_808_n 0.0129079f $X=8.235 $Y=3.38 $X2=4.08
+ $Y2=0.058
cc_462 N_CLK_c_658_n N_VPWR_c_808_n 0.00514727f $X=5.46 $Y=3.38 $X2=4.08
+ $Y2=0.058
cc_463 N_CLK_c_654_n N_VPWR_c_811_n 0.0211777f $X=8.235 $Y=3.38 $X2=9.84 $Y2=0
cc_464 N_CLK_c_654_n N_VPWR_c_812_n 0.0412835f $X=8.235 $Y=3.38 $X2=0 $Y2=0
cc_465 N_CLK_c_654_n N_VPWR_c_815_n 0.0251071f $X=8.235 $Y=3.38 $X2=0 $Y2=0
cc_466 N_CLK_c_661_n N_VPWR_c_816_n 0.00132264f $X=8.4 $Y=3.29 $X2=0 $Y2=0
cc_467 N_CLK_c_662_n N_VPWR_c_816_n 0.0677376f $X=8.417 $Y=3.125 $X2=0 $Y2=0
cc_468 N_CLK_M1011_g N_VPWR_c_816_n 0.00664218f $X=8.485 $Y=1.065 $X2=0 $Y2=0
cc_469 N_CLK_c_654_n N_VPWR_c_820_n 0.00723698f $X=8.235 $Y=3.38 $X2=0 $Y2=0
cc_470 N_CLK_c_654_n N_VPWR_c_823_n 0.0164637f $X=8.235 $Y=3.38 $X2=0 $Y2=0
cc_471 N_CLK_c_654_n N_VPWR_c_826_n 0.00685941f $X=8.235 $Y=3.38 $X2=0 $Y2=0
cc_472 N_CLK_c_654_n N_VPWR_c_833_n 0.00888031f $X=8.235 $Y=3.38 $X2=0 $Y2=0
cc_473 N_CLK_c_659_n N_VPWR_c_833_n 0.00303441f $X=8.485 $Y=3.095 $X2=0 $Y2=0
cc_474 N_CLK_c_660_n N_VPWR_c_833_n 0.0250527f $X=8.4 $Y=3.29 $X2=0 $Y2=0
cc_475 N_CLK_c_647_n N_VPWR_c_835_n 0.00567592f $X=3.555 $Y=2.21 $X2=0 $Y2=0
cc_476 N_CLK_c_650_n N_VPWR_c_835_n 0.0116752f $X=5.385 $Y=3.58 $X2=0 $Y2=0
cc_477 N_CLK_c_651_n N_VPWR_c_835_n 0.0032954f $X=4.295 $Y=3.58 $X2=0 $Y2=0
cc_478 N_CLK_c_654_n N_VPWR_c_835_n 0.0568213f $X=8.235 $Y=3.38 $X2=0 $Y2=0
cc_479 N_CLK_c_658_n N_VPWR_c_835_n 0.00530322f $X=5.46 $Y=3.38 $X2=0 $Y2=0
cc_480 N_CLK_c_659_n N_VPWR_c_835_n 0.00385655f $X=8.485 $Y=3.095 $X2=0 $Y2=0
cc_481 N_CLK_c_660_n N_VPWR_c_835_n 0.0133491f $X=8.4 $Y=3.29 $X2=0 $Y2=0
cc_482 N_CLK_M1011_g N_VGND_c_943_n 0.0063675f $X=8.485 $Y=1.065 $X2=4.08 $Y2=0
cc_483 N_CLK_M1011_g N_VGND_c_950_n 0.0215371f $X=8.485 $Y=1.065 $X2=0 $Y2=0
cc_484 N_CLK_M1005_g N_VGND_c_952_n 0.0301236f $X=3.555 $Y=0.87 $X2=0 $Y2=0
cc_485 N_CLK_M1005_g N_VGND_c_955_n 0.0079947f $X=3.555 $Y=0.87 $X2=0 $Y2=0
cc_486 N_CLK_M1011_g N_VGND_c_955_n 0.016429f $X=8.485 $Y=1.065 $X2=0 $Y2=0
cc_487 N_A_1438_171#_c_750_n N_VPWR_c_815_n 0.0250813f $X=8.095 $Y=2.36 $X2=0
+ $Y2=0
cc_488 N_A_1438_171#_M1016_g N_VPWR_c_816_n 0.033971f $X=9.325 $Y=2.965 $X2=0
+ $Y2=0
cc_489 N_A_1438_171#_c_752_n N_VPWR_c_816_n 0.00597948f $X=9.45 $Y=1.56 $X2=0
+ $Y2=0
cc_490 N_A_1438_171#_c_753_n N_VPWR_c_816_n 0.00249173f $X=9.45 $Y=1.56 $X2=0
+ $Y2=0
cc_491 N_A_1438_171#_c_754_n N_VPWR_c_816_n 0.00580055f $X=8.945 $Y=1.555 $X2=0
+ $Y2=0
cc_492 N_A_1438_171#_c_750_n N_VPWR_c_826_n 0.00153188f $X=8.095 $Y=2.36 $X2=0
+ $Y2=0
cc_493 N_A_1438_171#_c_750_n N_VPWR_c_833_n 9.74195e-19 $X=8.095 $Y=2.36 $X2=0
+ $Y2=0
cc_494 N_A_1438_171#_M1016_g N_VPWR_c_834_n 0.0277286f $X=9.325 $Y=2.965 $X2=0
+ $Y2=0
cc_495 N_A_1438_171#_M1016_g N_VPWR_c_835_n 0.0239408f $X=9.325 $Y=2.965 $X2=0
+ $Y2=0
cc_496 N_A_1438_171#_c_750_n N_VPWR_c_835_n 0.005784f $X=8.095 $Y=2.36 $X2=0
+ $Y2=0
cc_497 N_A_1438_171#_c_755_n N_GCLK_c_918_n 5.566e-19 $X=9.28 $Y=1.395 $X2=0
+ $Y2=0
cc_498 N_A_1438_171#_M1016_g GCLK 0.0195593f $X=9.325 $Y=2.965 $X2=0 $Y2=0
cc_499 N_A_1438_171#_M1016_g GCLK 0.00717157f $X=9.325 $Y=2.965 $X2=0 $Y2=0
cc_500 N_A_1438_171#_c_752_n GCLK 0.0277798f $X=9.45 $Y=1.56 $X2=0 $Y2=0
cc_501 N_A_1438_171#_c_753_n GCLK 0.00929555f $X=9.45 $Y=1.56 $X2=0 $Y2=0
cc_502 N_A_1438_171#_c_755_n GCLK 0.00675953f $X=9.28 $Y=1.395 $X2=0 $Y2=0
cc_503 N_A_1438_171#_c_753_n N_VGND_c_943_n 8.22277e-19 $X=9.45 $Y=1.56 $X2=4.08
+ $Y2=0
cc_504 N_A_1438_171#_c_754_n N_VGND_c_943_n 0.0237894f $X=8.945 $Y=1.555
+ $X2=4.08 $Y2=0
cc_505 N_A_1438_171#_c_755_n N_VGND_c_943_n 0.0154225f $X=9.28 $Y=1.395 $X2=4.08
+ $Y2=0
cc_506 N_A_1438_171#_c_748_n N_VGND_c_950_n 0.0430498f $X=7.955 $Y=1.05 $X2=0
+ $Y2=0
cc_507 N_A_1438_171#_c_755_n N_VGND_c_954_n 0.0290307f $X=9.28 $Y=1.395 $X2=0
+ $Y2=0
cc_508 N_A_1438_171#_c_748_n N_VGND_c_955_n 0.0294463f $X=7.955 $Y=1.05 $X2=0
+ $Y2=0
cc_509 N_A_1438_171#_c_755_n N_VGND_c_955_n 0.0243873f $X=9.28 $Y=1.395 $X2=0
+ $Y2=0
cc_510 N_A_1438_171#_c_748_n A_1591_171# 0.00283135f $X=7.955 $Y=1.05 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_835_n N_GCLK_M1016_d 0.00221032f $X=9.36 $Y=3.56 $X2=0 $Y2=0
cc_512 N_VPWR_c_816_n GCLK 0.0188494f $X=8.935 $Y=2.36 $X2=9.84 $Y2=4.07
cc_513 N_VPWR_c_834_n GCLK 0.0151461f $X=9.36 $Y=3.56 $X2=9.84 $Y2=4.07
cc_514 N_VPWR_c_835_n GCLK 0.0448072f $X=9.36 $Y=3.56 $X2=9.84 $Y2=4.07
cc_515 N_GCLK_c_918_n N_VGND_c_954_n 0.00592735f $X=9.715 $Y=0.68 $X2=0 $Y2=0
cc_516 N_GCLK_M1010_d N_VGND_c_955_n 0.00221032f $X=9.575 $Y=0.535 $X2=0 $Y2=0
cc_517 N_GCLK_c_918_n N_VGND_c_955_n 0.0349083f $X=9.715 $Y=0.68 $X2=0 $Y2=0
