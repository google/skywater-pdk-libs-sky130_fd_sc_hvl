* File: sky130_fd_sc_hvl__dfxtp_1.pex.spice
* Created: Fri Aug 28 09:34:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%VNB 5 7 11 25
c87 11 0 8.99003e-20 $X=0.24 $Y=0
c88 5 0 1.07121e-19 $X=-0.33 $Y=-0.265
r89 7 25 1.04167e-05 $w=1.2e-05 $l=1e-09 $layer=MET1_cond $X=6 $Y=0.057 $X2=6
+ $Y2=0.058
r90 7 11 0.00059375 $w=1.2e-05 $l=5.7e-08 $layer=MET1_cond $X=6 $Y=0.057 $X2=6
+ $Y2=0
r91 5 11 0.744 $w=1.7e-07 $l=2.125e-06 $layer=mcon $count=12 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r92 5 11 0.744 $w=1.7e-07 $l=2.125e-06 $layer=mcon $count=12 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%VPB 4 6 14 21
r108 10 21 0.00059375 $w=1.2e-05 $l=5.7e-08 $layer=MET1_cond $X=6 $Y=4.07 $X2=6
+ $Y2=4.013
r109 10 14 0.744 $w=1.7e-07 $l=2.125e-06 $layer=mcon $count=12 $X=11.76 $Y=4.07
+ $X2=11.76 $Y2=4.07
r110 9 14 751.572 $w=1.68e-07 $l=1.152e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=11.76 $Y2=4.07
r111 9 10 0.744 $w=1.7e-07 $l=2.125e-06 $layer=mcon $count=12 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r112 6 21 1.04167e-05 $w=1.2e-05 $l=1e-09 $layer=MET1_cond $X=6 $Y=4.012 $X2=6
+ $Y2=4.013
r113 4 14 14.56 $w=1.7e-07 $l=1.18024e-05 $layer=licon1_NTAP_notbjt $count=12
+ $X=0 $Y=3.985 $X2=11.76 $Y2=4.07
r114 4 9 14.56 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=12
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%CLK 3 7 8 9 11 12 13 17
c30 17 0 6.26942e-20 $X=0.705 $Y=2.07
r31 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=2.035
+ $X2=0.705 $Y2=2.405
r32 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.705
+ $Y=2.07 $X2=0.705 $Y2=2.07
r33 10 17 34.4682 $w=5.2e-07 $l=3.35e-07 $layer=POLY_cond $X=0.675 $Y=2.405
+ $X2=0.675 $Y2=2.07
r34 10 11 26.7515 $w=5.2e-07 $l=2.6e-07 $layer=POLY_cond $X=0.675 $Y=2.405
+ $X2=0.675 $Y2=2.665
r35 8 17 66.3642 $w=5.2e-07 $l=6.45e-07 $layer=POLY_cond $X=0.675 $Y=1.425
+ $X2=0.675 $Y2=2.07
r36 8 9 26.7515 $w=5.2e-07 $l=2.6e-07 $layer=POLY_cond $X=0.675 $Y=1.425
+ $X2=0.675 $Y2=1.165
r37 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.685 $Y=0.845 $X2=0.685
+ $Y2=1.165
r38 3 11 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.665 $Y=3.17 $X2=0.665
+ $Y2=2.665
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%A_30_127# 1 2 7 9 13 17 19 21 23 25 26 28
+ 30 32 37 41 43 45 46 47 49 53 58 61 62 63 66 70 75
c190 75 0 4.66275e-20 $X=6.87 $Y=2.39
c191 70 0 1.07121e-19 $X=2.735 $Y=1.845
c192 28 0 2.07934e-19 $X=8.185 $Y=1.115
c193 23 0 1.01852e-20 $X=7.025 $Y=2.605
c194 19 0 1.60989e-19 $X=4.66 $Y=2.585
r195 76 85 40.2282 $w=6.53e-07 $l=5.45e-07 $layer=POLY_cond $X=7.102 $Y=2.39
+ $X2=7.102 $Y2=1.845
r196 75 78 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=6.83 $Y=2.39 $X2=6.83
+ $Y2=2.47
r197 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.87
+ $Y=2.39 $X2=6.87 $Y2=2.39
r198 69 80 8.45614 $w=5.7e-07 $l=1e-07 $layer=POLY_cond $X=1.43 $Y=2.06 $X2=1.43
+ $Y2=1.96
r199 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.33
+ $Y=2.06 $X2=1.33 $Y2=2.06
r200 66 80 22.5276 $w=5.7e-07 $l=2.4e-07 $layer=POLY_cond $X=1.43 $Y=1.72
+ $X2=1.43 $Y2=1.96
r201 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.33
+ $Y=1.72 $X2=1.33 $Y2=1.72
r202 61 78 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.705 $Y=2.47
+ $X2=6.83 $Y2=2.47
r203 61 62 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=6.705 $Y=2.47
+ $X2=4.89 $Y2=2.47
r204 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.725
+ $Y=2.05 $X2=4.725 $Y2=2.05
r205 56 62 7.72402 $w=1.7e-07 $l=2.01057e-07 $layer=LI1_cond $X=4.727 $Y=2.385
+ $X2=4.89 $Y2=2.47
r206 56 58 11.879 $w=3.23e-07 $l=3.35e-07 $layer=LI1_cond $X=4.727 $Y=2.385
+ $X2=4.727 $Y2=2.05
r207 54 59 37.3303 $w=8.78e-07 $l=6.8e-07 $layer=POLY_cond $X=4.16 $Y=1.37
+ $X2=4.16 $Y2=2.05
r208 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.595
+ $Y=1.37 $X2=3.595 $Y2=1.37
r209 51 53 17.6256 $w=2.53e-07 $l=3.9e-07 $layer=LI1_cond $X=3.557 $Y=1.76
+ $X2=3.557 $Y2=1.37
r210 50 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.82 $Y=1.845
+ $X2=2.735 $Y2=1.845
r211 49 51 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=3.43 $Y=1.845
+ $X2=3.557 $Y2=1.76
r212 49 50 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.43 $Y=1.845
+ $X2=2.82 $Y2=1.845
r213 48 68 3.16044 $w=2.95e-07 $l=1.25e-07 $layer=LI1_cond $X=1.415 $Y=2.077
+ $X2=1.29 $Y2=2.077
r214 47 70 15.1358 $w=1.68e-07 $l=2.32e-07 $layer=LI1_cond $X=2.735 $Y=2.077
+ $X2=2.735 $Y2=1.845
r215 47 48 48.2463 $w=2.93e-07 $l=1.235e-06 $layer=LI1_cond $X=2.65 $Y=2.077
+ $X2=1.415 $Y2=2.077
r216 46 68 3.71667 $w=2.5e-07 $l=1.47e-07 $layer=LI1_cond $X=1.29 $Y=1.93
+ $X2=1.29 $Y2=2.077
r217 45 65 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.29 $Y=1.725
+ $X2=1.29 $Y2=1.64
r218 45 46 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=1.29 $Y=1.725
+ $X2=1.29 $Y2=1.93
r219 44 63 2.90867 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.38 $Y=1.64
+ $X2=0.245 $Y2=1.64
r220 43 65 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.165 $Y=1.64
+ $X2=1.29 $Y2=1.64
r221 43 44 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.165 $Y=1.64
+ $X2=0.38 $Y2=1.64
r222 39 63 3.58051 $w=2.6e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.235 $Y=1.725
+ $X2=0.245 $Y2=1.64
r223 39 41 56.0087 $w=2.48e-07 $l=1.215e-06 $layer=LI1_cond $X=0.235 $Y=1.725
+ $X2=0.235 $Y2=2.94
r224 35 63 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=1.555
+ $X2=0.245 $Y2=1.64
r225 35 37 30.305 $w=2.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.245 $Y=1.555
+ $X2=0.245 $Y2=0.845
r226 32 66 23.4662 $w=5.7e-07 $l=2.5e-07 $layer=POLY_cond $X=1.43 $Y=1.47
+ $X2=1.43 $Y2=1.72
r227 32 33 27.696 $w=5.7e-07 $l=2.85e-07 $layer=POLY_cond $X=1.43 $Y=1.47
+ $X2=1.43 $Y2=1.185
r228 28 34 67.9266 $w=5.18e-07 $l=7.37462e-07 $layer=POLY_cond $X=8.185 $Y=1.115
+ $X2=8.17 $Y2=1.845
r229 28 30 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=8.185 $Y=1.115
+ $X2=8.185 $Y2=0.775
r230 27 85 18.0178 $w=3.4e-07 $l=3.98e-07 $layer=POLY_cond $X=7.5 $Y=1.845
+ $X2=7.102 $Y2=1.845
r231 26 34 12.6477 $w=3.4e-07 $l=2.65e-07 $layer=POLY_cond $X=7.905 $Y=1.845
+ $X2=8.17 $Y2=1.845
r232 26 27 68.7359 $w=3.4e-07 $l=4.05e-07 $layer=POLY_cond $X=7.905 $Y=1.845
+ $X2=7.5 $Y2=1.845
r233 23 76 18.6366 $w=6.53e-07 $l=2.50559e-07 $layer=POLY_cond $X=7.025 $Y=2.605
+ $X2=7.102 $Y2=2.39
r234 23 25 58.804 $w=5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.025 $Y=2.605
+ $X2=7.025 $Y2=3.215
r235 19 59 38.2298 $w=8.78e-07 $l=7.44127e-07 $layer=POLY_cond $X=4.66 $Y=2.585
+ $X2=4.16 $Y2=2.05
r236 19 21 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.66 $Y=2.585 $X2=4.66
+ $Y2=2.925
r237 15 54 22.8585 $w=8.78e-07 $l=4.18509e-07 $layer=POLY_cond $X=3.85 $Y=1.115
+ $X2=4.16 $Y2=1.37
r238 15 17 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.85 $Y=1.115 $X2=3.85
+ $Y2=0.775
r239 13 33 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.465 $Y=0.845
+ $X2=1.465 $Y2=1.185
r240 7 69 52.8894 $w=5.58e-07 $l=6.12454e-07 $layer=POLY_cond $X=1.445 $Y=2.665
+ $X2=1.43 $Y2=2.06
r241 7 9 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.445 $Y=2.665
+ $X2=1.445 $Y2=3.17
r242 2 41 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.795 $X2=0.275 $Y2=2.94
r243 1 37 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.635 $X2=0.295 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%D 2 5 9 13 15 16 21 24
c56 24 0 9.13616e-20 $X=2.95 $Y=1.59
c57 21 0 6.26942e-20 $X=2.305 $Y=1.655
r58 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.305
+ $Y=1.655 $X2=2.305 $Y2=1.655
r59 16 21 8.24709 $w=1.93e-07 $l=1.45e-07 $layer=LI1_cond $X=2.16 $Y=1.652
+ $X2=2.305 $Y2=1.652
r60 15 16 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.652
+ $X2=2.16 $Y2=1.652
r61 7 24 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.95 $Y=1.34 $X2=2.95
+ $Y2=1.59
r62 7 9 60.4583 $w=5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.95 $Y=1.34 $X2=2.95
+ $Y2=0.775
r63 3 13 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.775 $Y=2.685
+ $X2=2.775 $Y2=2.435
r64 3 5 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.775 $Y=2.685 $X2=2.775
+ $Y2=3.025
r65 2 13 39.0572 $w=5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.41 $Y=2.435
+ $X2=2.775 $Y2=2.435
r66 1 24 57.7832 $w=5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.41 $Y=1.59 $X2=2.95
+ $Y2=1.59
r67 1 20 11.2356 $w=5e-07 $l=1.05e-07 $layer=POLY_cond $X=2.41 $Y=1.59 $X2=2.305
+ $Y2=1.59
r68 1 2 31.825 $w=5.8e-07 $l=3.45e-07 $layer=POLY_cond $X=2.41 $Y=1.84 $X2=2.41
+ $Y2=2.185
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%A_339_559# 1 2 7 9 12 16 18 19 20 21 23 24
+ 25 27 28 29 32 33 35 38 39 42 43 44 46 48 50 53 56 66 68 72 75 80
c217 75 0 2.3324e-19 $X=4.825 $Y=0.775
c218 66 0 1.40845e-19 $X=7.57 $Y=1.285
c219 53 0 8.73223e-20 $X=8.085 $Y=2.39
c220 46 0 4.89168e-20 $X=7.365 $Y=1.125
c221 38 0 1.60989e-19 $X=4.89 $Y=1.175
c222 18 0 6.43548e-20 $X=2.65 $Y=2.53
c223 7 0 1.84265e-19 $X=8.405 $Y=2.605
r224 65 80 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.405 $Y=1.28
+ $X2=7.405 $Y2=0.775
r225 64 66 4.50173 $w=3.18e-07 $l=1.25e-07 $layer=LI1_cond $X=7.445 $Y=1.285
+ $X2=7.57 $Y2=1.285
r226 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.445
+ $Y=1.28 $X2=7.445 $Y2=1.28
r227 61 64 2.88111 $w=3.18e-07 $l=8e-08 $layer=LI1_cond $X=7.365 $Y=1.285
+ $X2=7.445 $Y2=1.285
r228 60 75 51.8979 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.825 $Y=1.26
+ $X2=4.825 $Y2=0.775
r229 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.89
+ $Y=1.26 $X2=4.89 $Y2=1.26
r230 56 57 8.296 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=3.675 $Y=3.22
+ $X2=3.675 $Y2=3.39
r231 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.085
+ $Y=2.39 $X2=8.085 $Y2=2.39
r232 51 68 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.655 $Y=2.37
+ $X2=7.57 $Y2=2.37
r233 51 53 17.0879 $w=2.88e-07 $l=4.3e-07 $layer=LI1_cond $X=7.655 $Y=2.37
+ $X2=8.085 $Y2=2.37
r234 49 68 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.57 $Y=2.515
+ $X2=7.57 $Y2=2.37
r235 49 50 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.57 $Y=2.515
+ $X2=7.57 $Y2=3.135
r236 48 68 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.57 $Y=2.225
+ $X2=7.57 $Y2=2.37
r237 47 66 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=7.57 $Y=1.445
+ $X2=7.57 $Y2=1.285
r238 47 48 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=7.57 $Y=1.445
+ $X2=7.57 $Y2=2.225
r239 46 61 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=7.365 $Y=1.125
+ $X2=7.365 $Y2=1.285
r240 45 46 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.365 $Y=0.435
+ $X2=7.365 $Y2=1.125
r241 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.28 $Y=0.35
+ $X2=7.365 $Y2=0.435
r242 43 44 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.28 $Y=0.35
+ $X2=6.555 $Y2=0.35
r243 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.47 $Y=0.435
+ $X2=6.555 $Y2=0.35
r244 41 42 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.47 $Y=0.435
+ $X2=6.47 $Y2=1.175
r245 40 59 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.055 $Y=1.26
+ $X2=4.89 $Y2=1.26
r246 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.385 $Y=1.26
+ $X2=6.47 $Y2=1.175
r247 39 40 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=6.385 $Y=1.26
+ $X2=5.055 $Y2=1.26
r248 38 59 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.89 $Y=1.175
+ $X2=4.89 $Y2=1.26
r249 37 38 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=4.89 $Y=0.435
+ $X2=4.89 $Y2=1.175
r250 36 56 2.99516 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.84 $Y=3.22
+ $X2=3.675 $Y2=3.22
r251 35 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.485 $Y=3.22
+ $X2=7.57 $Y2=3.135
r252 35 36 237.802 $w=1.68e-07 $l=3.645e-06 $layer=LI1_cond $X=7.485 $Y=3.22
+ $X2=3.84 $Y2=3.22
r253 33 72 57.2482 $w=5e-07 $l=5.35e-07 $layer=POLY_cond $X=3.65 $Y=2.545
+ $X2=3.65 $Y2=3.08
r254 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.675
+ $Y=2.545 $X2=3.675 $Y2=2.545
r255 30 56 3.8884 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=3.135
+ $X2=3.675 $Y2=3.22
r256 30 32 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=3.675 $Y=3.135
+ $X2=3.675 $Y2=2.545
r257 28 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.725 $Y=0.35
+ $X2=4.89 $Y2=0.435
r258 28 29 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=4.725 $Y=0.35
+ $X2=3.115 $Y2=0.35
r259 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.03 $Y=0.435
+ $X2=3.115 $Y2=0.35
r260 26 27 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.03 $Y=0.435
+ $X2=3.03 $Y2=1.205
r261 24 57 2.99516 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.51 $Y=3.39
+ $X2=3.675 $Y2=3.39
r262 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.51 $Y=3.39
+ $X2=2.82 $Y2=3.39
r263 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.735 $Y=3.305
+ $X2=2.82 $Y2=3.39
r264 22 23 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.735 $Y=2.615
+ $X2=2.735 $Y2=3.305
r265 20 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.945 $Y=1.29
+ $X2=3.03 $Y2=1.205
r266 20 21 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=2.945 $Y=1.29
+ $X2=2.02 $Y2=1.29
r267 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.65 $Y=2.53
+ $X2=2.735 $Y2=2.615
r268 18 19 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.65 $Y=2.53 $X2=2
+ $Y2=2.53
r269 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.855 $Y=1.205
+ $X2=2.02 $Y2=1.29
r270 14 16 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.855 $Y=1.205
+ $X2=1.855 $Y2=0.845
r271 10 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.835 $Y=2.615
+ $X2=2 $Y2=2.53
r272 10 12 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.835 $Y=2.615
+ $X2=1.835 $Y2=2.94
r273 7 54 46.834 $w=3.8e-07 $l=3.2e-07 $layer=POLY_cond $X=8.405 $Y=2.415
+ $X2=8.085 $Y2=2.415
r274 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.405 $Y=2.605 $X2=8.405
+ $Y2=2.925
r275 2 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=2.795 $X2=1.835 $Y2=2.94
r276 1 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.715
+ $Y=0.635 $X2=1.855 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%A_1024_371# 1 2 9 13 15 17 23 28 29 33 36
c69 29 0 9.70108e-20 $X=5.6 $Y=1.96
c70 28 0 1.84265e-19 $X=7.22 $Y=2.755
r71 33 40 47.264 $w=6.65e-07 $l=5.45e-07 $layer=POLY_cond $X=5.452 $Y=2.04
+ $X2=5.452 $Y2=2.585
r72 33 39 18.3 $w=6.65e-07 $l=1.85e-07 $layer=POLY_cond $X=5.452 $Y=2.04
+ $X2=5.452 $Y2=1.855
r73 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.6
+ $Y=2.04 $X2=5.6 $Y2=2.04
r74 29 32 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.6 $Y=1.96 $X2=5.6
+ $Y2=2.04
r75 27 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.22 $Y=2.045
+ $X2=7.22 $Y2=1.96
r76 27 28 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=7.22 $Y=2.045
+ $X2=7.22 $Y2=2.755
r77 23 26 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=6.9 $Y=0.7 $X2=6.9
+ $Y2=1.19
r78 21 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.9 $Y=1.96 $X2=7.22
+ $Y2=1.96
r79 21 26 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=6.9 $Y=1.875
+ $X2=6.9 $Y2=1.19
r80 17 28 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=7.135 $Y=2.855
+ $X2=7.22 $Y2=2.755
r81 17 19 27.7273 $w=1.98e-07 $l=5e-07 $layer=LI1_cond $X=7.135 $Y=2.855
+ $X2=6.635 $Y2=2.855
r82 16 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.765 $Y=1.96
+ $X2=5.6 $Y2=1.96
r83 15 21 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.735 $Y=1.96
+ $X2=6.9 $Y2=1.96
r84 15 16 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=6.735 $Y=1.96
+ $X2=5.765 $Y2=1.96
r85 13 39 115.566 $w=5e-07 $l=1.08e-06 $layer=POLY_cond $X=5.535 $Y=0.775
+ $X2=5.535 $Y2=1.855
r86 9 40 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.37 $Y=2.925 $X2=5.37
+ $Y2=2.585
r87 2 19 600 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_PDIFF $count=1 $X=6.495
+ $Y=2.715 $X2=6.635 $Y2=2.855
r88 1 26 182 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_NDIFF $count=1 $X=6.76
+ $Y=0.565 $X2=6.9 $Y2=1.19
r89 1 23 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=6.76
+ $Y=0.565 $X2=6.9 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%A_780_574# 1 2 9 11 13 16 22 26 27 29
c72 22 0 1.01852e-20 $X=6.18 $Y=1.61
c73 11 0 2.84484e-19 $X=6.51 $Y=1.425
r74 26 27 8.98601 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=4.22 $Y=2.855
+ $X2=4.22 $Y2=2.675
r75 23 32 7.1705 $w=4.85e-07 $l=6.5e-08 $layer=POLY_cond $X=6.18 $Y=1.667
+ $X2=6.245 $Y2=1.667
r76 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.18
+ $Y=1.61 $X2=6.18 $Y2=1.61
r77 20 29 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.545 $Y=1.61
+ $X2=4.38 $Y2=1.61
r78 20 22 106.668 $w=1.68e-07 $l=1.635e-06 $layer=LI1_cond $X=4.545 $Y=1.61
+ $X2=6.18 $Y2=1.61
r79 18 29 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.3 $Y=1.695
+ $X2=4.38 $Y2=1.61
r80 18 27 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=4.3 $Y=1.695 $X2=4.3
+ $Y2=2.675
r81 14 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=1.525
+ $X2=4.38 $Y2=1.61
r82 14 16 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=4.38 $Y=1.525
+ $X2=4.38 $Y2=0.78
r83 11 32 29.2336 $w=4.85e-07 $l=2.65e-07 $layer=POLY_cond $X=6.51 $Y=1.667
+ $X2=6.245 $Y2=1.667
r84 11 13 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.51 $Y=1.425 $X2=6.51
+ $Y2=0.94
r85 7 32 2.09349 $w=5e-07 $l=2.43e-07 $layer=POLY_cond $X=6.245 $Y=1.91
+ $X2=6.245 $Y2=1.667
r86 7 9 139.643 $w=5e-07 $l=1.305e-06 $layer=POLY_cond $X=6.245 $Y=1.91
+ $X2=6.245 $Y2=3.215
r87 2 26 600 $w=1.7e-07 $l=3.27414e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=2.87 $X2=4.22 $Y2=2.855
r88 1 16 182 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_NDIFF $count=1 $X=4.1
+ $Y=0.565 $X2=4.38 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%A_1729_87# 1 2 9 13 17 21 23 25 28 32 34 36
+ 45 46 50 53
c79 53 0 1.92716e-19 $X=11.085 $Y=1.835
c80 25 0 5.1014e-20 $X=9.165 $Y=1.85
c81 23 0 1.08003e-19 $X=9.165 $Y=1.595
c82 13 0 2.63685e-19 $X=9.115 $Y=2.925
r83 51 52 12.3877 $w=3.25e-07 $l=3.3e-07 $layer=LI1_cond $X=10.362 $Y=1.51
+ $X2=10.362 $Y2=1.84
r84 50 57 18.0627 $w=7.2e-07 $l=1.85e-07 $layer=POLY_cond $X=9.005 $Y=1.51
+ $X2=9.005 $Y2=1.325
r85 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.165
+ $Y=1.51 $X2=9.165 $Y2=1.51
r86 46 53 5.30422 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=11.335 $Y=1.835
+ $X2=11.085 $Y2=1.835
r87 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=11.295
+ $Y=1.84 $X2=11.295 $Y2=1.84
r88 43 53 50.2928 $w=5e-07 $l=4.7e-07 $layer=POLY_cond $X=10.615 $Y=1.835
+ $X2=11.085 $Y2=1.835
r89 42 45 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.615 $Y=1.84
+ $X2=11.295 $Y2=1.84
r90 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=10.615
+ $Y=1.84 $X2=10.615 $Y2=1.84
r91 40 52 0.623162 $w=3.3e-07 $l=1.83e-07 $layer=LI1_cond $X=10.545 $Y=1.84
+ $X2=10.362 $Y2=1.84
r92 40 42 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=10.545 $Y=1.84
+ $X2=10.615 $Y2=1.84
r93 36 38 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=10.38 $Y=2.86
+ $X2=10.38 $Y2=3.57
r94 34 52 6.1 $w=3.3e-07 $l=1.73767e-07 $layer=LI1_cond $X=10.38 $Y=2.005
+ $X2=10.362 $Y2=1.84
r95 34 36 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=10.38 $Y=2.005
+ $X2=10.38 $Y2=2.86
r96 30 51 3.14242 $w=3.3e-07 $l=9.31128e-08 $layer=LI1_cond $X=10.345 $Y=1.425
+ $X2=10.362 $Y2=1.51
r97 30 32 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=10.345 $Y=1.425
+ $X2=10.345 $Y2=0.69
r98 29 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.33 $Y=1.51
+ $X2=9.165 $Y2=1.51
r99 28 51 4.53325 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.18 $Y=1.51
+ $X2=10.362 $Y2=1.51
r100 28 29 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=10.18 $Y=1.51
+ $X2=9.33 $Y2=1.51
r101 26 59 16.6344 $w=7.2e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=1.85
+ $X2=9.005 $Y2=2.015
r102 26 50 24.2803 $w=7.2e-07 $l=3.4e-07 $layer=POLY_cond $X=9.005 $Y=1.85
+ $X2=9.005 $Y2=1.51
r103 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.165
+ $Y=1.85 $X2=9.165 $Y2=1.85
r104 23 49 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.165 $Y=1.595
+ $X2=9.165 $Y2=1.51
r105 23 25 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=9.165 $Y=1.595
+ $X2=9.165 $Y2=1.85
r106 19 46 20.4101 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=11.335 $Y=2.085
+ $X2=11.335 $Y2=1.835
r107 19 21 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=11.335 $Y=2.085
+ $X2=11.335 $Y2=2.965
r108 15 46 20.4101 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=11.335 $Y=1.585
+ $X2=11.335 $Y2=1.835
r109 15 17 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=11.335 $Y=1.585
+ $X2=11.335 $Y2=1.08
r110 13 59 97.3754 $w=5e-07 $l=9.1e-07 $layer=POLY_cond $X=9.115 $Y=2.925
+ $X2=9.115 $Y2=2.015
r111 9 57 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=8.895 $Y=0.775
+ $X2=8.895 $Y2=1.325
r112 2 38 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=10.24
+ $Y=2.715 $X2=10.38 $Y2=3.57
r113 2 36 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.24
+ $Y=2.715 $X2=10.38 $Y2=2.86
r114 1 32 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=10.205
+ $Y=0.565 $X2=10.345 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%A_1455_543# 1 2 9 11 13 15 17 19 21 24 26
+ 27 31 35 39
c93 31 0 1.92716e-19 $X=9.87 $Y=1.94
c94 21 0 1.76363e-19 $X=8.43 $Y=2.78
r95 35 36 5.88596 $w=3.42e-07 $l=1.65e-07 $layer=LI1_cond $X=7.817 $Y=0.775
+ $X2=7.817 $Y2=0.94
r96 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.87
+ $Y=1.94 $X2=9.87 $Y2=1.94
r97 29 31 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.87 $Y=2.275
+ $X2=9.87 $Y2=1.94
r98 28 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.6 $Y=2.36 $X2=8.515
+ $Y2=2.36
r99 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.705 $Y=2.36
+ $X2=9.87 $Y2=2.275
r100 27 28 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=9.705 $Y=2.36
+ $X2=8.6 $Y2=2.36
r101 25 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.515 $Y=2.445
+ $X2=8.515 $Y2=2.36
r102 25 26 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.515 $Y=2.445
+ $X2=8.515 $Y2=2.695
r103 24 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.515 $Y=2.275
+ $X2=8.515 $Y2=2.36
r104 23 24 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=8.515 $Y=1.025
+ $X2=8.515 $Y2=2.275
r105 22 38 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.085 $Y=2.78
+ $X2=7.96 $Y2=2.78
r106 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.43 $Y=2.78
+ $X2=8.515 $Y2=2.695
r107 21 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.43 $Y=2.78
+ $X2=8.085 $Y2=2.78
r108 20 36 4.83608 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=8.005 $Y=0.94
+ $X2=7.817 $Y2=0.94
r109 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.43 $Y=0.94
+ $X2=8.515 $Y2=1.025
r110 19 20 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=8.43 $Y=0.94
+ $X2=8.005 $Y2=0.94
r111 15 38 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=2.865
+ $X2=7.96 $Y2=2.78
r112 15 17 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=7.96 $Y=2.865
+ $X2=7.96 $Y2=3.215
r113 11 32 46.6392 $w=5.48e-07 $l=5.38818e-07 $layer=POLY_cond $X=9.99 $Y=2.465
+ $X2=9.962 $Y2=1.94
r114 11 13 80.2544 $w=5e-07 $l=7.5e-07 $layer=POLY_cond $X=9.99 $Y=2.465
+ $X2=9.99 $Y2=3.215
r115 7 32 44.0006 $w=5.48e-07 $l=4.98488e-07 $layer=POLY_cond $X=9.955 $Y=1.445
+ $X2=9.962 $Y2=1.94
r116 7 9 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=9.955 $Y=1.445
+ $X2=9.955 $Y2=0.94
r117 2 38 600 $w=1.7e-07 $l=7.13828e-07 $layer=licon1_PDIFF $count=1 $X=7.275
+ $Y=2.715 $X2=7.92 $Y2=2.86
r118 2 17 300 $w=1.7e-07 $l=8.59375e-07 $layer=licon1_PDIFF $count=2 $X=7.275
+ $Y=2.715 $X2=7.92 $Y2=3.215
r119 1 35 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.655
+ $Y=0.565 $X2=7.795 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%VPWR 1 2 3 4 5 16 19 28 39 44 55 61
r74 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.2 $Y=3.59
+ $X2=11.2 $Y2=3.59
r75 58 60 0.40545 $w=5.88e-07 $l=2e-08 $layer=LI1_cond $X=11.02 $Y=3.57
+ $X2=11.02 $Y2=3.59
r76 55 58 24.5297 $w=5.88e-07 $l=1.21e-06 $layer=LI1_cond $X=11.02 $Y=2.36
+ $X2=11.02 $Y2=3.57
r77 52 61 0.595053 $w=3.7e-07 $l=1.55e-06 $layer=MET1_cond $X=9.65 $Y=3.63
+ $X2=11.2 $Y2=3.63
r78 50 52 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.93 $Y=3.63
+ $X2=9.65 $Y2=3.63
r79 49 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.65 $Y=3.59
+ $X2=9.65 $Y2=3.59
r80 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.93 $Y=3.59
+ $X2=8.93 $Y2=3.59
r81 47 49 4.81579 $w=9.48e-07 $l=3.75e-07 $layer=LI1_cond $X=9.29 $Y=3.215
+ $X2=9.29 $Y2=3.59
r82 44 47 4.55895 $w=9.48e-07 $l=3.55e-07 $layer=LI1_cond $X=9.29 $Y=2.86
+ $X2=9.29 $Y2=3.215
r83 39 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.905 $Y=3.6
+ $X2=5.905 $Y2=3.6
r84 36 41 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=5.185 $Y=3.63
+ $X2=5.905 $Y2=3.63
r85 35 39 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=5.185 $Y=3.61
+ $X2=5.855 $Y2=3.61
r86 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.185 $Y=3.6
+ $X2=5.185 $Y2=3.6
r87 32 36 1.09413 $w=3.7e-07 $l=2.85e-06 $layer=MET1_cond $X=2.335 $Y=3.63
+ $X2=5.185 $Y2=3.63
r88 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.335 $Y=3.59
+ $X2=2.335 $Y2=3.59
r89 28 31 26.0452 $w=2.48e-07 $l=5.65e-07 $layer=LI1_cond $X=2.345 $Y=3.025
+ $X2=2.345 $Y2=3.59
r90 25 32 0.368549 $w=3.7e-07 $l=9.6e-07 $layer=MET1_cond $X=1.375 $Y=3.63
+ $X2=2.335 $Y2=3.63
r91 23 25 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.655 $Y=3.63
+ $X2=1.375 $Y2=3.63
r92 22 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.375 $Y=3.59
+ $X2=1.375 $Y2=3.59
r93 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.655 $Y=3.59
+ $X2=0.655 $Y2=3.59
r94 19 22 8.60421 $w=9.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=2.92
+ $X2=1.015 $Y2=3.59
r95 16 50 1.12484 $w=3.7e-07 $l=2.93e-06 $layer=MET1_cond $X=6 $Y=3.63 $X2=8.93
+ $Y2=3.63
r96 16 41 0.036471 $w=3.7e-07 $l=9.5e-08 $layer=MET1_cond $X=6 $Y=3.63 $X2=5.905
+ $Y2=3.63
r97 5 58 300 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_PDIFF $count=2 $X=10.82
+ $Y=2.215 $X2=10.945 $Y2=3.57
r98 5 55 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=10.82
+ $Y=2.215 $X2=10.945 $Y2=2.36
r99 4 47 300 $w=1.7e-07 $l=6.06218e-07 $layer=licon1_PDIFF $count=2 $X=9.365
+ $Y=2.715 $X2=9.6 $Y2=3.215
r100 4 44 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=9.365
+ $Y=2.715 $X2=9.6 $Y2=2.86
r101 3 39 600 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=5.62
+ $Y=2.715 $X2=5.855 $Y2=3.57
r102 2 28 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=2.26
+ $Y=2.815 $X2=2.385 $Y2=3.025
r103 1 19 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.915
+ $Y=2.795 $X2=1.055 $Y2=2.92
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%A_605_563# 1 2 9 11 15 16 18
c39 18 0 1.70347e-19 $X=3.95 $Y=2.11
r40 17 18 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=3.95 $Y=1.025
+ $X2=3.95 $Y2=2.11
r41 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.865 $Y=2.195
+ $X2=3.95 $Y2=2.11
r42 15 16 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.865 $Y=2.195
+ $X2=3.33 $Y2=2.195
r43 11 17 8.45803 $w=4.1e-07 $l=2.43824e-07 $layer=LI1_cond $X=3.865 $Y=0.82
+ $X2=3.95 $Y2=1.025
r44 11 13 11.3839 $w=4.08e-07 $l=4.05e-07 $layer=LI1_cond $X=3.865 $Y=0.82
+ $X2=3.46 $Y2=0.82
r45 7 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.165 $Y=2.28
+ $X2=3.33 $Y2=2.195
r46 7 9 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=3.165 $Y=2.28
+ $X2=3.165 $Y2=3
r47 2 9 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=3.025
+ $Y=2.815 $X2=3.165 $Y2=3
r48 1 13 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.565 $X2=3.46 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%Q 1 2 7 8 9 10 11 12 13 36
r14 33 36 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=11.725 $Y=2.35
+ $X2=11.725 $Y2=2.36
r15 13 43 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=11.725 $Y=3.145
+ $X2=11.725 $Y2=3.57
r16 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=11.725 $Y=2.775
+ $X2=11.725 $Y2=3.145
r17 11 33 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=11.725 $Y=2.335
+ $X2=11.725 $Y2=2.35
r18 11 46 5.94304 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=11.725 $Y=2.335
+ $X2=11.725 $Y2=2.185
r19 11 12 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=11.725 $Y=2.42
+ $X2=11.725 $Y2=2.775
r20 11 36 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=11.725 $Y=2.42
+ $X2=11.725 $Y2=2.36
r21 10 46 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=11.765 $Y=2.035
+ $X2=11.765 $Y2=2.185
r22 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=11.765 $Y=1.665
+ $X2=11.765 $Y2=2.035
r23 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=11.765 $Y=1.295
+ $X2=11.765 $Y2=1.665
r24 7 8 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=11.765 $Y=0.85
+ $X2=11.765 $Y2=1.295
r25 2 43 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=11.585
+ $Y=2.215 $X2=11.725 $Y2=3.57
r26 2 36 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=11.585
+ $Y=2.215 $X2=11.725 $Y2=2.36
r27 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.585
+ $Y=0.705 $X2=11.725 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_HVL__DFXTP_1%VGND 1 2 3 4 5 16 19 28 35 44 53 54
r91 53 57 7.09538 $w=5.88e-07 $l=3.5e-07 $layer=LI1_cond $X=10.985 $Y=0.48
+ $X2=10.985 $Y2=0.83
r92 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.165 $Y=0.48
+ $X2=11.165 $Y2=0.48
r93 48 54 0.595053 $w=3.7e-07 $l=1.55e-06 $layer=MET1_cond $X=9.615 $Y=0.44
+ $X2=11.165 $Y2=0.44
r94 45 48 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=8.895 $Y=0.44
+ $X2=9.615 $Y2=0.44
r95 44 50 2.95368 $w=9.48e-07 $l=2.3e-07 $layer=LI1_cond $X=9.255 $Y=0.48
+ $X2=9.255 $Y2=0.71
r96 44 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.615 $Y=0.48
+ $X2=9.615 $Y2=0.48
r97 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.895 $Y=0.48
+ $X2=8.895 $Y2=0.48
r98 39 45 1.07685 $w=3.7e-07 $l=2.805e-06 $layer=MET1_cond $X=6.09 $Y=0.44
+ $X2=8.895 $Y2=0.44
r99 35 41 4.10947 $w=9.48e-07 $l=3.2e-07 $layer=LI1_cond $X=5.73 $Y=0.48
+ $X2=5.73 $Y2=0.8
r100 35 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.09 $Y=0.48
+ $X2=6.09 $Y2=0.48
r101 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.37 $Y=0.48
+ $X2=5.37 $Y2=0.48
r102 29 36 1.04038 $w=3.7e-07 $l=2.71e-06 $layer=MET1_cond $X=2.66 $Y=0.44
+ $X2=5.37 $Y2=0.44
r103 28 32 6.24501 $w=5.63e-07 $l=2.95e-07 $layer=LI1_cond $X=2.482 $Y=0.48
+ $X2=2.482 $Y2=0.775
r104 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.66 $Y=0.48
+ $X2=2.66 $Y2=0.48
r105 23 29 0.48564 $w=3.7e-07 $l=1.265e-06 $layer=MET1_cond $X=1.395 $Y=0.44
+ $X2=2.66 $Y2=0.44
r106 20 23 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.675 $Y=0.44
+ $X2=1.395 $Y2=0.44
r107 19 25 4.68737 $w=9.48e-07 $l=3.65e-07 $layer=LI1_cond $X=1.035 $Y=0.48
+ $X2=1.035 $Y2=0.845
r108 19 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.395 $Y=0.48
+ $X2=1.395 $Y2=0.48
r109 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.675 $Y=0.48
+ $X2=0.675 $Y2=0.48
r110 16 39 0.0345515 $w=3.7e-07 $l=9e-08 $layer=MET1_cond $X=6 $Y=0.44 $X2=6.09
+ $Y2=0.44
r111 16 36 0.24186 $w=3.7e-07 $l=6.3e-07 $layer=MET1_cond $X=6 $Y=0.44 $X2=5.37
+ $Y2=0.44
r112 5 57 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=10.8
+ $Y=0.705 $X2=10.945 $Y2=0.83
r113 4 50 91 $w=1.7e-07 $l=4.87134e-07 $layer=licon1_NDIFF $count=2 $X=9.145
+ $Y=0.565 $X2=9.565 $Y2=0.71
r114 3 41 182 $w=1.7e-07 $l=3.53483e-07 $layer=licon1_NDIFF $count=1 $X=5.785
+ $Y=0.565 $X2=6.04 $Y2=0.8
r115 2 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.565 $X2=2.56 $Y2=0.775
r116 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.935
+ $Y=0.635 $X2=1.075 $Y2=0.845
.ends

