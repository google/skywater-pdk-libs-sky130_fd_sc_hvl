* File: sky130_fd_sc_hvl__nor3_1.pex.spice
* Created: Wed Sep  2 09:08:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__NOR3_1%VNB 5 7 17 24
r23 11 24 0.769925 $w=2.3e-07 $l=1.2e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.44
+ $Y2=0
r24 7 17 0.92391 $w=2.3e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r25 7 24 0.153985 $w=2.3e-07 $l=2.4e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.44
+ $Y2=0
r26 5 17 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r27 5 11 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR3_1%VPB 4 6 14 15 21
r22 14 15 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=4.07
+ $X2=3.12 $Y2=4.07
r23 10 21 0.769925 $w=2.3e-07 $l=1.2e-06 $layer=MET1_cond $X=0.24 $Y=4.07
+ $X2=1.44 $Y2=4.07
r24 9 14 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=3.12 $Y2=4.07
r25 9 10 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r26 6 15 0.92391 $w=2.3e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=4.07
+ $X2=3.12 $Y2=4.07
r27 6 21 0.153985 $w=2.3e-07 $l=2.4e-07 $layer=MET1_cond $X=1.68 $Y=4.07
+ $X2=1.44 $Y2=4.07
r28 4 14 52 $w=1.7e-07 $l=3.16221e-06 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=3.12 $Y2=4.07
r29 4 9 52 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=3 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR3_1%A 3 7 9 10 18
r26 17 18 7.49041 $w=5e-07 $l=7e-08 $layer=POLY_cond $X=0.705 $Y=1.665 $X2=0.775
+ $Y2=1.665
r27 14 17 44.4074 $w=5e-07 $l=4.15e-07 $layer=POLY_cond $X=0.29 $Y=1.665
+ $X2=0.705 $Y2=1.665
r28 9 10 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.275 $Y=1.665
+ $X2=0.275 $Y2=2.035
r29 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.69 $X2=0.29 $Y2=1.69
r30 5 18 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.775 $Y=1.915
+ $X2=0.775 $Y2=1.665
r31 5 7 112.356 $w=5e-07 $l=1.05e-06 $layer=POLY_cond $X=0.775 $Y=1.915
+ $X2=0.775 $Y2=2.965
r32 1 17 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.705 $Y=1.415
+ $X2=0.705 $Y2=1.665
r33 1 3 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.705 $Y=1.415 $X2=0.705
+ $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR3_1%B 1 2 3 8 14
r28 11 14 115.031 $w=5e-07 $l=1.075e-06 $layer=POLY_cond $X=1.485 $Y=1.89
+ $X2=1.485 $Y2=2.965
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.89 $X2=1.42 $Y2=1.89
r30 8 11 104.866 $w=5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.485 $Y=0.91 $X2=1.485
+ $Y2=1.89
r31 3 12 8.68508 $w=3.43e-07 $l=2.6e-07 $layer=LI1_cond $X=1.68 $Y=1.947
+ $X2=1.42 $Y2=1.947
r32 2 12 7.34891 $w=3.43e-07 $l=2.2e-07 $layer=LI1_cond $X=1.2 $Y=1.947 $X2=1.42
+ $Y2=1.947
r33 1 2 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.947 $X2=1.2
+ $Y2=1.947
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR3_1%C 3 6 8 9 10 11 17 18 20
r26 17 20 21.1255 $w=5.7e-07 $l=2.15e-07 $layer=POLY_cond $X=2.23 $Y=1.89
+ $X2=2.23 $Y2=2.105
r27 17 19 27.696 $w=5.7e-07 $l=2.85e-07 $layer=POLY_cond $X=2.23 $Y=1.89
+ $X2=2.23 $Y2=1.605
r28 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.89 $X2=2.14 $Y2=1.89
r29 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.14 $Y=2.775
+ $X2=2.14 $Y2=3.145
r30 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.14 $Y=2.405
+ $X2=2.14 $Y2=2.775
r31 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.14 $Y=2.035 $X2=2.14
+ $Y2=2.405
r32 8 18 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.14 $Y=2.035
+ $X2=2.14 $Y2=1.89
r33 6 19 74.3691 $w=5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.265 $Y=0.91
+ $X2=2.265 $Y2=1.605
r34 3 20 82.904 $w=5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.195 $Y=2.965 $X2=2.195
+ $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR3_1%VPWR 1 4 7 19
r20 11 19 0.474123 $w=3.7e-07 $l=1.235e-06 $layer=MET1_cond $X=0.205 $Y=3.63
+ $X2=1.44 $Y2=3.63
r21 10 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.205 $Y=3.59
+ $X2=0.205 $Y2=3.59
r22 7 10 8.80299 $w=1.668e-06 $l=1.205e-06 $layer=LI1_cond $X=0.925 $Y=2.385
+ $X2=0.925 $Y2=3.59
r23 4 19 0.0787006 $w=3.7e-07 $l=2.05e-07 $layer=MET1_cond $X=1.645 $Y=3.63
+ $X2=1.44 $Y2=3.63
r24 4 10 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.645 $Y=3.59
+ $X2=1.645 $Y2=3.59
r25 1 10 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.24
+ $Y=2.215 $X2=0.385 $Y2=3.59
r26 1 7 300 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=2 $X=0.24
+ $Y=2.215 $X2=0.385 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR3_1%Y 1 2 3 12 14 15 18 20 21 22 23 24 33
r38 31 33 3.04419 $w=2.63e-07 $l=7e-08 $layer=LI1_cond $X=2.622 $Y=1.595
+ $X2=2.622 $Y2=1.665
r39 24 45 19.3523 $w=2.63e-07 $l=4.45e-07 $layer=LI1_cond $X=2.622 $Y=3.145
+ $X2=2.622 $Y2=3.59
r40 23 24 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=2.622 $Y=2.775
+ $X2=2.622 $Y2=3.145
r41 22 23 18.9175 $w=2.63e-07 $l=4.35e-07 $layer=LI1_cond $X=2.622 $Y=2.34
+ $X2=2.622 $Y2=2.775
r42 21 22 13.264 $w=2.63e-07 $l=3.05e-07 $layer=LI1_cond $X=2.622 $Y=2.035
+ $X2=2.622 $Y2=2.34
r43 20 31 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.622 $Y=1.51
+ $X2=2.622 $Y2=1.595
r44 20 21 15.7863 $w=2.63e-07 $l=3.63e-07 $layer=LI1_cond $X=2.622 $Y=1.672
+ $X2=2.622 $Y2=2.035
r45 20 33 0.304419 $w=2.63e-07 $l=7e-09 $layer=LI1_cond $X=2.622 $Y=1.672
+ $X2=2.622 $Y2=1.665
r46 16 20 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.622 $Y=1.425
+ $X2=2.622 $Y2=1.51
r47 16 18 32.3989 $w=2.63e-07 $l=7.45e-07 $layer=LI1_cond $X=2.622 $Y=1.425
+ $X2=2.622 $Y2=0.68
r48 14 20 2.98021 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.49 $Y=1.51
+ $X2=2.622 $Y2=1.51
r49 14 15 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=2.49 $Y=1.51
+ $X2=1.18 $Y2=1.51
r50 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.055 $Y=1.425
+ $X2=1.18 $Y2=1.51
r51 10 12 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=1.055 $Y=1.425
+ $X2=1.055 $Y2=0.66
r52 3 45 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.445
+ $Y=2.215 $X2=2.585 $Y2=3.59
r53 3 22 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.445
+ $Y=2.215 $X2=2.585 $Y2=2.34
r54 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.515
+ $Y=0.535 $X2=2.655 $Y2=0.68
r55 1 12 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.955
+ $Y=0.535 $X2=1.095 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__NOR3_1%VGND 1 2 7 10 17 21 28
r25 17 23 2.31158 $w=9.48e-07 $l=1.8e-07 $layer=LI1_cond $X=1.835 $Y=0.48
+ $X2=1.835 $Y2=0.66
r26 17 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.195 $Y=0.48
+ $X2=2.195 $Y2=0.48
r27 17 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.475 $Y=0.48
+ $X2=1.475 $Y2=0.48
r28 11 28 0.335917 $w=3.7e-07 $l=8.75e-07 $layer=MET1_cond $X=0.565 $Y=0.44
+ $X2=1.44 $Y2=0.44
r29 10 14 4.0545 $w=5.88e-07 $l=2e-07 $layer=LI1_cond $X=0.385 $Y=0.48 $X2=0.385
+ $Y2=0.68
r30 10 11 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.565 $Y=0.48
+ $X2=0.565 $Y2=0.48
r31 7 21 0.197711 $w=3.7e-07 $l=5.15e-07 $layer=MET1_cond $X=1.68 $Y=0.44
+ $X2=2.195 $Y2=0.44
r32 7 28 0.0921373 $w=3.7e-07 $l=2.4e-07 $layer=MET1_cond $X=1.68 $Y=0.44
+ $X2=1.44 $Y2=0.44
r33 2 23 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.735
+ $Y=0.535 $X2=1.875 $Y2=0.66
r34 1 14 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.19
+ $Y=0.535 $X2=0.315 $Y2=0.68
.ends

