* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
X0 a_1096_491# a_1138_81# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X1 a_775_491# a_345_107# a_917_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X2 a_1096_107# a_1138_81# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X3 a_917_107# a_462_107# a_1096_491# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X4 a_775_107# a_462_107# a_917_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X5 VPWR a_917_107# a_1138_81# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X6 a_462_107# a_345_107# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X7 a_1138_81# a_917_107# a_1512_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X8 a_917_107# a_345_107# a_1096_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X9 a_462_107# a_345_107# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X10 VPWR a_1138_81# Q VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 a_1138_81# RESET_B VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X12 a_32_107# D VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X13 VPWR a_32_107# a_775_491# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X14 VGND GATE a_345_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X15 a_32_107# D VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X16 VGND a_32_107# a_775_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X17 VGND a_1138_81# Q VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 VPWR GATE a_345_107# VPB sky130_fd_pr__pfet_g5v0d10v5 w=750000u l=500000u
X19 a_1512_107# RESET_B VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
.ends
