* File: sky130_fd_sc_hvl__sdfrbp_1.pxi.spice
* Created: Fri Aug 28 09:39:44 2020
* 
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%VNB N_VNB_M1029_b VNB N_VNB_c_3_p
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%VNB
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%VPB N_VPB_M1018_b VPB N_VPB_c_151_p
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%VPB
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%SCE N_SCE_M1018_g N_SCE_M1016_g N_SCE_c_378_n
+ N_SCE_M1031_g N_SCE_c_379_n N_SCE_c_360_n N_SCE_c_362_n N_SCE_c_364_n
+ N_SCE_c_365_n N_SCE_c_380_n N_SCE_c_366_n N_SCE_c_387_p N_SCE_c_381_n SCE SCE
+ N_SCE_M1029_g N_SCE_c_383_n N_SCE_c_370_n N_SCE_c_371_n
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%SCE
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%D N_D_c_484_n N_D_M1001_g N_D_M1040_g D
+ N_D_c_487_n PM_SKY130_FD_SC_HVL__SDFRBP_1%D
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%A_222_131# N_A_222_131#_M1029_d
+ N_A_222_131#_M1018_d N_A_222_131#_M1041_g N_A_222_131#_c_529_n
+ N_A_222_131#_M1006_g N_A_222_131#_c_524_n N_A_222_131#_c_525_n
+ N_A_222_131#_c_526_n N_A_222_131#_c_534_n N_A_222_131#_c_535_n
+ N_A_222_131#_c_538_n N_A_222_131#_c_527_n N_A_222_131#_c_528_n
+ N_A_222_131#_c_540_n N_A_222_131#_c_575_n N_A_222_131#_c_541_n
+ N_A_222_131#_c_542_n N_A_222_131#_c_606_p N_A_222_131#_c_543_n
+ N_A_222_131#_c_544_n N_A_222_131#_c_545_n N_A_222_131#_c_546_n
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%A_222_131#
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%SCD N_SCD_c_659_n N_SCD_M1033_g N_SCD_c_662_n
+ N_SCD_c_663_n N_SCD_c_664_n N_SCD_c_665_n SCD SCD N_SCD_M1035_g N_SCD_c_682_n
+ N_SCD_c_667_n PM_SKY130_FD_SC_HVL__SDFRBP_1%SCD
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%CLK N_CLK_M1026_g N_CLK_M1002_g CLK
+ N_CLK_c_726_n N_CLK_c_733_p PM_SKY130_FD_SC_HVL__SDFRBP_1%CLK
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%A_1569_126# N_A_1569_126#_M1000_d
+ N_A_1569_126#_M1019_d N_A_1569_126#_c_781_n N_A_1569_126#_M1017_g
+ N_A_1569_126#_M1028_g N_A_1569_126#_c_760_n N_A_1569_126#_c_761_n
+ N_A_1569_126#_c_762_n N_A_1569_126#_c_764_n N_A_1569_126#_c_766_n
+ N_A_1569_126#_c_810_p N_A_1569_126#_c_767_n N_A_1569_126#_c_828_p
+ N_A_1569_126#_c_768_n N_A_1569_126#_c_770_n N_A_1569_126#_c_801_p
+ N_A_1569_126#_c_772_n N_A_1569_126#_c_774_n N_A_1569_126#_c_786_n
+ N_A_1569_126#_c_775_n N_A_1569_126#_c_787_n N_A_1569_126#_c_872_p
+ N_A_1569_126#_c_776_n N_A_1569_126#_c_804_p N_A_1569_126#_c_778_n
+ N_A_1569_126#_M1004_g N_A_1569_126#_M1011_g N_A_1569_126#_c_780_n
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%A_1569_126#
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%A_1290_126# N_A_1290_126#_M1026_d
+ N_A_1290_126#_M1002_d N_A_1290_126#_M1000_g N_A_1290_126#_M1019_g
+ N_A_1290_126#_c_948_n N_A_1290_126#_c_949_n N_A_1290_126#_M1027_g
+ N_A_1290_126#_c_950_n N_A_1290_126#_M1037_g N_A_1290_126#_M1024_g
+ N_A_1290_126#_c_951_n N_A_1290_126#_c_952_n N_A_1290_126#_M1020_g
+ N_A_1290_126#_c_954_n N_A_1290_126#_c_955_n N_A_1290_126#_c_957_n
+ N_A_1290_126#_c_958_n N_A_1290_126#_c_974_n N_A_1290_126#_c_975_n
+ N_A_1290_126#_c_959_n N_A_1290_126#_c_960_n N_A_1290_126#_c_978_n
+ N_A_1290_126#_c_961_n N_A_1290_126#_c_1011_n N_A_1290_126#_c_1012_n
+ N_A_1290_126#_c_979_n N_A_1290_126#_c_1031_p N_A_1290_126#_c_962_n
+ N_A_1290_126#_c_963_n N_A_1290_126#_c_964_n
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%A_1290_126#
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%A_2014_537# N_A_2014_537#_M1039_d
+ N_A_2014_537#_M1003_d N_A_2014_537#_M1038_g N_A_2014_537#_c_1170_n
+ N_A_2014_537#_c_1171_n N_A_2014_537#_c_1163_n N_A_2014_537#_c_1164_n
+ N_A_2014_537#_c_1183_n N_A_2014_537#_c_1165_n N_A_2014_537#_c_1166_n
+ N_A_2014_537#_c_1167_n N_A_2014_537#_c_1177_n N_A_2014_537#_c_1180_n
+ N_A_2014_537#_c_1181_n N_A_2014_537#_c_1194_n N_A_2014_537#_c_1195_n
+ N_A_2014_537#_c_1168_n N_A_2014_537#_M1005_g
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%A_2014_537#
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%RESET_B N_RESET_B_M1012_g N_RESET_B_M1007_g
+ N_RESET_B_c_1286_n N_RESET_B_c_1287_n N_RESET_B_M1013_g N_RESET_B_c_1301_n
+ N_RESET_B_M1034_g N_RESET_B_c_1302_n N_RESET_B_c_1305_n N_RESET_B_c_1289_n
+ RESET_B RESET_B N_RESET_B_c_1308_n N_RESET_B_c_1309_n N_RESET_B_c_1310_n
+ N_RESET_B_c_1311_n N_RESET_B_c_1312_n N_RESET_B_c_1291_n N_RESET_B_M1008_g
+ N_RESET_B_c_1293_n N_RESET_B_M1014_g N_RESET_B_c_1296_n N_RESET_B_c_1297_n
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%RESET_B
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%A_1816_659# N_A_1816_659#_M1027_d
+ N_A_1816_659#_M1017_d N_A_1816_659#_M1013_d N_A_1816_659#_M1039_g
+ N_A_1816_659#_M1003_g N_A_1816_659#_c_1500_n N_A_1816_659#_c_1507_n
+ N_A_1816_659#_c_1510_n N_A_1816_659#_c_1511_n N_A_1816_659#_c_1512_n
+ N_A_1816_659#_c_1515_n N_A_1816_659#_c_1501_n N_A_1816_659#_c_1516_n
+ N_A_1816_659#_c_1517_n PM_SKY130_FD_SC_HVL__SDFRBP_1%A_1816_659#
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%A_2841_81# N_A_2841_81#_M1015_d
+ N_A_2841_81#_M1034_d N_A_2841_81#_M1030_g N_A_2841_81#_M1025_g
+ N_A_2841_81#_c_1618_n N_A_2841_81#_c_1620_n N_A_2841_81#_c_1625_n
+ N_A_2841_81#_c_1626_n N_A_2841_81#_c_1627_n N_A_2841_81#_c_1628_n
+ N_A_2841_81#_c_1669_p N_A_2841_81#_c_1629_n N_A_2841_81#_c_1621_n
+ N_A_2841_81#_c_1630_n N_A_2841_81#_c_1622_n N_A_2841_81#_c_1624_n
+ N_A_2841_81#_c_1632_n PM_SKY130_FD_SC_HVL__SDFRBP_1%A_2841_81#
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%A_2624_107# N_A_2624_107#_M1028_d
+ N_A_2624_107#_M1024_d N_A_2624_107#_c_1714_n N_A_2624_107#_M1015_g
+ N_A_2624_107#_M1021_g N_A_2624_107#_M1032_g N_A_2624_107#_c_1716_n
+ N_A_2624_107#_M1023_g N_A_2624_107#_c_1718_n N_A_2624_107#_c_1719_n
+ N_A_2624_107#_M1036_g N_A_2624_107#_M1009_g N_A_2624_107#_c_1722_n
+ N_A_2624_107#_c_1723_n N_A_2624_107#_c_1724_n N_A_2624_107#_c_1725_n
+ N_A_2624_107#_c_1736_n N_A_2624_107#_c_1739_n N_A_2624_107#_c_1752_n
+ N_A_2624_107#_c_1726_n N_A_2624_107#_c_1727_n N_A_2624_107#_c_1756_n
+ N_A_2624_107#_c_1757_n N_A_2624_107#_c_1789_n
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%A_2624_107#
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%A_3613_443# N_A_3613_443#_M1009_s
+ N_A_3613_443#_M1036_s N_A_3613_443#_M1022_g N_A_3613_443#_M1010_g
+ N_A_3613_443#_c_1879_n N_A_3613_443#_c_1885_n N_A_3613_443#_c_1880_n
+ N_A_3613_443#_c_1881_n N_A_3613_443#_c_1888_n
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%A_3613_443#
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%VPWR N_VPWR_M1018_s N_VPWR_M1016_d
+ N_VPWR_M1012_d N_VPWR_M1019_s N_VPWR_M1038_d N_VPWR_M1003_s N_VPWR_M1025_d
+ N_VPWR_M1021_d N_VPWR_M1036_d VPWR N_VPWR_c_1922_n N_VPWR_c_1925_n
+ N_VPWR_c_1928_n N_VPWR_c_1931_n N_VPWR_c_1934_n N_VPWR_c_1937_n
+ N_VPWR_c_1940_n N_VPWR_c_1943_n N_VPWR_c_1946_n N_VPWR_c_1949_n
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%VPWR
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%A_339_655# N_A_339_655#_M1041_d
+ N_A_339_655#_M1027_s N_A_339_655#_M1001_s N_A_339_655#_M1006_d
+ N_A_339_655#_M1017_s N_A_339_655#_c_2087_n N_A_339_655#_c_2088_n
+ N_A_339_655#_c_2080_n N_A_339_655#_c_2091_n N_A_339_655#_c_2081_n
+ N_A_339_655#_c_2095_n N_A_339_655#_c_2159_n N_A_339_655#_c_2096_n
+ N_A_339_655#_c_2099_n N_A_339_655#_c_2101_n N_A_339_655#_c_2082_n
+ N_A_339_655#_c_2083_n N_A_339_655#_c_2104_n N_A_339_655#_c_2105_n
+ N_A_339_655#_c_2107_n N_A_339_655#_c_2109_n N_A_339_655#_c_2084_n
+ N_A_339_655#_c_2085_n N_A_339_655#_c_2111_n N_A_339_655#_c_2112_n
+ N_A_339_655#_c_2086_n PM_SKY130_FD_SC_HVL__SDFRBP_1%A_339_655#
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%Q_N N_Q_N_M1023_d N_Q_N_M1032_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_2263_n PM_SKY130_FD_SC_HVL__SDFRBP_1%Q_N
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%Q N_Q_M1010_d N_Q_M1022_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%Q
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%VGND N_VGND_M1029_s N_VGND_M1007_d
+ N_VGND_M1000_s N_VGND_M1008_d N_VGND_M1030_d N_VGND_M1023_s N_VGND_M1009_d
+ VGND N_VGND_c_2294_n N_VGND_c_2296_n N_VGND_c_2298_n N_VGND_c_2300_n
+ N_VGND_c_2302_n N_VGND_c_2304_n N_VGND_c_2306_n N_VGND_c_2308_n
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%VGND
x_PM_SKY130_FD_SC_HVL__SDFRBP_1%noxref_25 N_noxref_25_M1040_s
+ N_noxref_25_M1035_d N_noxref_25_c_2431_n N_noxref_25_c_2432_n
+ N_noxref_25_c_2434_n N_noxref_25_c_2436_n
+ PM_SKY130_FD_SC_HVL__SDFRBP_1%noxref_25
cc_1 N_VNB_M1029_b N_SCE_M1031_g 0.0397909f $X=-0.33 $Y=-0.265 $X2=3.83
+ $Y2=0.745
cc_2 N_VNB_M1029_b N_SCE_c_360_n 0.0583843f $X=-0.33 $Y=-0.265 $X2=1.515
+ $Y2=0.35
cc_3 N_VNB_c_3_p N_SCE_c_360_n 0.00235285f $X=0.24 $Y=0 $X2=1.515 $Y2=0.35
cc_4 N_VNB_M1029_b N_SCE_c_362_n 0.0141601f $X=-0.33 $Y=-0.265 $X2=0.985
+ $Y2=0.35
cc_5 N_VNB_c_3_p N_SCE_c_362_n 5.63772e-19 $X=0.24 $Y=0 $X2=0.985 $Y2=0.35
cc_6 N_VNB_M1029_b N_SCE_c_364_n 0.0177304f $X=-0.33 $Y=-0.265 $X2=1.6 $Y2=1.275
cc_7 N_VNB_M1029_b N_SCE_c_365_n 0.00546025f $X=-0.33 $Y=-0.265 $X2=1.685
+ $Y2=1.36
cc_8 N_VNB_M1029_b N_SCE_c_366_n 0.00104405f $X=-0.33 $Y=-0.265 $X2=0.82
+ $Y2=1.295
cc_9 N_VNB_M1029_b SCE 0.00867222f $X=-0.33 $Y=-0.265 $X2=3.995 $Y2=1.58
cc_10 N_VNB_M1029_b N_SCE_M1029_g 0.139338f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=0.865
cc_11 N_VNB_c_3_p N_SCE_M1029_g 7.4229e-19 $X=0.24 $Y=0 $X2=0.86 $Y2=0.865
cc_12 N_VNB_M1029_b N_SCE_c_370_n 0.0807578f $X=-0.33 $Y=-0.265 $X2=3.765
+ $Y2=1.365
cc_13 N_VNB_M1029_b N_SCE_c_371_n 0.0407298f $X=-0.33 $Y=-0.265 $X2=3.485
+ $Y2=1.535
cc_14 N_VNB_M1029_b N_D_c_484_n 0.0674252f $X=-0.33 $Y=-0.265 $X2=0.86 $Y2=3.115
cc_15 N_VNB_M1029_b N_D_M1001_g 0.0109105f $X=-0.33 $Y=-0.265 $X2=0.86 $Y2=3.455
cc_16 N_VNB_M1029_b N_D_M1040_g 0.0491756f $X=-0.33 $Y=-0.265 $X2=2.94 $Y2=3.485
cc_17 N_VNB_M1029_b N_D_c_487_n 0.0082589f $X=-0.33 $Y=-0.265 $X2=3.83 $Y2=0.745
cc_18 N_VNB_M1029_b N_A_222_131#_M1041_g 0.0447569f $X=-0.33 $Y=-0.265 $X2=3.385
+ $Y2=1.89
cc_19 N_VNB_M1029_b N_A_222_131#_c_524_n 0.0148955f $X=-0.33 $Y=-0.265 $X2=0.82
+ $Y2=1.46
cc_20 N_VNB_M1029_b N_A_222_131#_c_525_n 0.0265527f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_21 N_VNB_M1029_b N_A_222_131#_c_526_n 0.0210341f $X=-0.33 $Y=-0.265 $X2=0.9
+ $Y2=1.295
cc_22 N_VNB_M1029_b N_A_222_131#_c_527_n 6.60714e-19 $X=-0.33 $Y=-0.265 $X2=0.82
+ $Y2=1.295
cc_23 N_VNB_M1029_b N_A_222_131#_c_528_n 0.020099f $X=-0.33 $Y=-0.265 $X2=1.64
+ $Y2=2.75
cc_24 N_VNB_M1029_b N_SCD_M1035_g 0.108951f $X=-0.33 $Y=-0.265 $X2=0.82 $Y2=1.46
cc_25 N_VNB_M1029_b N_CLK_M1026_g 0.0879884f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=3.455
cc_26 N_VNB_M1029_b N_CLK_c_726_n 0.0184059f $X=-0.33 $Y=-0.265 $X2=3.83
+ $Y2=0.745
cc_27 N_VNB_M1029_b N_A_1569_126#_c_760_n 0.00676569f $X=-0.33 $Y=-0.265
+ $X2=1.11 $Y2=2.865
cc_28 N_VNB_M1029_b N_A_1569_126#_c_761_n 0.00778358f $X=-0.33 $Y=-0.265
+ $X2=0.82 $Y2=1.46
cc_29 N_VNB_M1029_b N_A_1569_126#_c_762_n 0.128062f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_30 N_VNB_c_3_p N_A_1569_126#_c_762_n 0.00808919f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_31 N_VNB_M1029_b N_A_1569_126#_c_764_n 0.0171312f $X=-0.33 $Y=-0.265 $X2=0.82
+ $Y2=1.46
cc_32 N_VNB_c_3_p N_A_1569_126#_c_764_n 0.00120299f $X=0.24 $Y=0 $X2=0.82
+ $Y2=1.46
cc_33 N_VNB_M1029_b N_A_1569_126#_c_766_n 0.00164526f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_M1029_b N_A_1569_126#_c_767_n 0.0108199f $X=-0.33 $Y=-0.265 $X2=1.6
+ $Y2=1.275
cc_35 N_VNB_M1029_b N_A_1569_126#_c_768_n 0.0480975f $X=-0.33 $Y=-0.265
+ $X2=2.875 $Y2=2.75
cc_36 N_VNB_c_3_p N_A_1569_126#_c_768_n 0.00229582f $X=0.24 $Y=0 $X2=2.875
+ $Y2=2.75
cc_37 N_VNB_M1029_b N_A_1569_126#_c_770_n 0.0135505f $X=-0.33 $Y=-0.265
+ $X2=2.875 $Y2=2.75
cc_38 N_VNB_c_3_p N_A_1569_126#_c_770_n 5.63772e-19 $X=0.24 $Y=0 $X2=2.875
+ $Y2=2.75
cc_39 N_VNB_M1029_b N_A_1569_126#_c_772_n 0.0940638f $X=-0.33 $Y=-0.265 $X2=0.82
+ $Y2=1.295
cc_40 N_VNB_c_3_p N_A_1569_126#_c_772_n 0.00429538f $X=0.24 $Y=0 $X2=0.82
+ $Y2=1.295
cc_41 N_VNB_M1029_b N_A_1569_126#_c_774_n 0.0103952f $X=-0.33 $Y=-0.265 $X2=1.6
+ $Y2=2.83
cc_42 N_VNB_M1029_b N_A_1569_126#_c_775_n 0.0011164f $X=-0.33 $Y=-0.265
+ $X2=3.515 $Y2=1.58
cc_43 N_VNB_M1029_b N_A_1569_126#_c_776_n 0.0121104f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=1.46
cc_44 N_VNB_c_3_p N_A_1569_126#_c_776_n 5.63772e-19 $X=0.24 $Y=0 $X2=0.86
+ $Y2=1.46
cc_45 N_VNB_M1029_b N_A_1569_126#_c_778_n 0.0497584f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_M1029_b N_A_1569_126#_M1004_g 0.0887996f $X=-0.33 $Y=-0.265
+ $X2=3.385 $Y2=1.89
cc_47 N_VNB_M1029_b N_A_1569_126#_c_780_n 0.0369337f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_M1029_b N_A_1290_126#_M1019_g 0.0139856f $X=-0.33 $Y=-0.265 $X2=3.83
+ $Y2=0.745
cc_49 N_VNB_M1029_b N_A_1290_126#_c_948_n 0.0811246f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_M1029_b N_A_1290_126#_c_949_n 0.0256957f $X=-0.33 $Y=-0.265 $X2=1.11
+ $Y2=2.865
cc_51 N_VNB_M1029_b N_A_1290_126#_c_950_n 0.0269137f $X=-0.33 $Y=-0.265 $X2=0.82
+ $Y2=1.46
cc_52 N_VNB_M1029_b N_A_1290_126#_c_951_n 0.0256824f $X=-0.33 $Y=-0.265
+ $X2=3.485 $Y2=1.36
cc_53 N_VNB_M1029_b N_A_1290_126#_c_952_n 0.0376263f $X=-0.33 $Y=-0.265
+ $X2=1.685 $Y2=1.36
cc_54 N_VNB_M1029_b N_A_1290_126#_M1020_g 0.0389036f $X=-0.33 $Y=-0.265
+ $X2=2.875 $Y2=2.75
cc_55 N_VNB_M1029_b N_A_1290_126#_c_954_n 0.0370784f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_56 N_VNB_M1029_b N_A_1290_126#_c_955_n 0.0216169f $X=-0.33 $Y=-0.265 $X2=1.64
+ $Y2=2.83
cc_57 N_VNB_c_3_p N_A_1290_126#_c_955_n 3.93713e-19 $X=0.24 $Y=0 $X2=1.64
+ $Y2=2.83
cc_58 N_VNB_M1029_b N_A_1290_126#_c_957_n 0.00762054f $X=-0.33 $Y=-0.265
+ $X2=3.515 $Y2=1.58
cc_59 N_VNB_M1029_b N_A_1290_126#_c_958_n 0.0233746f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_60 N_VNB_M1029_b N_A_1290_126#_c_959_n 0.00330679f $X=-0.33 $Y=-0.265 $X2=1.6
+ $Y2=2.865
cc_61 N_VNB_M1029_b N_A_1290_126#_c_960_n 0.00246458f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_62 N_VNB_M1029_b N_A_1290_126#_c_961_n 0.00289881f $X=-0.33 $Y=-0.265
+ $X2=3.765 $Y2=1.507
cc_63 N_VNB_M1029_b N_A_1290_126#_c_962_n 0.0709499f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_64 N_VNB_M1029_b N_A_1290_126#_c_963_n 0.0284118f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_65 N_VNB_M1029_b N_A_1290_126#_c_964_n 0.0210915f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_66 N_VNB_M1029_b N_A_2014_537#_c_1163_n 0.017617f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=2.615
cc_67 N_VNB_M1029_b N_A_2014_537#_c_1164_n 0.010626f $X=-0.33 $Y=-0.265 $X2=0.82
+ $Y2=1.46
cc_68 N_VNB_M1029_b N_A_2014_537#_c_1165_n 0.00488948f $X=-0.33 $Y=-0.265
+ $X2=1.515 $Y2=0.35
cc_69 N_VNB_M1029_b N_A_2014_537#_c_1166_n 0.00769552f $X=-0.33 $Y=-0.265
+ $X2=0.985 $Y2=0.35
cc_70 N_VNB_M1029_b N_A_2014_537#_c_1167_n 6.11752e-19 $X=-0.33 $Y=-0.265
+ $X2=1.6 $Y2=0.435
cc_71 N_VNB_M1029_b N_A_2014_537#_c_1168_n 0.00108211f $X=-0.33 $Y=-0.265
+ $X2=1.6 $Y2=2.83
cc_72 N_VNB_M1029_b N_A_2014_537#_M1005_g 0.0703972f $X=-0.33 $Y=-0.265
+ $X2=3.515 $Y2=1.58
cc_73 N_VNB_M1029_b N_RESET_B_M1007_g 0.0467052f $X=-0.33 $Y=-0.265 $X2=2.94
+ $Y2=3.485
cc_74 N_VNB_M1029_b N_RESET_B_c_1286_n 0.331115f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_75 N_VNB_M1029_b N_RESET_B_c_1287_n 0.198346f $X=-0.33 $Y=-0.265 $X2=3.385
+ $Y2=1.89
cc_76 N_VNB_c_3_p N_RESET_B_c_1287_n 0.0914134f $X=0.24 $Y=0 $X2=3.385 $Y2=1.89
cc_77 N_VNB_M1029_b N_RESET_B_c_1289_n 0.00961225f $X=-0.33 $Y=-0.265 $X2=1.515
+ $Y2=0.35
cc_78 N_VNB_M1029_b RESET_B 0.00577786f $X=-0.33 $Y=-0.265 $X2=1.6 $Y2=1.275
cc_79 N_VNB_M1029_b N_RESET_B_c_1291_n 0.0293522f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=0.865
cc_80 N_VNB_M1029_b N_RESET_B_M1008_g 0.108032f $X=-0.33 $Y=-0.265 $X2=1.6
+ $Y2=2.865
cc_81 N_VNB_M1029_b N_RESET_B_c_1293_n 0.00200463f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_82 N_VNB_M1029_b N_RESET_B_M1014_g 0.0949481f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_83 N_VNB_c_3_p N_RESET_B_M1014_g 4.23569e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_84 N_VNB_M1029_b N_RESET_B_c_1296_n 0.0449916f $X=-0.33 $Y=-0.265 $X2=3.6
+ $Y2=1.535
cc_85 N_VNB_M1029_b N_RESET_B_c_1297_n 0.00369986f $X=-0.33 $Y=-0.265 $X2=3.485
+ $Y2=1.535
cc_86 N_VNB_M1029_b N_A_1816_659#_M1039_g 0.0876876f $X=-0.33 $Y=-0.265 $X2=3.83
+ $Y2=0.745
cc_87 N_VNB_c_3_p N_A_1816_659#_M1039_g 6.44563e-19 $X=0.24 $Y=0 $X2=3.83
+ $Y2=0.745
cc_88 N_VNB_M1029_b N_A_1816_659#_c_1500_n 0.00971348f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_89 N_VNB_M1029_b N_A_1816_659#_c_1501_n 0.00101051f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_90 N_VNB_M1029_b N_A_2841_81#_c_1618_n 0.0399529f $X=-0.33 $Y=-0.265 $X2=0.86
+ $Y2=2.615
cc_91 N_VNB_c_3_p N_A_2841_81#_c_1618_n 8.42484e-19 $X=0.24 $Y=0 $X2=0.86
+ $Y2=2.615
cc_92 N_VNB_M1029_b N_A_2841_81#_c_1620_n 0.0562197f $X=-0.33 $Y=-0.265 $X2=1.11
+ $Y2=2.865
cc_93 N_VNB_M1029_b N_A_2841_81#_c_1621_n 0.00918305f $X=-0.33 $Y=-0.265
+ $X2=1.765 $Y2=2.75
cc_94 N_VNB_M1029_b N_A_2841_81#_c_1622_n 0.015773f $X=-0.33 $Y=-0.265 $X2=0.82
+ $Y2=1.295
cc_95 N_VNB_c_3_p N_A_2841_81#_c_1622_n 8.97088e-19 $X=0.24 $Y=0 $X2=0.82
+ $Y2=1.295
cc_96 N_VNB_M1029_b N_A_2841_81#_c_1624_n 0.019429f $X=-0.33 $Y=-0.265 $X2=1.64
+ $Y2=2.83
cc_97 N_VNB_M1029_b N_A_2624_107#_c_1714_n 0.0512876f $X=-0.33 $Y=-0.265
+ $X2=2.94 $Y2=3.485
cc_98 N_VNB_c_3_p N_A_2624_107#_c_1714_n 0.0023273f $X=0.24 $Y=0 $X2=2.94
+ $Y2=3.485
cc_99 N_VNB_M1029_b N_A_2624_107#_c_1716_n 0.0495382f $X=-0.33 $Y=-0.265
+ $X2=0.82 $Y2=1.46
cc_100 N_VNB_c_3_p N_A_2624_107#_c_1716_n 0.00128467f $X=0.24 $Y=0 $X2=0.82
+ $Y2=1.46
cc_101 N_VNB_M1029_b N_A_2624_107#_c_1718_n 0.0549768f $X=-0.33 $Y=-0.265
+ $X2=0.82 $Y2=1.46
cc_102 N_VNB_M1029_b N_A_2624_107#_c_1719_n 0.137362f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_103 N_VNB_M1029_b N_A_2624_107#_M1009_g 0.0594077f $X=-0.33 $Y=-0.265
+ $X2=3.485 $Y2=1.36
cc_104 N_VNB_c_3_p N_A_2624_107#_M1009_g 7.93986e-19 $X=0.24 $Y=0 $X2=3.485
+ $Y2=1.36
cc_105 N_VNB_M1029_b N_A_2624_107#_c_1722_n 0.0363285f $X=-0.33 $Y=-0.265
+ $X2=1.765 $Y2=2.75
cc_106 N_VNB_M1029_b N_A_2624_107#_c_1723_n 0.00311731f $X=-0.33 $Y=-0.265
+ $X2=2.875 $Y2=2.75
cc_107 N_VNB_M1029_b N_A_2624_107#_c_1724_n 0.00162824f $X=-0.33 $Y=-0.265
+ $X2=2.875 $Y2=2.75
cc_108 N_VNB_M1029_b N_A_2624_107#_c_1725_n 8.96666e-19 $X=-0.33 $Y=-0.265
+ $X2=0.82 $Y2=1.295
cc_109 N_VNB_M1029_b N_A_2624_107#_c_1726_n 0.0022812f $X=-0.33 $Y=-0.265
+ $X2=0.86 $Y2=0.865
cc_110 N_VNB_M1029_b N_A_2624_107#_c_1727_n 0.0144999f $X=-0.33 $Y=-0.265
+ $X2=0.86 $Y2=0.865
cc_111 N_VNB_M1029_b N_A_3613_443#_M1010_g 0.0478348f $X=-0.33 $Y=-0.265
+ $X2=3.83 $Y2=0.745
cc_112 N_VNB_c_3_p N_A_3613_443#_M1010_g 8.51801e-19 $X=0.24 $Y=0 $X2=3.83
+ $Y2=0.745
cc_113 N_VNB_M1029_b N_A_3613_443#_c_1879_n 0.0158683f $X=-0.33 $Y=-0.265
+ $X2=0.86 $Y2=2.865
cc_114 N_VNB_M1029_b N_A_3613_443#_c_1880_n 0.00293136f $X=-0.33 $Y=-0.265
+ $X2=1.515 $Y2=0.35
cc_115 N_VNB_M1029_b N_A_3613_443#_c_1881_n 0.0329714f $X=-0.33 $Y=-0.265
+ $X2=0.985 $Y2=0.35
cc_116 N_VNB_M1029_b N_A_339_655#_c_2080_n 0.00820675f $X=-0.33 $Y=-0.265
+ $X2=0.82 $Y2=1.46
cc_117 N_VNB_M1029_b N_A_339_655#_c_2081_n 0.0149651f $X=-0.33 $Y=-0.265
+ $X2=1.515 $Y2=0.35
cc_118 N_VNB_M1029_b N_A_339_655#_c_2082_n 0.00372437f $X=-0.33 $Y=-0.265
+ $X2=2.875 $Y2=2.75
cc_119 N_VNB_M1029_b N_A_339_655#_c_2083_n 0.00202928f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_120 N_VNB_M1029_b N_A_339_655#_c_2084_n 0.00522997f $X=-0.33 $Y=-0.265
+ $X2=3.515 $Y2=1.58
cc_121 N_VNB_M1029_b N_A_339_655#_c_2085_n 0.00206288f $X=-0.33 $Y=-0.265
+ $X2=0.86 $Y2=0.865
cc_122 N_VNB_M1029_b N_A_339_655#_c_2086_n 0.0048957f $X=-0.33 $Y=-0.265
+ $X2=3.83 $Y2=1.507
cc_123 N_VNB_M1029_b N_Q_N_c_2263_n 0.0211237f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_124 N_VNB_c_3_p N_Q_N_c_2263_n 0.00110923f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_125 N_VNB_M1029_b Q 0.0562342f $X=-0.33 $Y=-0.265 $X2=2.94 $Y2=3.485
cc_126 N_VNB_M1029_b N_VGND_c_2294_n 0.0785992f $X=-0.33 $Y=-0.265 $X2=1.515
+ $Y2=0.35
cc_127 N_VNB_c_3_p N_VGND_c_2294_n 0.00154107f $X=0.24 $Y=0 $X2=1.515 $Y2=0.35
cc_128 N_VNB_M1029_b N_VGND_c_2296_n 0.0435124f $X=-0.33 $Y=-0.265 $X2=2.875
+ $Y2=2.75
cc_129 N_VNB_c_3_p N_VGND_c_2296_n 0.00342965f $X=0.24 $Y=0 $X2=2.875 $Y2=2.75
cc_130 N_VNB_M1029_b N_VGND_c_2298_n 0.0532326f $X=-0.33 $Y=-0.265 $X2=1.6
+ $Y2=2.83
cc_131 N_VNB_c_3_p N_VGND_c_2298_n 0.00241477f $X=0.24 $Y=0 $X2=1.6 $Y2=2.83
cc_132 N_VNB_M1029_b N_VGND_c_2300_n 0.0503771f $X=-0.33 $Y=-0.265 $X2=3.385
+ $Y2=2.685
cc_133 N_VNB_c_3_p N_VGND_c_2300_n 0.00377509f $X=0.24 $Y=0 $X2=3.385 $Y2=2.685
cc_134 N_VNB_M1029_b N_VGND_c_2302_n 0.0464657f $X=-0.33 $Y=-0.265 $X2=3.765
+ $Y2=1.507
cc_135 N_VNB_c_3_p N_VGND_c_2302_n 0.00270113f $X=0.24 $Y=0 $X2=3.765 $Y2=1.507
cc_136 N_VNB_M1029_b N_VGND_c_2304_n 0.0415113f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_137 N_VNB_c_3_p N_VGND_c_2304_n 0.0014985f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_138 N_VNB_M1029_b N_VGND_c_2306_n 0.0560138f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_139 N_VNB_c_3_p N_VGND_c_2306_n 0.00269049f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_140 N_VNB_M1029_b N_VGND_c_2308_n 0.238014f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_141 N_VNB_c_3_p N_VGND_c_2308_n 2.1442f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_142 N_VNB_M1029_b N_noxref_25_c_2431_n 0.00322716f $X=-0.33 $Y=-0.265
+ $X2=3.385 $Y2=1.89
cc_143 N_VNB_M1029_b N_noxref_25_c_2432_n 0.189113f $X=-0.33 $Y=-0.265 $X2=3.83
+ $Y2=1.125
cc_144 N_VNB_c_3_p N_noxref_25_c_2432_n 0.00895182f $X=0.24 $Y=0 $X2=3.83
+ $Y2=1.125
cc_145 N_VNB_M1029_b N_noxref_25_c_2434_n 0.0187012f $X=-0.33 $Y=-0.265 $X2=3.83
+ $Y2=0.745
cc_146 N_VNB_c_3_p N_noxref_25_c_2434_n 8.29076e-19 $X=0.24 $Y=0 $X2=3.83
+ $Y2=0.745
cc_147 N_VNB_M1029_b N_noxref_25_c_2436_n 0.0263861f $X=-0.33 $Y=-0.265 $X2=3.83
+ $Y2=0.745
cc_148 N_VNB_c_3_p N_noxref_25_c_2436_n 0.00109273f $X=0.24 $Y=0 $X2=3.83
+ $Y2=0.745
cc_149 N_VPB_M1018_b N_SCE_M1018_g 0.0482163f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=3.455
cc_150 VPB N_SCE_M1018_g 0.00274588f $X=0 $Y=3.955 $X2=0.86 $Y2=3.455
cc_151 N_VPB_c_151_p N_SCE_M1018_g 0.0104959f $X=19.92 $Y=4.07 $X2=0.86
+ $Y2=3.455
cc_152 N_VPB_M1018_b N_SCE_M1016_g 0.0644694f $X=-0.33 $Y=1.885 $X2=2.94
+ $Y2=3.485
cc_153 VPB N_SCE_M1016_g 0.00957431f $X=0 $Y=3.955 $X2=2.94 $Y2=3.485
cc_154 N_VPB_c_151_p N_SCE_M1016_g 0.0134742f $X=19.92 $Y=4.07 $X2=2.94
+ $Y2=3.485
cc_155 N_VPB_M1018_b N_SCE_c_378_n 0.0470954f $X=-0.33 $Y=1.885 $X2=3.385
+ $Y2=2.565
cc_156 N_VPB_M1018_b N_SCE_c_379_n 0.0541681f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=2.865
cc_157 N_VPB_M1018_b N_SCE_c_380_n 0.00824168f $X=-0.33 $Y=1.885 $X2=2.875
+ $Y2=2.75
cc_158 N_VPB_M1018_b N_SCE_c_381_n 0.0820548f $X=-0.33 $Y=1.885 $X2=1.6 $Y2=2.83
cc_159 N_VPB_M1018_b N_SCE_M1029_g 0.0950419f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=0.865
cc_160 N_VPB_M1018_b N_SCE_c_383_n 0.0469985f $X=-0.33 $Y=1.885 $X2=3.385
+ $Y2=2.685
cc_161 N_VPB_M1018_b N_SCE_c_370_n 0.0188907f $X=-0.33 $Y=1.885 $X2=3.765
+ $Y2=1.365
cc_162 N_VPB_M1018_b N_D_M1001_g 0.160269f $X=-0.33 $Y=1.885 $X2=0.86 $Y2=3.455
cc_163 VPB N_D_M1001_g 0.00957431f $X=0 $Y=3.955 $X2=0.86 $Y2=3.455
cc_164 N_VPB_c_151_p N_D_M1001_g 0.0176223f $X=19.92 $Y=4.07 $X2=0.86 $Y2=3.455
cc_165 N_VPB_M1018_b N_D_c_487_n 0.00763964f $X=-0.33 $Y=1.885 $X2=3.83
+ $Y2=0.745
cc_166 N_VPB_M1018_b N_A_222_131#_c_529_n 0.0266558f $X=-0.33 $Y=1.885 $X2=3.83
+ $Y2=0.745
cc_167 N_VPB_M1018_b N_A_222_131#_M1006_g 0.0438179f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=2.615
cc_168 VPB N_A_222_131#_M1006_g 0.00957431f $X=0 $Y=3.955 $X2=0.86 $Y2=2.615
cc_169 N_VPB_c_151_p N_A_222_131#_M1006_g 0.0188852f $X=19.92 $Y=4.07 $X2=0.86
+ $Y2=2.615
cc_170 N_VPB_M1018_b N_A_222_131#_c_526_n 0.0110198f $X=-0.33 $Y=1.885 $X2=0.9
+ $Y2=1.295
cc_171 N_VPB_M1018_b N_A_222_131#_c_534_n 0.00224254f $X=-0.33 $Y=1.885 $X2=1.6
+ $Y2=1.275
cc_172 N_VPB_M1018_b N_A_222_131#_c_535_n 0.00429695f $X=-0.33 $Y=1.885
+ $X2=1.685 $Y2=1.36
cc_173 VPB N_A_222_131#_c_535_n 7.04937e-19 $X=0 $Y=3.955 $X2=1.685 $Y2=1.36
cc_174 N_VPB_c_151_p N_A_222_131#_c_535_n 0.0107078f $X=19.92 $Y=4.07 $X2=1.685
+ $Y2=1.36
cc_175 N_VPB_M1018_b N_A_222_131#_c_538_n 0.0302366f $X=-0.33 $Y=1.885 $X2=2.875
+ $Y2=2.75
cc_176 N_VPB_M1018_b N_A_222_131#_c_528_n 0.0340948f $X=-0.33 $Y=1.885 $X2=1.64
+ $Y2=2.75
cc_177 N_VPB_M1018_b N_A_222_131#_c_540_n 0.00896362f $X=-0.33 $Y=1.885 $X2=1.64
+ $Y2=2.83
cc_178 N_VPB_M1018_b N_A_222_131#_c_541_n 0.0167101f $X=-0.33 $Y=1.885 $X2=3.515
+ $Y2=1.58
cc_179 N_VPB_M1018_b N_A_222_131#_c_542_n 0.00173311f $X=-0.33 $Y=1.885
+ $X2=3.995 $Y2=1.58
cc_180 N_VPB_M1018_b N_A_222_131#_c_543_n 0.0465796f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=0.865
cc_181 N_VPB_M1018_b N_A_222_131#_c_544_n 0.00258443f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=1.46
cc_182 N_VPB_M1018_b N_A_222_131#_c_545_n 0.00496696f $X=-0.33 $Y=1.885 $X2=1.6
+ $Y2=2.865
cc_183 N_VPB_M1018_b N_A_222_131#_c_546_n 0.00205601f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_184 N_VPB_M1018_b N_SCD_c_659_n 0.0502154f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=3.115
cc_185 VPB N_SCD_c_659_n 0.00957431f $X=0 $Y=3.955 $X2=0.86 $Y2=3.115
cc_186 N_VPB_c_151_p N_SCD_c_659_n 0.0188741f $X=19.92 $Y=4.07 $X2=0.86
+ $Y2=3.115
cc_187 N_VPB_M1018_b N_SCD_c_662_n 0.0289753f $X=-0.33 $Y=1.885 $X2=2.94
+ $Y2=3.485
cc_188 N_VPB_M1018_b N_SCD_c_663_n 0.00909535f $X=-0.33 $Y=1.885 $X2=2.94
+ $Y2=3.485
cc_189 N_VPB_M1018_b N_SCD_c_664_n 0.00398331f $X=-0.33 $Y=1.885 $X2=3.385
+ $Y2=1.89
cc_190 N_VPB_M1018_b N_SCD_c_665_n 0.0395386f $X=-0.33 $Y=1.885 $X2=3.83
+ $Y2=0.745
cc_191 N_VPB_M1018_b N_SCD_M1035_g 0.0233766f $X=-0.33 $Y=1.885 $X2=0.82
+ $Y2=1.46
cc_192 N_VPB_M1018_b N_SCD_c_667_n 0.00397201f $X=-0.33 $Y=1.885 $X2=1.685
+ $Y2=1.36
cc_193 N_VPB_M1018_b N_CLK_M1002_g 0.0699386f $X=-0.33 $Y=1.885 $X2=2.94
+ $Y2=3.485
cc_194 VPB N_CLK_M1002_g 0.00970178f $X=0 $Y=3.955 $X2=2.94 $Y2=3.485
cc_195 N_VPB_c_151_p N_CLK_M1002_g 0.0157135f $X=19.92 $Y=4.07 $X2=2.94
+ $Y2=3.485
cc_196 N_VPB_M1018_b N_CLK_c_726_n 0.0741291f $X=-0.33 $Y=1.885 $X2=3.83
+ $Y2=0.745
cc_197 N_VPB_M1018_b N_A_1569_126#_c_781_n 0.158573f $X=-0.33 $Y=1.885 $X2=2.94
+ $Y2=3.485
cc_198 VPB N_A_1569_126#_c_781_n 0.00970178f $X=0 $Y=3.955 $X2=2.94 $Y2=3.485
cc_199 N_VPB_c_151_p N_A_1569_126#_c_781_n 0.0161942f $X=19.92 $Y=4.07 $X2=2.94
+ $Y2=3.485
cc_200 N_VPB_M1018_b N_A_1569_126#_c_761_n 0.00501221f $X=-0.33 $Y=1.885
+ $X2=0.82 $Y2=1.46
cc_201 N_VPB_M1018_b N_A_1569_126#_c_774_n 0.00425379f $X=-0.33 $Y=1.885 $X2=1.6
+ $Y2=2.83
cc_202 N_VPB_M1018_b N_A_1569_126#_c_786_n 0.0872477f $X=-0.33 $Y=1.885 $X2=1.6
+ $Y2=2.83
cc_203 N_VPB_M1018_b N_A_1569_126#_c_787_n 0.00677117f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_204 N_VPB_M1018_b N_A_1290_126#_M1019_g 0.0677537f $X=-0.33 $Y=1.885 $X2=3.83
+ $Y2=0.745
cc_205 N_VPB_M1018_b N_A_1290_126#_c_950_n 0.00954664f $X=-0.33 $Y=1.885
+ $X2=0.82 $Y2=1.46
cc_206 N_VPB_M1018_b N_A_1290_126#_M1037_g 0.095731f $X=-0.33 $Y=1.885 $X2=0.9
+ $Y2=0.435
cc_207 VPB N_A_1290_126#_M1037_g 0.00970178f $X=0 $Y=3.955 $X2=0.9 $Y2=0.435
cc_208 N_VPB_c_151_p N_A_1290_126#_M1037_g 0.0193887f $X=19.92 $Y=4.07 $X2=0.9
+ $Y2=0.435
cc_209 N_VPB_M1018_b N_A_1290_126#_M1024_g 0.0373671f $X=-0.33 $Y=1.885 $X2=1.6
+ $Y2=0.435
cc_210 VPB N_A_1290_126#_M1024_g 0.00970178f $X=0 $Y=3.955 $X2=1.6 $Y2=0.435
cc_211 N_VPB_c_151_p N_A_1290_126#_M1024_g 0.0191024f $X=19.92 $Y=4.07 $X2=1.6
+ $Y2=0.435
cc_212 N_VPB_M1018_b N_A_1290_126#_c_957_n 0.0243125f $X=-0.33 $Y=1.885
+ $X2=3.515 $Y2=1.58
cc_213 N_VPB_M1018_b N_A_1290_126#_c_974_n 0.015459f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=0.865
cc_214 N_VPB_M1018_b N_A_1290_126#_c_975_n 0.00439753f $X=-0.33 $Y=1.885
+ $X2=0.86 $Y2=1.46
cc_215 N_VPB_M1018_b N_A_1290_126#_c_959_n 0.00220421f $X=-0.33 $Y=1.885 $X2=1.6
+ $Y2=2.865
cc_216 N_VPB_M1018_b N_A_1290_126#_c_960_n 0.00174719f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_217 N_VPB_M1018_b N_A_1290_126#_c_978_n 0.00446596f $X=-0.33 $Y=1.885
+ $X2=3.385 $Y2=2.685
cc_218 N_VPB_M1018_b N_A_1290_126#_c_979_n 0.0944008f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_219 N_VPB_M1018_b N_A_1290_126#_c_964_n 0.106126f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_220 N_VPB_M1018_b N_A_2014_537#_c_1170_n 0.0595339f $X=-0.33 $Y=1.885
+ $X2=3.83 $Y2=0.745
cc_221 N_VPB_M1018_b N_A_2014_537#_c_1171_n 0.0826595f $X=-0.33 $Y=1.885
+ $X2=3.83 $Y2=0.745
cc_222 VPB N_A_2014_537#_c_1171_n 0.00970178f $X=0 $Y=3.955 $X2=3.83 $Y2=0.745
cc_223 N_VPB_c_151_p N_A_2014_537#_c_1171_n 0.013715f $X=19.92 $Y=4.07 $X2=3.83
+ $Y2=0.745
cc_224 N_VPB_M1018_b N_A_2014_537#_c_1163_n 0.0113858f $X=-0.33 $Y=1.885
+ $X2=0.86 $Y2=2.615
cc_225 N_VPB_M1018_b N_A_2014_537#_c_1166_n 0.0051335f $X=-0.33 $Y=1.885
+ $X2=0.985 $Y2=0.35
cc_226 N_VPB_M1018_b N_A_2014_537#_c_1167_n 0.00140118f $X=-0.33 $Y=1.885
+ $X2=1.6 $Y2=0.435
cc_227 N_VPB_M1018_b N_A_2014_537#_c_1177_n 0.00156545f $X=-0.33 $Y=1.885
+ $X2=1.685 $Y2=1.36
cc_228 VPB N_A_2014_537#_c_1177_n 8.01732e-19 $X=0 $Y=3.955 $X2=1.685 $Y2=1.36
cc_229 N_VPB_c_151_p N_A_2014_537#_c_1177_n 0.0130099f $X=19.92 $Y=4.07
+ $X2=1.685 $Y2=1.36
cc_230 N_VPB_M1018_b N_A_2014_537#_c_1180_n 0.00178063f $X=-0.33 $Y=1.885
+ $X2=2.875 $Y2=2.75
cc_231 N_VPB_M1018_b N_A_2014_537#_c_1181_n 0.00317366f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_232 N_VPB_M1018_b N_RESET_B_M1013_g 0.0393042f $X=-0.33 $Y=1.885 $X2=3.83
+ $Y2=0.745
cc_233 VPB N_RESET_B_M1013_g 0.00970178f $X=0 $Y=3.955 $X2=3.83 $Y2=0.745
cc_234 N_VPB_c_151_p N_RESET_B_M1013_g 0.0190953f $X=19.92 $Y=4.07 $X2=3.83
+ $Y2=0.745
cc_235 N_VPB_M1018_b N_RESET_B_c_1301_n 0.0364991f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_236 N_VPB_M1018_b N_RESET_B_c_1302_n 0.0889846f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_237 VPB N_RESET_B_c_1302_n 0.00957431f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_238 N_VPB_c_151_p N_RESET_B_c_1302_n 0.0143649f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_239 N_VPB_M1018_b N_RESET_B_c_1305_n 0.0551429f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_240 N_VPB_M1018_b N_RESET_B_c_1289_n 0.0770446f $X=-0.33 $Y=1.885 $X2=1.515
+ $Y2=0.35
cc_241 N_VPB_M1018_b RESET_B 0.00425288f $X=-0.33 $Y=1.885 $X2=1.6 $Y2=1.275
cc_242 N_VPB_M1018_b N_RESET_B_c_1308_n 0.073365f $X=-0.33 $Y=1.885 $X2=1.765
+ $Y2=2.75
cc_243 N_VPB_M1018_b N_RESET_B_c_1309_n 0.00414252f $X=-0.33 $Y=1.885 $X2=2.875
+ $Y2=2.75
cc_244 N_VPB_M1018_b N_RESET_B_c_1310_n 0.0307562f $X=-0.33 $Y=1.885 $X2=2.875
+ $Y2=2.75
cc_245 N_VPB_M1018_b N_RESET_B_c_1311_n 0.00252623f $X=-0.33 $Y=1.885 $X2=2.875
+ $Y2=2.75
cc_246 N_VPB_M1018_b N_RESET_B_c_1312_n 0.00389375f $X=-0.33 $Y=1.885 $X2=3.515
+ $Y2=1.58
cc_247 N_VPB_M1018_b N_RESET_B_c_1291_n 0.074179f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=0.865
cc_248 N_VPB_M1018_b N_RESET_B_M1008_g 0.0682592f $X=-0.33 $Y=1.885 $X2=1.6
+ $Y2=2.865
cc_249 N_VPB_M1018_b N_RESET_B_c_1293_n 0.00301579f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_250 N_VPB_M1018_b N_RESET_B_c_1297_n 0.00192363f $X=-0.33 $Y=1.885 $X2=3.485
+ $Y2=1.535
cc_251 N_VPB_M1018_b N_A_1816_659#_M1039_g 0.0191722f $X=-0.33 $Y=1.885 $X2=3.83
+ $Y2=0.745
cc_252 N_VPB_M1018_b N_A_1816_659#_M1003_g 0.0393182f $X=-0.33 $Y=1.885 $X2=1.11
+ $Y2=2.865
cc_253 VPB N_A_1816_659#_M1003_g 0.00970178f $X=0 $Y=3.955 $X2=1.11 $Y2=2.865
cc_254 N_VPB_c_151_p N_A_1816_659#_M1003_g 0.0154024f $X=19.92 $Y=4.07 $X2=1.11
+ $Y2=2.865
cc_255 N_VPB_M1018_b N_A_1816_659#_c_1500_n 0.00968768f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_256 N_VPB_M1018_b N_A_1816_659#_c_1507_n 0.0030332f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_257 VPB N_A_1816_659#_c_1507_n 8.01732e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_258 N_VPB_c_151_p N_A_1816_659#_c_1507_n 0.0130099f $X=19.92 $Y=4.07 $X2=0
+ $Y2=0
cc_259 N_VPB_M1018_b N_A_1816_659#_c_1510_n 0.00943946f $X=-0.33 $Y=1.885
+ $X2=0.9 $Y2=1.295
cc_260 N_VPB_M1018_b N_A_1816_659#_c_1511_n 0.0124034f $X=-0.33 $Y=1.885
+ $X2=0.985 $Y2=0.35
cc_261 N_VPB_M1018_b N_A_1816_659#_c_1512_n 0.00978305f $X=-0.33 $Y=1.885
+ $X2=1.6 $Y2=1.275
cc_262 VPB N_A_1816_659#_c_1512_n 0.00137465f $X=0 $Y=3.955 $X2=1.6 $Y2=1.275
cc_263 N_VPB_c_151_p N_A_1816_659#_c_1512_n 0.0216688f $X=19.92 $Y=4.07 $X2=1.6
+ $Y2=1.275
cc_264 N_VPB_M1018_b N_A_1816_659#_c_1515_n 0.00168656f $X=-0.33 $Y=1.885
+ $X2=2.875 $Y2=2.75
cc_265 N_VPB_M1018_b N_A_1816_659#_c_1516_n 0.00208646f $X=-0.33 $Y=1.885
+ $X2=1.6 $Y2=2.83
cc_266 N_VPB_M1018_b N_A_1816_659#_c_1517_n 0.10089f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_267 N_VPB_M1018_b N_A_2841_81#_c_1625_n 0.00566963f $X=-0.33 $Y=1.885
+ $X2=0.86 $Y2=2.865
cc_268 N_VPB_M1018_b N_A_2841_81#_c_1626_n 0.0438305f $X=-0.33 $Y=1.885 $X2=0.82
+ $Y2=1.46
cc_269 N_VPB_M1018_b N_A_2841_81#_c_1627_n 0.00555045f $X=-0.33 $Y=1.885 $X2=0.9
+ $Y2=1.295
cc_270 N_VPB_M1018_b N_A_2841_81#_c_1628_n 0.00264205f $X=-0.33 $Y=1.885 $X2=1.6
+ $Y2=0.435
cc_271 N_VPB_M1018_b N_A_2841_81#_c_1629_n 9.66992e-19 $X=-0.33 $Y=1.885
+ $X2=3.485 $Y2=1.36
cc_272 N_VPB_M1018_b N_A_2841_81#_c_1630_n 9.27498e-19 $X=-0.33 $Y=1.885
+ $X2=2.875 $Y2=2.75
cc_273 N_VPB_M1018_b N_A_2841_81#_c_1624_n 0.023567f $X=-0.33 $Y=1.885 $X2=1.64
+ $Y2=2.83
cc_274 N_VPB_M1018_b N_A_2841_81#_c_1632_n 0.036297f $X=-0.33 $Y=1.885 $X2=1.6
+ $Y2=2.83
cc_275 N_VPB_M1018_b N_A_2624_107#_M1021_g 0.0966071f $X=-0.33 $Y=1.885 $X2=3.83
+ $Y2=0.745
cc_276 N_VPB_M1018_b N_A_2624_107#_M1032_g 0.0436592f $X=-0.33 $Y=1.885 $X2=1.11
+ $Y2=2.865
cc_277 VPB N_A_2624_107#_M1032_g 0.00116559f $X=0 $Y=3.955 $X2=1.11 $Y2=2.865
cc_278 N_VPB_c_151_p N_A_2624_107#_M1032_g 0.00661471f $X=19.92 $Y=4.07 $X2=1.11
+ $Y2=2.865
cc_279 N_VPB_M1018_b N_A_2624_107#_c_1718_n 0.0361702f $X=-0.33 $Y=1.885
+ $X2=0.82 $Y2=1.46
cc_280 N_VPB_M1018_b N_A_2624_107#_c_1719_n 0.0421483f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_281 N_VPB_M1018_b N_A_2624_107#_M1036_g 0.0431139f $X=-0.33 $Y=1.885
+ $X2=1.515 $Y2=0.35
cc_282 N_VPB_M1018_b N_A_2624_107#_c_1722_n 0.0202503f $X=-0.33 $Y=1.885
+ $X2=1.765 $Y2=2.75
cc_283 N_VPB_M1018_b N_A_2624_107#_c_1736_n 0.0138797f $X=-0.33 $Y=1.885 $X2=1.6
+ $Y2=2.83
cc_284 VPB N_A_2624_107#_c_1736_n 0.00104693f $X=0 $Y=3.955 $X2=1.6 $Y2=2.83
cc_285 N_VPB_c_151_p N_A_2624_107#_c_1736_n 0.0172373f $X=19.92 $Y=4.07 $X2=1.6
+ $Y2=2.83
cc_286 N_VPB_M1018_b N_A_2624_107#_c_1739_n 0.00539052f $X=-0.33 $Y=1.885
+ $X2=3.515 $Y2=1.58
cc_287 N_VPB_M1018_b N_A_2624_107#_c_1726_n 0.00532175f $X=-0.33 $Y=1.885
+ $X2=0.86 $Y2=0.865
cc_288 N_VPB_M1018_b N_A_3613_443#_M1022_g 0.0425385f $X=-0.33 $Y=1.885
+ $X2=3.385 $Y2=1.89
cc_289 VPB N_A_3613_443#_M1022_g 0.00970178f $X=0 $Y=3.955 $X2=3.385 $Y2=1.89
cc_290 N_VPB_c_151_p N_A_3613_443#_M1022_g 0.0162989f $X=19.92 $Y=4.07 $X2=3.385
+ $Y2=1.89
cc_291 N_VPB_M1018_b N_A_3613_443#_c_1885_n 0.0147452f $X=-0.33 $Y=1.885
+ $X2=0.82 $Y2=1.46
cc_292 N_VPB_M1018_b N_A_3613_443#_c_1880_n 0.00298737f $X=-0.33 $Y=1.885
+ $X2=1.515 $Y2=0.35
cc_293 N_VPB_M1018_b N_A_3613_443#_c_1881_n 0.0228896f $X=-0.33 $Y=1.885
+ $X2=0.985 $Y2=0.35
cc_294 N_VPB_M1018_b N_A_3613_443#_c_1888_n 4.99077e-19 $X=-0.33 $Y=1.885
+ $X2=1.6 $Y2=1.275
cc_295 N_VPB_M1018_b N_VPWR_c_1922_n 0.040862f $X=-0.33 $Y=1.885 $X2=1.765
+ $Y2=2.75
cc_296 VPB N_VPWR_c_1922_n 0.00320333f $X=0 $Y=3.955 $X2=1.765 $Y2=2.75
cc_297 N_VPB_c_151_p N_VPWR_c_1922_n 0.0369986f $X=19.92 $Y=4.07 $X2=1.765
+ $Y2=2.75
cc_298 N_VPB_M1018_b N_VPWR_c_1925_n 0.00231721f $X=-0.33 $Y=1.885 $X2=3.995
+ $Y2=1.58
cc_299 VPB N_VPWR_c_1925_n 0.00365012f $X=0 $Y=3.955 $X2=3.995 $Y2=1.58
cc_300 N_VPB_c_151_p N_VPWR_c_1925_n 0.0436237f $X=19.92 $Y=4.07 $X2=3.995
+ $Y2=1.58
cc_301 N_VPB_M1018_b N_VPWR_c_1928_n 0.00214168f $X=-0.33 $Y=1.885 $X2=2.875
+ $Y2=2.685
cc_302 VPB N_VPWR_c_1928_n 0.00340168f $X=0 $Y=3.955 $X2=2.875 $Y2=2.685
cc_303 N_VPB_c_151_p N_VPWR_c_1928_n 0.0448224f $X=19.92 $Y=4.07 $X2=2.875
+ $Y2=2.685
cc_304 N_VPB_M1018_b N_VPWR_c_1931_n 0.0200833f $X=-0.33 $Y=1.885 $X2=3.765
+ $Y2=1.507
cc_305 VPB N_VPWR_c_1931_n 4.76796e-19 $X=0 $Y=3.955 $X2=3.765 $Y2=1.507
cc_306 N_VPB_c_151_p N_VPWR_c_1931_n 0.00726526f $X=19.92 $Y=4.07 $X2=3.765
+ $Y2=1.507
cc_307 N_VPB_M1018_b N_VPWR_c_1934_n 0.00638817f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_1934_n 0.00375873f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_309 N_VPB_c_151_p N_VPWR_c_1934_n 0.0477601f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_310 N_VPB_M1018_b N_VPWR_c_1937_n 0.00117792f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_1937_n 0.00241469f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_312 N_VPB_c_151_p N_VPWR_c_1937_n 0.0271364f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_313 N_VPB_M1018_b N_VPWR_c_1940_n 0.0312271f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_1940_n 0.00260535f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_315 N_VPB_c_151_p N_VPWR_c_1940_n 0.0396995f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_316 N_VPB_M1018_b N_VPWR_c_1943_n 0.0183294f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_317 VPB N_VPWR_c_1943_n 0.00261954f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_318 N_VPB_c_151_p N_VPWR_c_1943_n 0.0399157f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_319 N_VPB_M1018_b N_VPWR_c_1946_n 0.0322743f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_320 VPB N_VPWR_c_1946_n 0.00335473f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_321 N_VPB_c_151_p N_VPWR_c_1946_n 0.0490696f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_322 N_VPB_M1018_b N_VPWR_c_1949_n 0.172006f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_323 VPB N_VPWR_c_1949_n 2.14549f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_324 N_VPB_c_151_p N_VPWR_c_1949_n 0.103238f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_325 N_VPB_M1018_b N_A_339_655#_c_2087_n 0.0124523f $X=-0.33 $Y=1.885 $X2=1.11
+ $Y2=2.865
cc_326 N_VPB_M1018_b N_A_339_655#_c_2088_n 0.0118364f $X=-0.33 $Y=1.885 $X2=0.86
+ $Y2=2.865
cc_327 VPB N_A_339_655#_c_2088_n 0.0015589f $X=0 $Y=3.955 $X2=0.86 $Y2=2.865
cc_328 N_VPB_c_151_p N_A_339_655#_c_2088_n 0.0207778f $X=19.92 $Y=4.07 $X2=0.86
+ $Y2=2.865
cc_329 N_VPB_M1018_b N_A_339_655#_c_2091_n 0.00213583f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_330 VPB N_A_339_655#_c_2091_n 7.80441e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_331 N_VPB_c_151_p N_A_339_655#_c_2091_n 0.0119623f $X=19.92 $Y=4.07 $X2=0
+ $Y2=0
cc_332 N_VPB_M1018_b N_A_339_655#_c_2081_n 0.0208764f $X=-0.33 $Y=1.885
+ $X2=1.515 $Y2=0.35
cc_333 N_VPB_M1018_b N_A_339_655#_c_2095_n 0.00405521f $X=-0.33 $Y=1.885
+ $X2=0.985 $Y2=0.35
cc_334 N_VPB_M1018_b N_A_339_655#_c_2096_n 0.00728213f $X=-0.33 $Y=1.885
+ $X2=1.685 $Y2=1.36
cc_335 VPB N_A_339_655#_c_2096_n 0.00248257f $X=0 $Y=3.955 $X2=1.685 $Y2=1.36
cc_336 N_VPB_c_151_p N_A_339_655#_c_2096_n 0.0459346f $X=19.92 $Y=4.07 $X2=1.685
+ $Y2=1.36
cc_337 VPB N_A_339_655#_c_2099_n 8.21022e-19 $X=0 $Y=3.955 $X2=1.765 $Y2=2.75
cc_338 N_VPB_c_151_p N_A_339_655#_c_2099_n 0.0108189f $X=19.92 $Y=4.07 $X2=1.765
+ $Y2=2.75
cc_339 N_VPB_M1018_b N_A_339_655#_c_2101_n 0.0326832f $X=-0.33 $Y=1.885
+ $X2=2.875 $Y2=2.75
cc_340 N_VPB_M1018_b N_A_339_655#_c_2082_n 0.00477457f $X=-0.33 $Y=1.885
+ $X2=2.875 $Y2=2.75
cc_341 N_VPB_M1018_b N_A_339_655#_c_2083_n 0.00166376f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_342 N_VPB_M1018_b N_A_339_655#_c_2104_n 0.00437969f $X=-0.33 $Y=1.885
+ $X2=1.64 $Y2=2.75
cc_343 N_VPB_M1018_b N_A_339_655#_c_2105_n 0.0147851f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_344 N_VPB_c_151_p N_A_339_655#_c_2105_n 0.0078046f $X=19.92 $Y=4.07 $X2=0
+ $Y2=0
cc_345 N_VPB_M1018_b N_A_339_655#_c_2107_n 0.00426083f $X=-0.33 $Y=1.885
+ $X2=1.64 $Y2=2.83
cc_346 N_VPB_c_151_p N_A_339_655#_c_2107_n 0.00266145f $X=19.92 $Y=4.07 $X2=1.64
+ $Y2=2.83
cc_347 N_VPB_c_151_p N_A_339_655#_c_2109_n 0.00466818f $X=19.92 $Y=4.07 $X2=1.6
+ $Y2=2.83
cc_348 N_VPB_M1018_b N_A_339_655#_c_2084_n 0.00929154f $X=-0.33 $Y=1.885
+ $X2=3.515 $Y2=1.58
cc_349 N_VPB_M1018_b N_A_339_655#_c_2111_n 0.00977095f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_350 N_VPB_M1018_b N_A_339_655#_c_2112_n 0.00913981f $X=-0.33 $Y=1.885
+ $X2=2.875 $Y2=2.685
cc_351 VPB N_A_339_655#_c_2112_n 0.0010482f $X=0 $Y=3.955 $X2=2.875 $Y2=2.685
cc_352 N_VPB_c_151_p N_A_339_655#_c_2112_n 0.017156f $X=19.92 $Y=4.07 $X2=2.875
+ $Y2=2.685
cc_353 N_VPB_M1018_b N_Q_N_c_2263_n 0.030692f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_354 VPB N_Q_N_c_2263_n 0.00106329f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_355 N_VPB_c_151_p N_Q_N_c_2263_n 0.0107605f $X=19.92 $Y=4.07 $X2=0 $Y2=0
cc_356 N_VPB_M1018_b Q 0.0670661f $X=-0.33 $Y=1.885 $X2=2.94 $Y2=3.485
cc_357 VPB Q 0.00107758f $X=0 $Y=3.955 $X2=2.94 $Y2=3.485
cc_358 N_VPB_c_151_p Q 0.0177658f $X=19.92 $Y=4.07 $X2=2.94 $Y2=3.485
cc_359 N_SCE_c_371_n N_D_c_484_n 0.049474f $X=3.485 $Y=1.535 $X2=0 $Y2=0
cc_360 N_SCE_c_380_n N_D_M1001_g 0.0250491f $X=2.875 $Y=2.75 $X2=0 $Y2=0
cc_361 N_SCE_c_387_p N_D_M1001_g 0.00128763f $X=1.64 $Y=2.75 $X2=0 $Y2=0
cc_362 N_SCE_c_381_n N_D_M1001_g 0.0351805f $X=1.6 $Y=2.83 $X2=0 $Y2=0
cc_363 N_SCE_c_383_n N_D_M1001_g 0.0897974f $X=3.385 $Y=2.685 $X2=0 $Y2=0
cc_364 N_SCE_c_364_n N_D_M1040_g 0.00981955f $X=1.6 $Y=1.275 $X2=0 $Y2=0
cc_365 N_SCE_c_365_n N_D_c_487_n 0.0105212f $X=1.685 $Y=1.36 $X2=0 $Y2=0
cc_366 N_SCE_c_371_n N_D_c_487_n 0.0483839f $X=3.485 $Y=1.535 $X2=0 $Y2=0
cc_367 N_SCE_M1031_g N_A_222_131#_M1041_g 0.0166023f $X=3.83 $Y=0.745 $X2=0
+ $Y2=0
cc_368 N_SCE_c_370_n N_A_222_131#_M1041_g 0.017773f $X=3.765 $Y=1.365 $X2=0
+ $Y2=0
cc_369 SCE N_A_222_131#_c_524_n 0.00405447f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_370 N_SCE_c_370_n N_A_222_131#_c_524_n 0.00421201f $X=3.765 $Y=1.365 $X2=0
+ $Y2=0
cc_371 N_SCE_c_371_n N_A_222_131#_c_524_n 0.00490853f $X=3.485 $Y=1.535 $X2=0
+ $Y2=0
cc_372 N_SCE_c_370_n N_A_222_131#_c_525_n 0.00200107f $X=3.765 $Y=1.365 $X2=0
+ $Y2=0
cc_373 N_SCE_c_371_n N_A_222_131#_c_525_n 0.0341293f $X=3.485 $Y=1.535 $X2=0
+ $Y2=0
cc_374 N_SCE_c_360_n N_A_222_131#_c_526_n 0.0115077f $X=1.515 $Y=0.35 $X2=0
+ $Y2=0
cc_375 N_SCE_c_364_n N_A_222_131#_c_526_n 0.0470714f $X=1.6 $Y=1.275 $X2=0 $Y2=0
cc_376 N_SCE_c_365_n N_A_222_131#_c_526_n 0.0137874f $X=1.685 $Y=1.36 $X2=0
+ $Y2=0
cc_377 N_SCE_c_366_n N_A_222_131#_c_526_n 0.0794443f $X=0.82 $Y=1.295 $X2=0
+ $Y2=0
cc_378 N_SCE_M1029_g N_A_222_131#_c_526_n 0.0425357f $X=0.86 $Y=0.865 $X2=0
+ $Y2=0
cc_379 N_SCE_c_381_n N_A_222_131#_c_534_n 0.00383716f $X=1.6 $Y=2.83 $X2=0 $Y2=0
cc_380 N_SCE_c_380_n N_A_222_131#_c_538_n 0.0657963f $X=2.875 $Y=2.75 $X2=0
+ $Y2=0
cc_381 N_SCE_c_387_p N_A_222_131#_c_538_n 0.0179351f $X=1.64 $Y=2.75 $X2=0 $Y2=0
cc_382 N_SCE_c_381_n N_A_222_131#_c_538_n 0.0140105f $X=1.6 $Y=2.83 $X2=0 $Y2=0
cc_383 N_SCE_c_383_n N_A_222_131#_c_538_n 0.00117449f $X=3.385 $Y=2.685 $X2=0
+ $Y2=0
cc_384 SCE N_A_222_131#_c_527_n 0.00644306f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_385 N_SCE_c_370_n N_A_222_131#_c_527_n 0.00353685f $X=3.765 $Y=1.365 $X2=0
+ $Y2=0
cc_386 N_SCE_c_371_n N_A_222_131#_c_527_n 0.0241199f $X=3.485 $Y=1.535 $X2=0
+ $Y2=0
cc_387 N_SCE_c_378_n N_A_222_131#_c_528_n 0.0225466f $X=3.385 $Y=2.565 $X2=0
+ $Y2=0
cc_388 N_SCE_c_380_n N_A_222_131#_c_528_n 2.5052e-19 $X=2.875 $Y=2.75 $X2=0
+ $Y2=0
cc_389 SCE N_A_222_131#_c_528_n 4.11596e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_390 N_SCE_c_383_n N_A_222_131#_c_528_n 0.0173127f $X=3.385 $Y=2.685 $X2=0
+ $Y2=0
cc_391 N_SCE_c_370_n N_A_222_131#_c_528_n 0.0225466f $X=3.765 $Y=1.365 $X2=0
+ $Y2=0
cc_392 N_SCE_c_371_n N_A_222_131#_c_528_n 4.74455e-19 $X=3.485 $Y=1.535 $X2=0
+ $Y2=0
cc_393 N_SCE_c_378_n N_A_222_131#_c_540_n 0.0168532f $X=3.385 $Y=2.565 $X2=0
+ $Y2=0
cc_394 N_SCE_c_383_n N_A_222_131#_c_540_n 0.0065882f $X=3.385 $Y=2.685 $X2=0
+ $Y2=0
cc_395 N_SCE_c_378_n N_A_222_131#_c_575_n 0.00508459f $X=3.385 $Y=2.565 $X2=0
+ $Y2=0
cc_396 N_SCE_c_383_n N_A_222_131#_c_575_n 0.00703784f $X=3.385 $Y=2.685 $X2=0
+ $Y2=0
cc_397 N_SCE_c_383_n N_A_222_131#_c_541_n 0.00514119f $X=3.385 $Y=2.685 $X2=0
+ $Y2=0
cc_398 N_SCE_M1016_g N_A_222_131#_c_542_n 4.2355e-19 $X=2.94 $Y=3.485 $X2=0
+ $Y2=0
cc_399 N_SCE_c_380_n N_A_222_131#_c_542_n 0.0112422f $X=2.875 $Y=2.75 $X2=0
+ $Y2=0
cc_400 N_SCE_c_383_n N_A_222_131#_c_542_n 0.00707069f $X=3.385 $Y=2.685 $X2=0
+ $Y2=0
cc_401 N_SCE_M1029_g N_A_222_131#_c_544_n 0.00895276f $X=0.86 $Y=0.865 $X2=0
+ $Y2=0
cc_402 N_SCE_M1018_g N_A_222_131#_c_545_n 0.00694551f $X=0.86 $Y=3.455 $X2=0
+ $Y2=0
cc_403 N_SCE_c_387_p N_A_222_131#_c_545_n 0.0220177f $X=1.64 $Y=2.75 $X2=0 $Y2=0
cc_404 N_SCE_c_381_n N_A_222_131#_c_545_n 0.0452113f $X=1.6 $Y=2.83 $X2=0 $Y2=0
cc_405 N_SCE_M1029_g N_A_222_131#_c_545_n 0.00578772f $X=0.86 $Y=0.865 $X2=0
+ $Y2=0
cc_406 N_SCE_c_380_n N_A_222_131#_c_546_n 0.0239577f $X=2.875 $Y=2.75 $X2=0
+ $Y2=0
cc_407 N_SCE_c_383_n N_A_222_131#_c_546_n 0.003102f $X=3.385 $Y=2.685 $X2=0
+ $Y2=0
cc_408 N_SCE_M1016_g N_SCD_c_659_n 0.0222883f $X=2.94 $Y=3.485 $X2=0 $Y2=0
cc_409 N_SCE_c_383_n N_SCD_c_659_n 0.00199942f $X=3.385 $Y=2.685 $X2=0 $Y2=0
cc_410 N_SCE_M1016_g N_SCD_c_662_n 0.00643804f $X=2.94 $Y=3.485 $X2=0 $Y2=0
cc_411 N_SCE_c_383_n N_SCD_c_662_n 0.0217794f $X=3.385 $Y=2.685 $X2=0 $Y2=0
cc_412 SCE N_SCD_c_663_n 0.0121162f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_413 N_SCE_c_370_n N_SCD_c_663_n 0.00117175f $X=3.765 $Y=1.365 $X2=0 $Y2=0
cc_414 N_SCE_c_378_n N_SCD_c_664_n 0.00529159f $X=3.385 $Y=2.565 $X2=0 $Y2=0
cc_415 SCE N_SCD_c_664_n 0.0267f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_416 N_SCE_c_370_n N_SCD_c_664_n 0.00277646f $X=3.765 $Y=1.365 $X2=0 $Y2=0
cc_417 N_SCE_c_378_n N_SCD_c_665_n 0.0217794f $X=3.385 $Y=2.565 $X2=0 $Y2=0
cc_418 SCE N_SCD_c_665_n 2.69084e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_419 N_SCE_c_370_n N_SCD_c_665_n 0.0182974f $X=3.765 $Y=1.365 $X2=0 $Y2=0
cc_420 N_SCE_M1031_g N_SCD_M1035_g 0.104206f $X=3.83 $Y=0.745 $X2=10.08 $Y2=0
cc_421 SCE N_SCD_M1035_g 0.00440584f $X=3.995 $Y=1.58 $X2=10.08 $Y2=0
cc_422 SCE N_SCD_c_682_n 0.0404057f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_423 N_SCE_c_370_n N_SCD_c_682_n 0.00104263f $X=3.765 $Y=1.365 $X2=0 $Y2=0
cc_424 N_SCE_M1018_g N_VPWR_c_1922_n 0.0442032f $X=0.86 $Y=3.455 $X2=0 $Y2=0
cc_425 N_SCE_M1016_g N_VPWR_c_1925_n 0.0295211f $X=2.94 $Y=3.485 $X2=0 $Y2=0
cc_426 N_SCE_M1018_g N_VPWR_c_1949_n 0.0133887f $X=0.86 $Y=3.455 $X2=0 $Y2=0
cc_427 N_SCE_M1016_g N_VPWR_c_1949_n 0.00205099f $X=2.94 $Y=3.485 $X2=0 $Y2=0
cc_428 N_SCE_c_380_n N_VPWR_c_1949_n 0.00137427f $X=2.875 $Y=2.75 $X2=0 $Y2=0
cc_429 N_SCE_c_387_p N_VPWR_c_1949_n 0.00628336f $X=1.64 $Y=2.75 $X2=0 $Y2=0
cc_430 N_SCE_c_381_n N_VPWR_c_1949_n 0.00852263f $X=1.6 $Y=2.83 $X2=0 $Y2=0
cc_431 N_SCE_M1016_g N_A_339_655#_c_2087_n 0.0266484f $X=2.94 $Y=3.485 $X2=19.92
+ $Y2=0
cc_432 N_SCE_c_380_n N_A_339_655#_c_2087_n 0.0597401f $X=2.875 $Y=2.75 $X2=19.92
+ $Y2=0
cc_433 N_SCE_c_383_n N_A_339_655#_c_2087_n 0.00320259f $X=3.385 $Y=2.685
+ $X2=19.92 $Y2=0
cc_434 N_SCE_M1018_g N_A_339_655#_c_2088_n 0.00115309f $X=0.86 $Y=3.455
+ $X2=19.92 $Y2=0
cc_435 N_SCE_M1016_g N_A_339_655#_c_2088_n 0.00107129f $X=2.94 $Y=3.485
+ $X2=19.92 $Y2=0
cc_436 N_SCE_c_380_n N_A_339_655#_c_2088_n 0.0195714f $X=2.875 $Y=2.75 $X2=19.92
+ $Y2=0
cc_437 N_SCE_c_387_p N_A_339_655#_c_2088_n 0.00523649f $X=1.64 $Y=2.75 $X2=19.92
+ $Y2=0
cc_438 N_SCE_c_381_n N_A_339_655#_c_2088_n 0.00394668f $X=1.6 $Y=2.83 $X2=19.92
+ $Y2=0
cc_439 N_SCE_M1031_g N_A_339_655#_c_2080_n 0.0272142f $X=3.83 $Y=0.745 $X2=0
+ $Y2=0
cc_440 SCE N_A_339_655#_c_2080_n 0.0427121f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_441 N_SCE_M1031_g N_A_339_655#_c_2085_n 0.0106383f $X=3.83 $Y=0.745 $X2=0
+ $Y2=0
cc_442 N_SCE_c_370_n N_A_339_655#_c_2085_n 0.00120044f $X=3.765 $Y=1.365 $X2=0
+ $Y2=0
cc_443 N_SCE_c_371_n N_A_339_655#_c_2085_n 0.0260738f $X=3.485 $Y=1.535 $X2=0
+ $Y2=0
cc_444 N_SCE_c_362_n N_VGND_c_2294_n 0.00488232f $X=0.985 $Y=0.35 $X2=0 $Y2=0
cc_445 N_SCE_c_366_n N_VGND_c_2294_n 0.0470194f $X=0.82 $Y=1.295 $X2=0 $Y2=0
cc_446 N_SCE_M1029_g N_VGND_c_2294_n 0.0155663f $X=0.86 $Y=0.865 $X2=0 $Y2=0
cc_447 N_SCE_M1031_g N_VGND_c_2308_n 0.00877628f $X=3.83 $Y=0.745 $X2=0 $Y2=0
cc_448 N_SCE_c_360_n N_VGND_c_2308_n 0.0280262f $X=1.515 $Y=0.35 $X2=0 $Y2=0
cc_449 N_SCE_c_362_n N_VGND_c_2308_n 0.00777234f $X=0.985 $Y=0.35 $X2=0 $Y2=0
cc_450 N_SCE_c_364_n N_VGND_c_2308_n 0.0194693f $X=1.6 $Y=1.275 $X2=0 $Y2=0
cc_451 N_SCE_c_366_n N_VGND_c_2308_n 0.0192322f $X=0.82 $Y=1.295 $X2=0 $Y2=0
cc_452 N_SCE_M1029_g N_VGND_c_2308_n 0.0192291f $X=0.86 $Y=0.865 $X2=0 $Y2=0
cc_453 N_SCE_c_364_n N_noxref_25_c_2431_n 0.0396594f $X=1.6 $Y=1.275 $X2=0 $Y2=0
cc_454 N_SCE_c_371_n N_noxref_25_c_2431_n 0.0145801f $X=3.485 $Y=1.535 $X2=0
+ $Y2=0
cc_455 N_SCE_M1031_g N_noxref_25_c_2432_n 0.0190332f $X=3.83 $Y=0.745 $X2=0.24
+ $Y2=0
cc_456 N_SCE_c_360_n N_noxref_25_c_2434_n 0.0119651f $X=1.515 $Y=0.35 $X2=0
+ $Y2=0
cc_457 N_SCE_M1031_g N_noxref_25_c_2436_n 0.00125914f $X=3.83 $Y=0.745 $X2=0
+ $Y2=0
cc_458 N_D_M1040_g N_A_222_131#_M1041_g 0.0371346f $X=2.34 $Y=0.745 $X2=0 $Y2=0
cc_459 N_D_c_484_n N_A_222_131#_c_525_n 0.0474352f $X=2.23 $Y=1.775 $X2=0 $Y2=0
cc_460 N_D_c_484_n N_A_222_131#_c_526_n 0.00397721f $X=2.23 $Y=1.775 $X2=0 $Y2=0
cc_461 N_D_M1001_g N_A_222_131#_c_526_n 0.00437459f $X=2.23 $Y=3.485 $X2=0 $Y2=0
cc_462 N_D_c_487_n N_A_222_131#_c_526_n 0.0346976f $X=2.165 $Y=1.71 $X2=0 $Y2=0
cc_463 N_D_M1001_g N_A_222_131#_c_534_n 9.36896e-19 $X=2.23 $Y=3.485 $X2=0 $Y2=0
cc_464 N_D_M1001_g N_A_222_131#_c_538_n 0.0348898f $X=2.23 $Y=3.485 $X2=0 $Y2=0
cc_465 N_D_c_487_n N_A_222_131#_c_538_n 0.0574705f $X=2.165 $Y=1.71 $X2=0 $Y2=0
cc_466 N_D_c_484_n N_A_222_131#_c_527_n 0.00353229f $X=2.23 $Y=1.775 $X2=0 $Y2=0
cc_467 N_D_c_487_n N_A_222_131#_c_527_n 0.0202537f $X=2.165 $Y=1.71 $X2=0 $Y2=0
cc_468 N_D_c_484_n N_A_222_131#_c_528_n 0.018581f $X=2.23 $Y=1.775 $X2=0 $Y2=0
cc_469 N_D_M1001_g N_A_222_131#_c_528_n 0.018581f $X=2.23 $Y=3.485 $X2=0 $Y2=0
cc_470 N_D_c_487_n N_A_222_131#_c_528_n 0.00150468f $X=2.165 $Y=1.71 $X2=0 $Y2=0
cc_471 N_D_M1001_g N_A_222_131#_c_545_n 0.00389178f $X=2.23 $Y=3.485 $X2=0 $Y2=0
cc_472 N_D_M1001_g N_VPWR_c_1925_n 0.00370609f $X=2.23 $Y=3.485 $X2=0 $Y2=0
cc_473 N_D_M1001_g N_VPWR_c_1949_n 0.0120734f $X=2.23 $Y=3.485 $X2=0 $Y2=0
cc_474 N_D_M1001_g N_A_339_655#_c_2087_n 0.0184504f $X=2.23 $Y=3.485 $X2=19.92
+ $Y2=0
cc_475 N_D_M1001_g N_A_339_655#_c_2088_n 0.0253152f $X=2.23 $Y=3.485 $X2=19.92
+ $Y2=0
cc_476 N_D_M1040_g N_A_339_655#_c_2085_n 0.00147895f $X=2.34 $Y=0.745 $X2=0
+ $Y2=0
cc_477 N_D_M1040_g N_VGND_c_2308_n 0.023887f $X=2.34 $Y=0.745 $X2=0 $Y2=0
cc_478 N_D_M1040_g N_noxref_25_c_2431_n 0.0170961f $X=2.34 $Y=0.745 $X2=0 $Y2=0
cc_479 N_D_M1040_g N_noxref_25_c_2432_n 0.0210753f $X=2.34 $Y=0.745 $X2=0.24
+ $Y2=0
cc_480 N_D_M1040_g N_noxref_25_c_2434_n 0.00106498f $X=2.34 $Y=0.745 $X2=0 $Y2=0
cc_481 N_A_222_131#_M1006_g N_SCD_c_659_n 0.0380025f $X=4.43 $Y=3.485 $X2=0
+ $Y2=0
cc_482 N_A_222_131#_c_541_n N_SCD_c_659_n 0.00567281f $X=4.35 $Y=2.75 $X2=0
+ $Y2=0
cc_483 N_A_222_131#_c_529_n N_SCD_c_662_n 0.0380025f $X=4.43 $Y=3.02 $X2=0 $Y2=0
cc_484 N_A_222_131#_c_541_n N_SCD_c_662_n 0.0153286f $X=4.35 $Y=2.75 $X2=0 $Y2=0
cc_485 N_A_222_131#_c_606_p N_SCD_c_662_n 6.46987e-19 $X=4.515 $Y=2.41 $X2=0
+ $Y2=0
cc_486 N_A_222_131#_c_543_n N_SCD_c_662_n 0.00690443f $X=4.515 $Y=2.41 $X2=0
+ $Y2=0
cc_487 N_A_222_131#_c_529_n N_SCD_c_663_n 7.88027e-19 $X=4.43 $Y=3.02 $X2=0
+ $Y2=0
cc_488 N_A_222_131#_c_541_n N_SCD_c_663_n 0.0109417f $X=4.35 $Y=2.75 $X2=0 $Y2=0
cc_489 N_A_222_131#_c_606_p N_SCD_c_663_n 0.0018443f $X=4.515 $Y=2.41 $X2=0
+ $Y2=0
cc_490 N_A_222_131#_c_543_n N_SCD_c_663_n 2.10134e-19 $X=4.515 $Y=2.41 $X2=0
+ $Y2=0
cc_491 N_A_222_131#_c_527_n N_SCD_c_664_n 0.00890027f $X=2.895 $Y=1.79 $X2=0
+ $Y2=0
cc_492 N_A_222_131#_c_540_n N_SCD_c_664_n 0.00908468f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_493 N_A_222_131#_c_541_n N_SCD_c_664_n 0.0230282f $X=4.35 $Y=2.75 $X2=0 $Y2=0
cc_494 N_A_222_131#_c_606_p N_SCD_c_664_n 0.0071927f $X=4.515 $Y=2.41 $X2=0
+ $Y2=0
cc_495 N_A_222_131#_c_543_n N_SCD_c_664_n 0.00115523f $X=4.515 $Y=2.41 $X2=0
+ $Y2=0
cc_496 N_A_222_131#_c_540_n N_SCD_c_665_n 5.5474e-19 $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_497 N_A_222_131#_c_575_n N_SCD_c_665_n 0.00109688f $X=3.355 $Y=2.665 $X2=0
+ $Y2=0
cc_498 N_A_222_131#_c_541_n N_SCD_c_665_n 0.00181832f $X=4.35 $Y=2.75 $X2=0
+ $Y2=0
cc_499 N_A_222_131#_c_606_p N_SCD_c_665_n 0.00115523f $X=4.515 $Y=2.41 $X2=0
+ $Y2=0
cc_500 N_A_222_131#_c_543_n N_SCD_c_665_n 0.0130598f $X=4.515 $Y=2.41 $X2=0
+ $Y2=0
cc_501 N_A_222_131#_c_541_n N_SCD_M1035_g 2.42746e-19 $X=4.35 $Y=2.75 $X2=10.08
+ $Y2=0
cc_502 N_A_222_131#_c_606_p N_SCD_M1035_g 2.73118e-19 $X=4.515 $Y=2.41 $X2=10.08
+ $Y2=0
cc_503 N_A_222_131#_c_543_n N_SCD_M1035_g 0.0164614f $X=4.515 $Y=2.41 $X2=10.08
+ $Y2=0
cc_504 N_A_222_131#_c_606_p N_SCD_c_667_n 0.026549f $X=4.515 $Y=2.41 $X2=0 $Y2=0
cc_505 N_A_222_131#_c_543_n N_SCD_c_667_n 0.00271367f $X=4.515 $Y=2.41 $X2=0
+ $Y2=0
cc_506 N_A_222_131#_c_529_n N_RESET_B_c_1302_n 0.015004f $X=4.43 $Y=3.02 $X2=0
+ $Y2=0
cc_507 N_A_222_131#_c_543_n N_RESET_B_c_1302_n 0.015004f $X=4.515 $Y=2.41 $X2=0
+ $Y2=0
cc_508 N_A_222_131#_c_543_n N_RESET_B_c_1291_n 0.0107124f $X=4.515 $Y=2.41 $X2=0
+ $Y2=0
cc_509 N_A_222_131#_c_534_n N_VPWR_c_1922_n 0.0241554f $X=1.29 $Y=3.33 $X2=0
+ $Y2=0
cc_510 N_A_222_131#_M1006_g N_VPWR_c_1925_n 0.0016215f $X=4.43 $Y=3.485 $X2=0
+ $Y2=0
cc_511 N_A_222_131#_M1006_g N_VPWR_c_1928_n 4.28529e-19 $X=4.43 $Y=3.485 $X2=0
+ $Y2=0
cc_512 N_A_222_131#_M1018_d N_VPWR_c_1949_n 9.58863e-19 $X=1.11 $Y=3.245 $X2=0
+ $Y2=0
cc_513 N_A_222_131#_M1006_g N_VPWR_c_1949_n 0.0149341f $X=4.43 $Y=3.485 $X2=0
+ $Y2=0
cc_514 N_A_222_131#_c_535_n N_VPWR_c_1949_n 0.022651f $X=1.25 $Y=3.455 $X2=0
+ $Y2=0
cc_515 N_A_222_131#_c_541_n N_VPWR_c_1949_n 5.32817e-19 $X=4.35 $Y=2.75 $X2=0
+ $Y2=0
cc_516 N_A_222_131#_c_529_n N_A_339_655#_c_2087_n 0.00684817f $X=4.43 $Y=3.02
+ $X2=19.92 $Y2=0
cc_517 N_A_222_131#_M1006_g N_A_339_655#_c_2087_n 0.0166119f $X=4.43 $Y=3.485
+ $X2=19.92 $Y2=0
cc_518 N_A_222_131#_c_540_n N_A_339_655#_c_2087_n 0.00661822f $X=3.27 $Y=2.4
+ $X2=19.92 $Y2=0
cc_519 N_A_222_131#_c_541_n N_A_339_655#_c_2087_n 0.0808255f $X=4.35 $Y=2.75
+ $X2=19.92 $Y2=0
cc_520 N_A_222_131#_c_542_n N_A_339_655#_c_2087_n 0.013083f $X=3.44 $Y=2.75
+ $X2=19.92 $Y2=0
cc_521 N_A_222_131#_c_546_n N_A_339_655#_c_2087_n 6.86039e-19 $X=2.895 $Y=2.4
+ $X2=19.92 $Y2=0
cc_522 N_A_222_131#_c_534_n N_A_339_655#_c_2088_n 0.0265055f $X=1.29 $Y=3.33
+ $X2=19.92 $Y2=0
cc_523 N_A_222_131#_c_545_n N_A_339_655#_c_2088_n 0.00609345f $X=1.29 $Y=3.205
+ $X2=19.92 $Y2=0
cc_524 N_A_222_131#_M1006_g N_A_339_655#_c_2091_n 0.0150613f $X=4.43 $Y=3.485
+ $X2=0 $Y2=0
cc_525 N_A_222_131#_c_529_n N_A_339_655#_c_2081_n 0.00382155f $X=4.43 $Y=3.02
+ $X2=0 $Y2=0
cc_526 N_A_222_131#_c_541_n N_A_339_655#_c_2081_n 0.0117527f $X=4.35 $Y=2.75
+ $X2=0 $Y2=0
cc_527 N_A_222_131#_c_606_p N_A_339_655#_c_2081_n 0.0221705f $X=4.515 $Y=2.41
+ $X2=0 $Y2=0
cc_528 N_A_222_131#_c_543_n N_A_339_655#_c_2081_n 0.00483217f $X=4.515 $Y=2.41
+ $X2=0 $Y2=0
cc_529 N_A_222_131#_M1041_g N_A_339_655#_c_2085_n 0.0138204f $X=3.05 $Y=0.745
+ $X2=0 $Y2=0
cc_530 N_A_222_131#_c_529_n N_A_339_655#_c_2111_n 4.24501e-19 $X=4.43 $Y=3.02
+ $X2=0 $Y2=0
cc_531 N_A_222_131#_M1006_g N_A_339_655#_c_2111_n 0.00256019f $X=4.43 $Y=3.485
+ $X2=0 $Y2=0
cc_532 N_A_222_131#_c_541_n N_A_339_655#_c_2111_n 0.00193497f $X=4.35 $Y=2.75
+ $X2=0 $Y2=0
cc_533 N_A_222_131#_M1041_g N_VGND_c_2308_n 0.0247522f $X=3.05 $Y=0.745 $X2=0
+ $Y2=0
cc_534 N_A_222_131#_c_526_n N_VGND_c_2308_n 0.0118584f $X=1.25 $Y=0.865 $X2=0
+ $Y2=0
cc_535 N_A_222_131#_M1041_g N_noxref_25_c_2431_n 0.00196443f $X=3.05 $Y=0.745
+ $X2=0 $Y2=0
cc_536 N_A_222_131#_M1041_g N_noxref_25_c_2432_n 0.0221759f $X=3.05 $Y=0.745
+ $X2=0.24 $Y2=0
cc_537 N_SCD_M1035_g N_RESET_B_M1007_g 0.0199951f $X=4.54 $Y=0.745 $X2=0 $Y2=0
cc_538 N_SCD_M1035_g N_RESET_B_c_1296_n 0.0338529f $X=4.54 $Y=0.745 $X2=0 $Y2=0
cc_539 N_SCD_c_659_n N_VPWR_c_1925_n 0.0102333f $X=3.72 $Y=3.265 $X2=0 $Y2=0
cc_540 N_SCD_c_659_n N_VPWR_c_1949_n 0.0146093f $X=3.72 $Y=3.265 $X2=0 $Y2=0
cc_541 N_SCD_c_659_n N_A_339_655#_c_2087_n 0.0244898f $X=3.72 $Y=3.265 $X2=19.92
+ $Y2=0
cc_542 N_SCD_M1035_g N_A_339_655#_c_2080_n 0.0351796f $X=4.54 $Y=0.745 $X2=0
+ $Y2=0
cc_543 N_SCD_c_682_n N_A_339_655#_c_2080_n 0.0219216f $X=4.54 $Y=1.46 $X2=0
+ $Y2=0
cc_544 N_SCD_c_659_n N_A_339_655#_c_2091_n 0.00206755f $X=3.72 $Y=3.265 $X2=0
+ $Y2=0
cc_545 N_SCD_M1035_g N_A_339_655#_c_2081_n 0.0102824f $X=4.54 $Y=0.745 $X2=0
+ $Y2=0
cc_546 N_SCD_c_682_n N_A_339_655#_c_2081_n 0.0489102f $X=4.54 $Y=1.46 $X2=0
+ $Y2=0
cc_547 N_SCD_c_667_n N_A_339_655#_c_2081_n 0.0145257f $X=4.54 $Y=1.975 $X2=0
+ $Y2=0
cc_548 N_SCD_M1035_g N_A_339_655#_c_2085_n 9.9266e-19 $X=4.54 $Y=0.745 $X2=0
+ $Y2=0
cc_549 N_SCD_M1035_g N_VGND_c_2296_n 8.67218e-19 $X=4.54 $Y=0.745 $X2=0 $Y2=0
cc_550 N_SCD_M1035_g N_VGND_c_2308_n 0.00791759f $X=4.54 $Y=0.745 $X2=0 $Y2=0
cc_551 N_SCD_M1035_g N_noxref_25_c_2432_n 0.0180005f $X=4.54 $Y=0.745 $X2=0.24
+ $Y2=0
cc_552 N_SCD_M1035_g N_noxref_25_c_2436_n 0.0103626f $X=4.54 $Y=0.745 $X2=0
+ $Y2=0
cc_553 N_CLK_M1026_g N_A_1290_126#_c_955_n 0.0241246f $X=6.2 $Y=0.84 $X2=0 $Y2=0
cc_554 N_CLK_M1026_g N_A_1290_126#_c_957_n 0.0500142f $X=6.2 $Y=0.84 $X2=0 $Y2=0
cc_555 N_CLK_c_733_p N_A_1290_126#_c_957_n 0.0308305f $X=6.035 $Y=2.015 $X2=0
+ $Y2=0
cc_556 N_CLK_M1026_g N_A_1290_126#_c_961_n 0.00895276f $X=6.2 $Y=0.84 $X2=0
+ $Y2=0
cc_557 N_CLK_M1026_g N_RESET_B_M1007_g 0.03685f $X=6.2 $Y=0.84 $X2=0 $Y2=0
cc_558 N_CLK_M1026_g N_RESET_B_c_1286_n 0.0344733f $X=6.2 $Y=0.84 $X2=0 $Y2=0
cc_559 N_CLK_M1002_g N_RESET_B_c_1302_n 0.0130586f $X=6.2 $Y=3.34 $X2=0 $Y2=0
cc_560 N_CLK_c_726_n N_RESET_B_c_1308_n 0.0260183f $X=6.035 $Y=2.015 $X2=0 $Y2=0
cc_561 N_CLK_c_733_p N_RESET_B_c_1308_n 0.0392651f $X=6.035 $Y=2.015 $X2=0 $Y2=0
cc_562 N_CLK_c_726_n N_RESET_B_c_1309_n 0.00144293f $X=6.035 $Y=2.015 $X2=0
+ $Y2=0
cc_563 N_CLK_c_733_p N_RESET_B_c_1309_n 0.00255234f $X=6.035 $Y=2.015 $X2=0
+ $Y2=0
cc_564 N_CLK_M1026_g N_RESET_B_c_1291_n 0.00668895f $X=6.2 $Y=0.84 $X2=0 $Y2=0
cc_565 N_CLK_M1002_g N_RESET_B_c_1291_n 0.0277678f $X=6.2 $Y=3.34 $X2=0 $Y2=0
cc_566 N_CLK_c_726_n N_RESET_B_c_1291_n 0.0419581f $X=6.035 $Y=2.015 $X2=0 $Y2=0
cc_567 N_CLK_c_733_p N_RESET_B_c_1291_n 0.00298598f $X=6.035 $Y=2.015 $X2=0
+ $Y2=0
cc_568 N_CLK_M1026_g N_RESET_B_c_1297_n 0.00640002f $X=6.2 $Y=0.84 $X2=0 $Y2=0
cc_569 N_CLK_c_726_n N_RESET_B_c_1297_n 0.00381943f $X=6.035 $Y=2.015 $X2=0
+ $Y2=0
cc_570 N_CLK_c_733_p N_RESET_B_c_1297_n 0.015539f $X=6.035 $Y=2.015 $X2=0 $Y2=0
cc_571 N_CLK_M1002_g N_VPWR_c_1928_n 0.00560162f $X=6.2 $Y=3.34 $X2=0 $Y2=0
cc_572 N_CLK_M1002_g N_VPWR_c_1949_n 0.0126791f $X=6.2 $Y=3.34 $X2=0 $Y2=0
cc_573 N_CLK_M1002_g N_A_339_655#_c_2095_n 0.0259541f $X=6.2 $Y=3.34 $X2=0 $Y2=0
cc_574 N_CLK_c_726_n N_A_339_655#_c_2095_n 0.00208994f $X=6.035 $Y=2.015 $X2=0
+ $Y2=0
cc_575 N_CLK_c_733_p N_A_339_655#_c_2095_n 0.00979145f $X=6.035 $Y=2.015 $X2=0
+ $Y2=0
cc_576 N_CLK_M1002_g N_A_339_655#_c_2159_n 0.0173152f $X=6.2 $Y=3.34 $X2=0 $Y2=0
cc_577 N_CLK_M1002_g N_A_339_655#_c_2096_n 0.00907311f $X=6.2 $Y=3.34 $X2=0
+ $Y2=0
cc_578 N_CLK_M1002_g N_A_339_655#_c_2099_n 0.00503226f $X=6.2 $Y=3.34 $X2=0
+ $Y2=0
cc_579 N_CLK_M1002_g N_A_339_655#_c_2101_n 0.00440111f $X=6.2 $Y=3.34 $X2=0
+ $Y2=0
cc_580 N_CLK_M1026_g N_VGND_c_2296_n 0.0360595f $X=6.2 $Y=0.84 $X2=0 $Y2=0
cc_581 N_CLK_M1026_g N_VGND_c_2308_n 0.0138207f $X=6.2 $Y=0.84 $X2=0 $Y2=0
cc_582 N_A_1569_126#_c_781_n N_A_1290_126#_M1019_g 0.0174791f $X=8.83 $Y=3.185
+ $X2=0 $Y2=0
cc_583 N_A_1569_126#_c_761_n N_A_1290_126#_M1019_g 0.0172042f $X=8.027 $Y=2.225
+ $X2=0 $Y2=0
cc_584 N_A_1569_126#_c_787_n N_A_1290_126#_M1019_g 0.0157755f $X=8.07 $Y=2.39
+ $X2=0 $Y2=0
cc_585 N_A_1569_126#_c_761_n N_A_1290_126#_c_948_n 0.0301468f $X=8.027 $Y=2.225
+ $X2=0 $Y2=0
cc_586 N_A_1569_126#_c_762_n N_A_1290_126#_c_948_n 0.00480986f $X=9.7 $Y=0.35
+ $X2=0 $Y2=0
cc_587 N_A_1569_126#_c_787_n N_A_1290_126#_c_948_n 0.0125734f $X=8.07 $Y=2.39
+ $X2=0 $Y2=0
cc_588 N_A_1569_126#_c_760_n N_A_1290_126#_c_949_n 0.00245398f $X=7.985 $Y=0.83
+ $X2=19.92 $Y2=0
cc_589 N_A_1569_126#_c_762_n N_A_1290_126#_c_949_n 0.00537992f $X=9.7 $Y=0.35
+ $X2=19.92 $Y2=0
cc_590 N_A_1569_126#_c_766_n N_A_1290_126#_c_949_n 8.71057e-19 $X=9.837 $Y=0.925
+ $X2=19.92 $Y2=0
cc_591 N_A_1569_126#_c_775_n N_A_1290_126#_c_949_n 0.00166583f $X=8.025 $Y=0.995
+ $X2=19.92 $Y2=0
cc_592 N_A_1569_126#_M1004_g N_A_1290_126#_c_949_n 0.0113842f $X=9.745 $Y=0.84
+ $X2=19.92 $Y2=0
cc_593 N_A_1569_126#_c_781_n N_A_1290_126#_M1037_g 0.0372221f $X=8.83 $Y=3.185
+ $X2=10.08 $Y2=0.057
cc_594 N_A_1569_126#_c_786_n N_A_1290_126#_M1024_g 0.0134603f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_595 N_A_1569_126#_c_801_p N_A_1290_126#_c_951_n 0.00109626f $X=12.91 $Y=1.475
+ $X2=0 $Y2=0
cc_596 N_A_1569_126#_c_772_n N_A_1290_126#_c_951_n 7.2024e-19 $X=14.1 $Y=0.35
+ $X2=0 $Y2=0
cc_597 N_A_1569_126#_c_780_n N_A_1290_126#_c_951_n 0.00779509f $X=12.897
+ $Y=1.395 $X2=0 $Y2=0
cc_598 N_A_1569_126#_c_804_p N_A_1290_126#_c_952_n 7.8279e-19 $X=12.99 $Y=1.56
+ $X2=0 $Y2=0
cc_599 N_A_1569_126#_c_778_n N_A_1290_126#_c_952_n 0.0173552f $X=12.99 $Y=1.56
+ $X2=0 $Y2=0
cc_600 N_A_1569_126#_c_801_p N_A_1290_126#_M1020_g 0.00131853f $X=12.91 $Y=1.475
+ $X2=0 $Y2=0
cc_601 N_A_1569_126#_c_772_n N_A_1290_126#_M1020_g 0.0226495f $X=14.1 $Y=0.35
+ $X2=0 $Y2=0
cc_602 N_A_1569_126#_c_774_n N_A_1290_126#_M1020_g 0.0172514f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_603 N_A_1569_126#_c_780_n N_A_1290_126#_M1020_g 0.0135696f $X=12.897 $Y=1.395
+ $X2=0 $Y2=0
cc_604 N_A_1569_126#_c_810_p N_A_1290_126#_c_954_n 5.81374e-19 $X=9.81 $Y=1.44
+ $X2=0 $Y2=0
cc_605 N_A_1569_126#_M1004_g N_A_1290_126#_c_954_n 0.0421262f $X=9.745 $Y=0.84
+ $X2=0 $Y2=0
cc_606 N_A_1569_126#_c_810_p N_A_1290_126#_c_974_n 0.0017612f $X=9.81 $Y=1.44
+ $X2=0 $Y2=0
cc_607 N_A_1569_126#_M1004_g N_A_1290_126#_c_974_n 0.00288548f $X=9.745 $Y=0.84
+ $X2=0 $Y2=0
cc_608 N_A_1569_126#_c_761_n N_A_1290_126#_c_1011_n 0.0204469f $X=8.027 $Y=2.225
+ $X2=0 $Y2=0
cc_609 N_A_1569_126#_c_810_p N_A_1290_126#_c_1012_n 0.00595897f $X=9.81 $Y=1.44
+ $X2=0 $Y2=0
cc_610 N_A_1569_126#_M1004_g N_A_1290_126#_c_1012_n 0.00305668f $X=9.745 $Y=0.84
+ $X2=0 $Y2=0
cc_611 N_A_1569_126#_c_781_n N_A_1290_126#_c_979_n 0.0189818f $X=8.83 $Y=3.185
+ $X2=0 $Y2=0
cc_612 N_A_1569_126#_c_810_p N_A_1290_126#_c_979_n 4.6244e-19 $X=9.81 $Y=1.44
+ $X2=0 $Y2=0
cc_613 N_A_1569_126#_c_787_n N_A_1290_126#_c_979_n 9.89963e-19 $X=8.07 $Y=2.39
+ $X2=0 $Y2=0
cc_614 N_A_1569_126#_M1004_g N_A_1290_126#_c_979_n 0.0260242f $X=9.745 $Y=0.84
+ $X2=0 $Y2=0
cc_615 N_A_1569_126#_c_761_n N_A_1290_126#_c_962_n 0.02458f $X=8.027 $Y=2.225
+ $X2=0 $Y2=0
cc_616 N_A_1569_126#_c_760_n N_A_1290_126#_c_963_n 0.00297952f $X=7.985 $Y=0.83
+ $X2=0 $Y2=0
cc_617 N_A_1569_126#_c_761_n N_A_1290_126#_c_963_n 0.00522537f $X=8.027 $Y=2.225
+ $X2=0 $Y2=0
cc_618 N_A_1569_126#_c_786_n N_A_1290_126#_c_964_n 0.030583f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_619 N_A_1569_126#_c_778_n N_A_1290_126#_c_964_n 0.0234479f $X=12.99 $Y=1.56
+ $X2=0 $Y2=0
cc_620 N_A_1569_126#_c_767_n N_A_2014_537#_c_1164_n 0.107644f $X=11.975 $Y=1.01
+ $X2=0 $Y2=0
cc_621 N_A_1569_126#_c_767_n N_A_2014_537#_c_1183_n 0.0135702f $X=11.975 $Y=1.01
+ $X2=0 $Y2=0
cc_622 N_A_1569_126#_c_828_p N_A_2014_537#_c_1183_n 0.0220406f $X=12.06 $Y=0.925
+ $X2=0 $Y2=0
cc_623 N_A_1569_126#_c_768_n N_A_2014_537#_c_1183_n 0.0199321f $X=12.825 $Y=0.35
+ $X2=0 $Y2=0
cc_624 N_A_1569_126#_c_801_p N_A_2014_537#_c_1183_n 0.0449134f $X=12.91 $Y=1.475
+ $X2=0 $Y2=0
cc_625 N_A_1569_126#_c_780_n N_A_2014_537#_c_1183_n 0.011946f $X=12.897 $Y=1.395
+ $X2=0 $Y2=0
cc_626 N_A_1569_126#_c_801_p N_A_2014_537#_c_1165_n 0.00190994f $X=12.91
+ $Y=1.475 $X2=0 $Y2=0
cc_627 N_A_1569_126#_c_804_p N_A_2014_537#_c_1165_n 0.0115167f $X=12.99 $Y=1.56
+ $X2=0 $Y2=0
cc_628 N_A_1569_126#_c_778_n N_A_2014_537#_c_1165_n 0.0121443f $X=12.99 $Y=1.56
+ $X2=0 $Y2=0
cc_629 N_A_1569_126#_c_804_p N_A_2014_537#_c_1166_n 0.021033f $X=12.99 $Y=1.56
+ $X2=0 $Y2=0
cc_630 N_A_1569_126#_c_778_n N_A_2014_537#_c_1166_n 0.012388f $X=12.99 $Y=1.56
+ $X2=0 $Y2=0
cc_631 N_A_1569_126#_c_786_n N_A_2014_537#_c_1180_n 4.34669e-19 $X=14.185
+ $Y=2.39 $X2=0 $Y2=0
cc_632 N_A_1569_126#_c_786_n N_A_2014_537#_c_1194_n 3.14784e-19 $X=14.185
+ $Y=2.39 $X2=0 $Y2=0
cc_633 N_A_1569_126#_c_810_p N_A_2014_537#_c_1195_n 0.0264198f $X=9.81 $Y=1.44
+ $X2=0 $Y2=0
cc_634 N_A_1569_126#_c_767_n N_A_2014_537#_c_1195_n 0.0203427f $X=11.975 $Y=1.01
+ $X2=0 $Y2=0
cc_635 N_A_1569_126#_M1004_g N_A_2014_537#_c_1195_n 0.00191729f $X=9.745 $Y=0.84
+ $X2=0 $Y2=0
cc_636 N_A_1569_126#_c_801_p N_A_2014_537#_c_1168_n 0.0122935f $X=12.91 $Y=1.475
+ $X2=0 $Y2=0
cc_637 N_A_1569_126#_c_778_n N_A_2014_537#_c_1168_n 0.00145978f $X=12.99 $Y=1.56
+ $X2=0 $Y2=0
cc_638 N_A_1569_126#_c_780_n N_A_2014_537#_c_1168_n 0.00334023f $X=12.897
+ $Y=1.395 $X2=0 $Y2=0
cc_639 N_A_1569_126#_c_766_n N_A_2014_537#_M1005_g 0.00344233f $X=9.837 $Y=0.925
+ $X2=0 $Y2=0
cc_640 N_A_1569_126#_c_810_p N_A_2014_537#_M1005_g 0.00304607f $X=9.81 $Y=1.44
+ $X2=0 $Y2=0
cc_641 N_A_1569_126#_c_767_n N_A_2014_537#_M1005_g 0.0225786f $X=11.975 $Y=1.01
+ $X2=0 $Y2=0
cc_642 N_A_1569_126#_M1004_g N_A_2014_537#_M1005_g 0.0875347f $X=9.745 $Y=0.84
+ $X2=0 $Y2=0
cc_643 N_A_1569_126#_c_762_n N_RESET_B_c_1286_n 0.0344961f $X=9.7 $Y=0.35 $X2=0
+ $Y2=0
cc_644 N_A_1569_126#_c_764_n N_RESET_B_c_1286_n 0.00841261f $X=8.15 $Y=0.35
+ $X2=0 $Y2=0
cc_645 N_A_1569_126#_c_767_n N_RESET_B_c_1286_n 0.00409475f $X=11.975 $Y=1.01
+ $X2=0 $Y2=0
cc_646 N_A_1569_126#_c_770_n N_RESET_B_c_1286_n 0.0016256f $X=12.145 $Y=0.35
+ $X2=0 $Y2=0
cc_647 N_A_1569_126#_M1004_g N_RESET_B_c_1286_n 0.0333124f $X=9.745 $Y=0.84
+ $X2=0 $Y2=0
cc_648 N_A_1569_126#_c_781_n N_RESET_B_c_1308_n 0.00487693f $X=8.83 $Y=3.185
+ $X2=0 $Y2=0
cc_649 N_A_1569_126#_c_761_n N_RESET_B_c_1308_n 0.0313447f $X=8.027 $Y=2.225
+ $X2=0 $Y2=0
cc_650 N_A_1569_126#_c_810_p N_RESET_B_c_1308_n 0.00764222f $X=9.81 $Y=1.44
+ $X2=0 $Y2=0
cc_651 N_A_1569_126#_c_787_n N_RESET_B_c_1308_n 0.0252208f $X=8.07 $Y=2.39 $X2=0
+ $Y2=0
cc_652 N_A_1569_126#_M1004_g N_RESET_B_c_1308_n 0.00843496f $X=9.745 $Y=0.84
+ $X2=0 $Y2=0
cc_653 N_A_1569_126#_c_774_n N_RESET_B_c_1310_n 0.0168807f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_654 N_A_1569_126#_c_786_n N_RESET_B_c_1310_n 0.00572173f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_655 N_A_1569_126#_c_804_p N_RESET_B_c_1310_n 0.00168243f $X=12.99 $Y=1.56
+ $X2=0 $Y2=0
cc_656 N_A_1569_126#_c_767_n N_RESET_B_M1008_g 0.026117f $X=11.975 $Y=1.01 $X2=0
+ $Y2=0
cc_657 N_A_1569_126#_c_828_p N_RESET_B_M1008_g 0.00118983f $X=12.06 $Y=0.925
+ $X2=0 $Y2=0
cc_658 N_A_1569_126#_c_767_n N_A_1816_659#_M1039_g 0.0166108f $X=11.975 $Y=1.01
+ $X2=0 $Y2=0
cc_659 N_A_1569_126#_c_828_p N_A_1816_659#_M1039_g 0.0203472f $X=12.06 $Y=0.925
+ $X2=0 $Y2=0
cc_660 N_A_1569_126#_c_768_n N_A_1816_659#_M1039_g 0.0084765f $X=12.825 $Y=0.35
+ $X2=0 $Y2=0
cc_661 N_A_1569_126#_c_770_n N_A_1816_659#_M1039_g 0.00354446f $X=12.145 $Y=0.35
+ $X2=0 $Y2=0
cc_662 N_A_1569_126#_c_801_p N_A_1816_659#_M1039_g 0.00134252f $X=12.91 $Y=1.475
+ $X2=0 $Y2=0
cc_663 N_A_1569_126#_c_780_n N_A_1816_659#_M1039_g 0.0320979f $X=12.897 $Y=1.395
+ $X2=0 $Y2=0
cc_664 N_A_1569_126#_c_781_n N_A_1816_659#_c_1500_n 0.00192063f $X=8.83 $Y=3.185
+ $X2=0 $Y2=0
cc_665 N_A_1569_126#_c_810_p N_A_1816_659#_c_1500_n 0.026024f $X=9.81 $Y=1.44
+ $X2=0 $Y2=0
cc_666 N_A_1569_126#_c_872_p N_A_1816_659#_c_1500_n 0.00415011f $X=9.837 $Y=1.01
+ $X2=0 $Y2=0
cc_667 N_A_1569_126#_M1004_g N_A_1816_659#_c_1500_n 0.00619435f $X=9.745 $Y=0.84
+ $X2=0 $Y2=0
cc_668 N_A_1569_126#_c_781_n N_A_1816_659#_c_1507_n 0.00342635f $X=8.83 $Y=3.185
+ $X2=0 $Y2=0
cc_669 N_A_1569_126#_c_762_n N_A_1816_659#_c_1501_n 0.0256136f $X=9.7 $Y=0.35
+ $X2=0 $Y2=0
cc_670 N_A_1569_126#_c_766_n N_A_1816_659#_c_1501_n 0.0220895f $X=9.837 $Y=0.925
+ $X2=0 $Y2=0
cc_671 N_A_1569_126#_c_872_p N_A_1816_659#_c_1501_n 0.00534495f $X=9.837 $Y=1.01
+ $X2=0 $Y2=0
cc_672 N_A_1569_126#_M1004_g N_A_1816_659#_c_1501_n 0.00790084f $X=9.745 $Y=0.84
+ $X2=0 $Y2=0
cc_673 N_A_1569_126#_c_781_n N_A_1816_659#_c_1516_n 0.00171697f $X=8.83 $Y=3.185
+ $X2=0 $Y2=0
cc_674 N_A_1569_126#_c_778_n N_A_1816_659#_c_1517_n 0.00269412f $X=12.99 $Y=1.56
+ $X2=0 $Y2=0
cc_675 N_A_1569_126#_c_772_n N_A_2841_81#_c_1618_n 0.00180985f $X=14.1 $Y=0.35
+ $X2=0 $Y2=0
cc_676 N_A_1569_126#_c_774_n N_A_2841_81#_c_1618_n 0.0188799f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_677 N_A_1569_126#_c_774_n N_A_2841_81#_c_1620_n 0.0138399f $X=14.185 $Y=2.39
+ $X2=19.92 $Y2=0
cc_678 N_A_1569_126#_c_786_n N_A_2841_81#_c_1620_n 0.00247062f $X=14.185 $Y=2.39
+ $X2=19.92 $Y2=0
cc_679 N_A_1569_126#_c_774_n N_A_2841_81#_c_1624_n 0.00261922f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_680 N_A_1569_126#_c_786_n N_A_2841_81#_c_1624_n 0.07036f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_681 N_A_1569_126#_c_801_p N_A_2624_107#_c_1723_n 0.00593071f $X=12.91
+ $Y=1.475 $X2=0 $Y2=0
cc_682 N_A_1569_126#_c_801_p N_A_2624_107#_c_1724_n 0.016659f $X=12.91 $Y=1.475
+ $X2=0 $Y2=0
cc_683 N_A_1569_126#_c_772_n N_A_2624_107#_c_1724_n 0.0166099f $X=14.1 $Y=0.35
+ $X2=0 $Y2=0
cc_684 N_A_1569_126#_c_774_n N_A_2624_107#_c_1724_n 0.013651f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_685 N_A_1569_126#_c_774_n N_A_2624_107#_c_1725_n 0.0130062f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_686 N_A_1569_126#_c_786_n N_A_2624_107#_c_1736_n 0.00635253f $X=14.185
+ $Y=2.39 $X2=0 $Y2=0
cc_687 N_A_1569_126#_c_774_n N_A_2624_107#_c_1739_n 0.084941f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_688 N_A_1569_126#_c_786_n N_A_2624_107#_c_1739_n 0.0207129f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_689 N_A_1569_126#_c_804_p N_A_2624_107#_c_1739_n 0.00426493f $X=12.99 $Y=1.56
+ $X2=0 $Y2=0
cc_690 N_A_1569_126#_c_778_n N_A_2624_107#_c_1739_n 0.00138611f $X=12.99 $Y=1.56
+ $X2=0 $Y2=0
cc_691 N_A_1569_126#_c_780_n N_A_2624_107#_c_1739_n 4.13625e-19 $X=12.897
+ $Y=1.395 $X2=0 $Y2=0
cc_692 N_A_1569_126#_c_774_n N_A_2624_107#_c_1752_n 0.00769616f $X=14.185
+ $Y=2.39 $X2=0 $Y2=0
cc_693 N_A_1569_126#_c_786_n N_A_2624_107#_c_1752_n 0.0307386f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_694 N_A_1569_126#_c_774_n N_A_2624_107#_c_1726_n 0.090153f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_695 N_A_1569_126#_c_786_n N_A_2624_107#_c_1726_n 0.00576163f $X=14.185
+ $Y=2.39 $X2=0 $Y2=0
cc_696 N_A_1569_126#_c_774_n N_A_2624_107#_c_1756_n 0.0123662f $X=14.185 $Y=2.39
+ $X2=0 $Y2=0
cc_697 N_A_1569_126#_c_786_n N_A_2624_107#_c_1757_n 0.00500048f $X=14.185
+ $Y=2.39 $X2=0 $Y2=0
cc_698 N_A_1569_126#_c_786_n N_VPWR_c_1940_n 0.00114203f $X=14.185 $Y=2.39 $X2=0
+ $Y2=0
cc_699 N_A_1569_126#_c_781_n N_VPWR_c_1949_n 0.0171301f $X=8.83 $Y=3.185 $X2=0
+ $Y2=0
cc_700 N_A_1569_126#_c_786_n N_VPWR_c_1949_n 0.0156697f $X=14.185 $Y=2.39 $X2=0
+ $Y2=0
cc_701 N_A_1569_126#_c_787_n N_VPWR_c_1949_n 0.00290267f $X=8.07 $Y=2.39 $X2=0
+ $Y2=0
cc_702 N_A_1569_126#_c_761_n N_A_339_655#_c_2082_n 0.0119116f $X=8.027 $Y=2.225
+ $X2=0 $Y2=0
cc_703 N_A_1569_126#_c_781_n N_A_339_655#_c_2104_n 0.00251646f $X=8.83 $Y=3.185
+ $X2=0 $Y2=0
cc_704 N_A_1569_126#_c_761_n N_A_339_655#_c_2104_n 0.0128081f $X=8.027 $Y=2.225
+ $X2=0 $Y2=0
cc_705 N_A_1569_126#_c_787_n N_A_339_655#_c_2104_n 0.0590207f $X=8.07 $Y=2.39
+ $X2=0 $Y2=0
cc_706 N_A_1569_126#_c_781_n N_A_339_655#_c_2105_n 3.35152e-19 $X=8.83 $Y=3.185
+ $X2=0 $Y2=0
cc_707 N_A_1569_126#_c_787_n N_A_339_655#_c_2105_n 0.0219463f $X=8.07 $Y=2.39
+ $X2=0 $Y2=0
cc_708 N_A_1569_126#_c_781_n N_A_339_655#_c_2109_n 0.0221467f $X=8.83 $Y=3.185
+ $X2=0 $Y2=0
cc_709 N_A_1569_126#_c_781_n N_A_339_655#_c_2084_n 0.0331461f $X=8.83 $Y=3.185
+ $X2=0 $Y2=0
cc_710 N_A_1569_126#_c_761_n N_A_339_655#_c_2084_n 0.0320403f $X=8.027 $Y=2.225
+ $X2=0 $Y2=0
cc_711 N_A_1569_126#_c_787_n N_A_339_655#_c_2084_n 0.064118f $X=8.07 $Y=2.39
+ $X2=0 $Y2=0
cc_712 N_A_1569_126#_c_781_n N_A_339_655#_c_2112_n 0.0200951f $X=8.83 $Y=3.185
+ $X2=0 $Y2=0
cc_713 N_A_1569_126#_c_787_n N_A_339_655#_c_2112_n 0.0242542f $X=8.07 $Y=2.39
+ $X2=0 $Y2=0
cc_714 N_A_1569_126#_c_760_n N_A_339_655#_c_2086_n 0.0237605f $X=7.985 $Y=0.83
+ $X2=0 $Y2=0
cc_715 N_A_1569_126#_c_762_n N_A_339_655#_c_2086_n 0.0359366f $X=9.7 $Y=0.35
+ $X2=0 $Y2=0
cc_716 N_A_1569_126#_c_767_n N_VGND_M1008_d 0.00590299f $X=11.975 $Y=1.01 $X2=0
+ $Y2=0
cc_717 N_A_1569_126#_c_760_n N_VGND_c_2298_n 0.0242531f $X=7.985 $Y=0.83 $X2=0
+ $Y2=0
cc_718 N_A_1569_126#_c_764_n N_VGND_c_2298_n 0.00489946f $X=8.15 $Y=0.35 $X2=0
+ $Y2=0
cc_719 N_A_1569_126#_c_767_n N_VGND_c_2300_n 0.0594447f $X=11.975 $Y=1.01 $X2=0
+ $Y2=0
cc_720 N_A_1569_126#_c_828_p N_VGND_c_2300_n 0.0155808f $X=12.06 $Y=0.925 $X2=0
+ $Y2=0
cc_721 N_A_1569_126#_c_770_n N_VGND_c_2300_n 0.00502463f $X=12.145 $Y=0.35 $X2=0
+ $Y2=0
cc_722 N_A_1569_126#_c_772_n N_VGND_c_2302_n 0.00465917f $X=14.1 $Y=0.35 $X2=0
+ $Y2=0
cc_723 N_A_1569_126#_c_774_n N_VGND_c_2302_n 0.0311598f $X=14.185 $Y=2.39 $X2=0
+ $Y2=0
cc_724 N_A_1569_126#_c_760_n N_VGND_c_2308_n 0.0221323f $X=7.985 $Y=0.83 $X2=0
+ $Y2=0
cc_725 N_A_1569_126#_c_762_n N_VGND_c_2308_n 0.07018f $X=9.7 $Y=0.35 $X2=0 $Y2=0
cc_726 N_A_1569_126#_c_764_n N_VGND_c_2308_n 0.00921692f $X=8.15 $Y=0.35 $X2=0
+ $Y2=0
cc_727 N_A_1569_126#_c_766_n N_VGND_c_2308_n 0.032529f $X=9.837 $Y=0.925 $X2=0
+ $Y2=0
cc_728 N_A_1569_126#_c_767_n N_VGND_c_2308_n 0.0430075f $X=11.975 $Y=1.01 $X2=0
+ $Y2=0
cc_729 N_A_1569_126#_c_828_p N_VGND_c_2308_n 0.0190071f $X=12.06 $Y=0.925 $X2=0
+ $Y2=0
cc_730 N_A_1569_126#_c_768_n N_VGND_c_2308_n 0.0234961f $X=12.825 $Y=0.35 $X2=0
+ $Y2=0
cc_731 N_A_1569_126#_c_770_n N_VGND_c_2308_n 0.00773045f $X=12.145 $Y=0.35 $X2=0
+ $Y2=0
cc_732 N_A_1569_126#_c_801_p N_VGND_c_2308_n 0.0229942f $X=12.91 $Y=1.475 $X2=0
+ $Y2=0
cc_733 N_A_1569_126#_c_772_n N_VGND_c_2308_n 0.050422f $X=14.1 $Y=0.35 $X2=0
+ $Y2=0
cc_734 N_A_1569_126#_c_774_n N_VGND_c_2308_n 0.021187f $X=14.185 $Y=2.39 $X2=0
+ $Y2=0
cc_735 N_A_1569_126#_c_776_n N_VGND_c_2308_n 0.00355762f $X=12.91 $Y=0.35 $X2=0
+ $Y2=0
cc_736 N_A_1569_126#_M1004_g N_VGND_c_2308_n 0.010862f $X=9.745 $Y=0.84 $X2=0
+ $Y2=0
cc_737 N_A_1569_126#_c_780_n N_VGND_c_2308_n 0.0156595f $X=12.897 $Y=1.395 $X2=0
+ $Y2=0
cc_738 N_A_1569_126#_c_767_n A_1999_126# 6.46584e-19 $X=11.975 $Y=1.01 $X2=0
+ $Y2=0
cc_739 N_A_1569_126#_c_767_n A_2141_126# 9.12575e-19 $X=11.975 $Y=1.01 $X2=0
+ $Y2=0
cc_740 N_A_1569_126#_c_774_n A_2799_107# 0.00627186f $X=14.185 $Y=2.39 $X2=0
+ $Y2=0
cc_741 N_A_1290_126#_c_974_n N_A_2014_537#_c_1170_n 0.028997f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_742 N_A_1290_126#_c_1012_n N_A_2014_537#_c_1170_n 0.00361239f $X=9.675
+ $Y=2.17 $X2=0 $Y2=0
cc_743 N_A_1290_126#_c_979_n N_A_2014_537#_c_1170_n 0.0287404f $X=9.675 $Y=2.17
+ $X2=0 $Y2=0
cc_744 N_A_1290_126#_M1037_g N_A_2014_537#_c_1171_n 0.0826493f $X=9.61 $Y=3.505
+ $X2=0 $Y2=0
cc_745 N_A_1290_126#_c_974_n N_A_2014_537#_c_1171_n 0.00378335f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_746 N_A_1290_126#_c_974_n N_A_2014_537#_c_1163_n 0.00127949f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_747 N_A_1290_126#_c_959_n N_A_2014_537#_c_1164_n 0.015633f $X=12.125 $Y=1.96
+ $X2=0 $Y2=0
cc_748 N_A_1290_126#_c_960_n N_A_2014_537#_c_1164_n 0.00633621f $X=11.595
+ $Y=1.96 $X2=0 $Y2=0
cc_749 N_A_1290_126#_c_1031_p N_A_2014_537#_c_1164_n 0.0049359f $X=12.21 $Y=1.96
+ $X2=0 $Y2=0
cc_750 N_A_1290_126#_c_978_n N_A_2014_537#_c_1166_n 0.0339151f $X=13.055 $Y=2.26
+ $X2=0 $Y2=0
cc_751 N_A_1290_126#_c_964_n N_A_2014_537#_c_1166_n 0.0218358f $X=13.21 $Y=2.16
+ $X2=0 $Y2=0
cc_752 N_A_1290_126#_c_978_n N_A_2014_537#_c_1167_n 0.0101722f $X=13.055 $Y=2.26
+ $X2=0 $Y2=0
cc_753 N_A_1290_126#_c_1031_p N_A_2014_537#_c_1167_n 0.00892504f $X=12.21
+ $Y=1.96 $X2=0 $Y2=0
cc_754 N_A_1290_126#_M1024_g N_A_2014_537#_c_1177_n 0.0294098f $X=13.21 $Y=3.215
+ $X2=0 $Y2=0
cc_755 N_A_1290_126#_M1024_g N_A_2014_537#_c_1180_n 0.0262283f $X=13.21 $Y=3.215
+ $X2=0 $Y2=0
cc_756 N_A_1290_126#_c_978_n N_A_2014_537#_c_1180_n 0.0143734f $X=13.055 $Y=2.26
+ $X2=0 $Y2=0
cc_757 N_A_1290_126#_c_964_n N_A_2014_537#_c_1180_n 0.0127465f $X=13.21 $Y=2.16
+ $X2=0 $Y2=0
cc_758 N_A_1290_126#_M1024_g N_A_2014_537#_c_1181_n 0.00124565f $X=13.21
+ $Y=3.215 $X2=0 $Y2=0
cc_759 N_A_1290_126#_c_978_n N_A_2014_537#_c_1181_n 0.0183425f $X=13.055 $Y=2.26
+ $X2=0 $Y2=0
cc_760 N_A_1290_126#_c_964_n N_A_2014_537#_c_1181_n 0.00403757f $X=13.21 $Y=2.16
+ $X2=0 $Y2=0
cc_761 N_A_1290_126#_c_978_n N_A_2014_537#_c_1194_n 0.0122207f $X=13.055 $Y=2.26
+ $X2=0 $Y2=0
cc_762 N_A_1290_126#_c_964_n N_A_2014_537#_c_1194_n 0.0264059f $X=13.21 $Y=2.16
+ $X2=0 $Y2=0
cc_763 N_A_1290_126#_c_974_n N_A_2014_537#_c_1195_n 0.00592128f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_764 N_A_1290_126#_c_949_n N_RESET_B_c_1286_n 0.0342495f $X=8.965 $Y=1.125
+ $X2=0 $Y2=0
cc_765 N_A_1290_126#_c_955_n N_RESET_B_c_1286_n 0.00282274f $X=6.59 $Y=0.83
+ $X2=0 $Y2=0
cc_766 N_A_1290_126#_c_963_n N_RESET_B_c_1286_n 0.034112f $X=7.637 $Y=1.125
+ $X2=0 $Y2=0
cc_767 N_A_1290_126#_c_974_n N_RESET_B_c_1305_n 0.0018663f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_768 N_A_1290_126#_M1019_g N_RESET_B_c_1308_n 0.0214164f $X=7.68 $Y=2.62 $X2=0
+ $Y2=0
cc_769 N_A_1290_126#_c_948_n N_RESET_B_c_1308_n 0.0144666f $X=8.715 $Y=1.345
+ $X2=0 $Y2=0
cc_770 N_A_1290_126#_c_950_n N_RESET_B_c_1308_n 0.00747799f $X=9.1 $Y=1.985
+ $X2=0 $Y2=0
cc_771 N_A_1290_126#_c_957_n N_RESET_B_c_1308_n 0.0242997f $X=6.59 $Y=3.19 $X2=0
+ $Y2=0
cc_772 N_A_1290_126#_c_958_n N_RESET_B_c_1308_n 0.0102287f $X=7.365 $Y=1.59
+ $X2=0 $Y2=0
cc_773 N_A_1290_126#_c_974_n N_RESET_B_c_1308_n 0.0264053f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_774 N_A_1290_126#_c_1011_n N_RESET_B_c_1308_n 0.00188853f $X=7.53 $Y=1.51
+ $X2=0 $Y2=0
cc_775 N_A_1290_126#_c_1012_n N_RESET_B_c_1308_n 0.0283132f $X=9.675 $Y=2.17
+ $X2=0 $Y2=0
cc_776 N_A_1290_126#_c_979_n N_RESET_B_c_1308_n 0.0152992f $X=9.675 $Y=2.17
+ $X2=0 $Y2=0
cc_777 N_A_1290_126#_c_974_n N_RESET_B_c_1310_n 0.00857117f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_778 N_A_1290_126#_c_975_n N_RESET_B_c_1310_n 0.00622931f $X=11.51 $Y=2.315
+ $X2=0 $Y2=0
cc_779 N_A_1290_126#_c_959_n N_RESET_B_c_1310_n 0.0189341f $X=12.125 $Y=1.96
+ $X2=0 $Y2=0
cc_780 N_A_1290_126#_c_960_n N_RESET_B_c_1310_n 0.00515656f $X=11.595 $Y=1.96
+ $X2=0 $Y2=0
cc_781 N_A_1290_126#_c_978_n N_RESET_B_c_1310_n 0.0265913f $X=13.055 $Y=2.26
+ $X2=0 $Y2=0
cc_782 N_A_1290_126#_c_1031_p N_RESET_B_c_1310_n 0.0175683f $X=12.21 $Y=1.96
+ $X2=0 $Y2=0
cc_783 N_A_1290_126#_c_964_n N_RESET_B_c_1310_n 0.0235204f $X=13.21 $Y=2.16
+ $X2=0 $Y2=0
cc_784 N_A_1290_126#_c_974_n N_RESET_B_c_1311_n 0.00853574f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_785 N_A_1290_126#_c_975_n N_RESET_B_c_1311_n 6.37106e-19 $X=11.51 $Y=2.315
+ $X2=0 $Y2=0
cc_786 N_A_1290_126#_c_960_n N_RESET_B_c_1311_n 2.05628e-19 $X=11.595 $Y=1.96
+ $X2=0 $Y2=0
cc_787 N_A_1290_126#_c_974_n N_RESET_B_M1008_g 0.0289032f $X=11.425 $Y=2.4 $X2=0
+ $Y2=0
cc_788 N_A_1290_126#_c_975_n N_RESET_B_M1008_g 0.00553442f $X=11.51 $Y=2.315
+ $X2=0 $Y2=0
cc_789 N_A_1290_126#_c_960_n N_RESET_B_M1008_g 0.00199016f $X=11.595 $Y=1.96
+ $X2=0 $Y2=0
cc_790 N_A_1290_126#_c_974_n N_RESET_B_c_1293_n 0.0355449f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_791 N_A_1290_126#_c_975_n N_RESET_B_c_1293_n 0.00592676f $X=11.51 $Y=2.315
+ $X2=0 $Y2=0
cc_792 N_A_1290_126#_c_960_n N_RESET_B_c_1293_n 0.0127276f $X=11.595 $Y=1.96
+ $X2=0 $Y2=0
cc_793 N_A_1290_126#_c_975_n N_A_1816_659#_M1039_g 2.93198e-19 $X=11.51 $Y=2.315
+ $X2=0 $Y2=0
cc_794 N_A_1290_126#_c_959_n N_A_1816_659#_M1039_g 0.0190703f $X=12.125 $Y=1.96
+ $X2=0 $Y2=0
cc_795 N_A_1290_126#_c_1031_p N_A_1816_659#_M1039_g 0.0103687f $X=12.21 $Y=1.96
+ $X2=0 $Y2=0
cc_796 N_A_1290_126#_c_964_n N_A_1816_659#_M1039_g 0.00205077f $X=13.21 $Y=2.16
+ $X2=0 $Y2=0
cc_797 N_A_1290_126#_M1024_g N_A_1816_659#_M1003_g 0.0125691f $X=13.21 $Y=3.215
+ $X2=19.92 $Y2=0
cc_798 N_A_1290_126#_c_949_n N_A_1816_659#_c_1500_n 0.00370969f $X=8.965
+ $Y=1.125 $X2=0 $Y2=0
cc_799 N_A_1290_126#_c_950_n N_A_1816_659#_c_1500_n 0.0149831f $X=9.1 $Y=1.985
+ $X2=0 $Y2=0
cc_800 N_A_1290_126#_M1037_g N_A_1816_659#_c_1500_n 0.00865443f $X=9.61 $Y=3.505
+ $X2=0 $Y2=0
cc_801 N_A_1290_126#_c_954_n N_A_1816_659#_c_1500_n 0.0143349f $X=9 $Y=1.345
+ $X2=0 $Y2=0
cc_802 N_A_1290_126#_c_1012_n N_A_1816_659#_c_1500_n 0.0410391f $X=9.675 $Y=2.17
+ $X2=0 $Y2=0
cc_803 N_A_1290_126#_c_979_n N_A_1816_659#_c_1500_n 0.0257266f $X=9.675 $Y=2.17
+ $X2=0 $Y2=0
cc_804 N_A_1290_126#_M1037_g N_A_1816_659#_c_1507_n 0.0176938f $X=9.61 $Y=3.505
+ $X2=0 $Y2=0
cc_805 N_A_1290_126#_M1037_g N_A_1816_659#_c_1510_n 0.0294258f $X=9.61 $Y=3.505
+ $X2=0 $Y2=0
cc_806 N_A_1290_126#_c_974_n N_A_1816_659#_c_1510_n 0.052443f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_807 N_A_1290_126#_c_1012_n N_A_1816_659#_c_1510_n 0.019574f $X=9.675 $Y=2.17
+ $X2=0 $Y2=0
cc_808 N_A_1290_126#_c_974_n N_A_1816_659#_c_1511_n 0.0217277f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_809 N_A_1290_126#_c_959_n N_A_1816_659#_c_1511_n 0.00331029f $X=12.125
+ $Y=1.96 $X2=0 $Y2=0
cc_810 N_A_1290_126#_c_974_n N_A_1816_659#_c_1515_n 0.0131381f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_811 N_A_1290_126#_c_975_n N_A_1816_659#_c_1515_n 0.00612965f $X=11.51
+ $Y=2.315 $X2=0 $Y2=0
cc_812 N_A_1290_126#_c_959_n N_A_1816_659#_c_1515_n 0.0104922f $X=12.125 $Y=1.96
+ $X2=0 $Y2=0
cc_813 N_A_1290_126#_c_1031_p N_A_1816_659#_c_1515_n 0.00776925f $X=12.21
+ $Y=1.96 $X2=0 $Y2=0
cc_814 N_A_1290_126#_c_949_n N_A_1816_659#_c_1501_n 0.00932056f $X=8.965
+ $Y=1.125 $X2=0 $Y2=0
cc_815 N_A_1290_126#_c_954_n N_A_1816_659#_c_1501_n 3.88979e-19 $X=9 $Y=1.345
+ $X2=0 $Y2=0
cc_816 N_A_1290_126#_M1037_g N_A_1816_659#_c_1516_n 0.00324065f $X=9.61 $Y=3.505
+ $X2=0 $Y2=0
cc_817 N_A_1290_126#_c_979_n N_A_1816_659#_c_1516_n 0.00194951f $X=9.675 $Y=2.17
+ $X2=0 $Y2=0
cc_818 N_A_1290_126#_c_974_n N_A_1816_659#_c_1517_n 0.0015681f $X=11.425 $Y=2.4
+ $X2=0 $Y2=0
cc_819 N_A_1290_126#_c_975_n N_A_1816_659#_c_1517_n 0.00241026f $X=11.51
+ $Y=2.315 $X2=0 $Y2=0
cc_820 N_A_1290_126#_c_959_n N_A_1816_659#_c_1517_n 0.00415454f $X=12.125
+ $Y=1.96 $X2=0 $Y2=0
cc_821 N_A_1290_126#_c_978_n N_A_1816_659#_c_1517_n 0.0256665f $X=13.055 $Y=2.26
+ $X2=0 $Y2=0
cc_822 N_A_1290_126#_c_1031_p N_A_1816_659#_c_1517_n 0.0158405f $X=12.21 $Y=1.96
+ $X2=0 $Y2=0
cc_823 N_A_1290_126#_c_964_n N_A_1816_659#_c_1517_n 0.0372373f $X=13.21 $Y=2.16
+ $X2=0 $Y2=0
cc_824 N_A_1290_126#_M1020_g N_A_2841_81#_c_1618_n 0.0376325f $X=13.745 $Y=0.745
+ $X2=0 $Y2=0
cc_825 N_A_1290_126#_c_951_n N_A_2841_81#_c_1620_n 0.0376325f $X=13.727 $Y=1.352
+ $X2=19.92 $Y2=0
cc_826 N_A_1290_126#_c_952_n N_A_2841_81#_c_1624_n 0.00642895f $X=13.727
+ $Y=1.735 $X2=0 $Y2=0
cc_827 N_A_1290_126#_c_964_n N_A_2624_107#_c_1723_n 9.30023e-19 $X=13.21 $Y=2.16
+ $X2=0 $Y2=0
cc_828 N_A_1290_126#_c_951_n N_A_2624_107#_c_1724_n 6.70233e-19 $X=13.727
+ $Y=1.352 $X2=0 $Y2=0
cc_829 N_A_1290_126#_M1020_g N_A_2624_107#_c_1724_n 0.00763432f $X=13.745
+ $Y=0.745 $X2=0 $Y2=0
cc_830 N_A_1290_126#_c_951_n N_A_2624_107#_c_1725_n 0.0317498f $X=13.727
+ $Y=1.352 $X2=0 $Y2=0
cc_831 N_A_1290_126#_c_964_n N_A_2624_107#_c_1725_n 7.61011e-19 $X=13.21 $Y=2.16
+ $X2=0 $Y2=0
cc_832 N_A_1290_126#_M1024_g N_A_2624_107#_c_1736_n 0.0212656f $X=13.21 $Y=3.215
+ $X2=0 $Y2=0
cc_833 N_A_1290_126#_M1024_g N_A_2624_107#_c_1739_n 0.003354f $X=13.21 $Y=3.215
+ $X2=0 $Y2=0
cc_834 N_A_1290_126#_c_951_n N_A_2624_107#_c_1739_n 0.00231926f $X=13.727
+ $Y=1.352 $X2=0 $Y2=0
cc_835 N_A_1290_126#_c_952_n N_A_2624_107#_c_1739_n 0.0159297f $X=13.727
+ $Y=1.735 $X2=0 $Y2=0
cc_836 N_A_1290_126#_c_964_n N_A_2624_107#_c_1739_n 0.0212945f $X=13.21 $Y=2.16
+ $X2=0 $Y2=0
cc_837 N_A_1290_126#_M1024_g N_A_2624_107#_c_1757_n 0.00496761f $X=13.21
+ $Y=3.215 $X2=0 $Y2=0
cc_838 N_A_1290_126#_c_964_n N_A_2624_107#_c_1757_n 0.00221223f $X=13.21 $Y=2.16
+ $X2=0 $Y2=0
cc_839 N_A_1290_126#_M1019_g N_VPWR_c_1931_n 0.00755044f $X=7.68 $Y=2.62 $X2=0
+ $Y2=0
cc_840 N_A_1290_126#_M1037_g N_VPWR_c_1934_n 0.0060057f $X=9.61 $Y=3.505 $X2=0
+ $Y2=0
cc_841 N_A_1290_126#_M1024_g N_VPWR_c_1937_n 3.53617e-19 $X=13.21 $Y=3.215 $X2=0
+ $Y2=0
cc_842 N_A_1290_126#_c_978_n N_VPWR_c_1937_n 0.00603631f $X=13.055 $Y=2.26 $X2=0
+ $Y2=0
cc_843 N_A_1290_126#_c_1031_p N_VPWR_c_1937_n 0.00364476f $X=12.21 $Y=1.96 $X2=0
+ $Y2=0
cc_844 N_A_1290_126#_M1002_d N_VPWR_c_1949_n 0.00479598f $X=6.45 $Y=2.965 $X2=0
+ $Y2=0
cc_845 N_A_1290_126#_M1019_g N_VPWR_c_1949_n 0.00363935f $X=7.68 $Y=2.62 $X2=0
+ $Y2=0
cc_846 N_A_1290_126#_M1037_g N_VPWR_c_1949_n 0.0149876f $X=9.61 $Y=3.505 $X2=0
+ $Y2=0
cc_847 N_A_1290_126#_M1024_g N_VPWR_c_1949_n 0.0270666f $X=13.21 $Y=3.215 $X2=0
+ $Y2=0
cc_848 N_A_1290_126#_c_957_n N_VPWR_c_1949_n 0.0117486f $X=6.59 $Y=3.19 $X2=0
+ $Y2=0
cc_849 N_A_1290_126#_c_957_n N_A_339_655#_c_2159_n 0.00885538f $X=6.59 $Y=3.19
+ $X2=0 $Y2=0
cc_850 N_A_1290_126#_M1002_d N_A_339_655#_c_2096_n 0.00233214f $X=6.45 $Y=2.965
+ $X2=0 $Y2=0
cc_851 N_A_1290_126#_c_957_n N_A_339_655#_c_2096_n 0.0110919f $X=6.59 $Y=3.19
+ $X2=0 $Y2=0
cc_852 N_A_1290_126#_M1019_g N_A_339_655#_c_2101_n 0.00452167f $X=7.68 $Y=2.62
+ $X2=0 $Y2=0
cc_853 N_A_1290_126#_c_957_n N_A_339_655#_c_2101_n 0.10222f $X=6.59 $Y=3.19
+ $X2=0 $Y2=0
cc_854 N_A_1290_126#_M1019_g N_A_339_655#_c_2082_n 0.019087f $X=7.68 $Y=2.62
+ $X2=0 $Y2=0
cc_855 N_A_1290_126#_c_958_n N_A_339_655#_c_2082_n 0.0225571f $X=7.365 $Y=1.59
+ $X2=0 $Y2=0
cc_856 N_A_1290_126#_c_1011_n N_A_339_655#_c_2082_n 0.0219721f $X=7.53 $Y=1.51
+ $X2=0 $Y2=0
cc_857 N_A_1290_126#_c_962_n N_A_339_655#_c_2082_n 0.00251713f $X=7.637 $Y=1.345
+ $X2=0 $Y2=0
cc_858 N_A_1290_126#_c_957_n N_A_339_655#_c_2083_n 0.0130312f $X=6.59 $Y=3.19
+ $X2=0 $Y2=0
cc_859 N_A_1290_126#_c_958_n N_A_339_655#_c_2083_n 0.0128271f $X=7.365 $Y=1.59
+ $X2=0 $Y2=0
cc_860 N_A_1290_126#_M1019_g N_A_339_655#_c_2104_n 0.0464784f $X=7.68 $Y=2.62
+ $X2=0 $Y2=0
cc_861 N_A_1290_126#_M1019_g N_A_339_655#_c_2105_n 0.00849609f $X=7.68 $Y=2.62
+ $X2=0 $Y2=0
cc_862 N_A_1290_126#_c_949_n N_A_339_655#_c_2084_n 0.00715188f $X=8.965 $Y=1.125
+ $X2=0 $Y2=0
cc_863 N_A_1290_126#_c_950_n N_A_339_655#_c_2084_n 0.0142555f $X=9.1 $Y=1.985
+ $X2=0 $Y2=0
cc_864 N_A_1290_126#_M1037_g N_A_339_655#_c_2084_n 2.61951e-19 $X=9.61 $Y=3.505
+ $X2=0 $Y2=0
cc_865 N_A_1290_126#_c_954_n N_A_339_655#_c_2084_n 0.0262507f $X=9 $Y=1.345
+ $X2=0 $Y2=0
cc_866 N_A_1290_126#_c_979_n N_A_339_655#_c_2084_n 0.015674f $X=9.675 $Y=2.17
+ $X2=0 $Y2=0
cc_867 N_A_1290_126#_c_948_n N_A_339_655#_c_2086_n 0.00953385f $X=8.715 $Y=1.345
+ $X2=0 $Y2=0
cc_868 N_A_1290_126#_c_949_n N_A_339_655#_c_2086_n 0.0194403f $X=8.965 $Y=1.125
+ $X2=0 $Y2=0
cc_869 N_A_1290_126#_c_955_n N_VGND_c_2296_n 0.0157653f $X=6.59 $Y=0.83 $X2=0
+ $Y2=0
cc_870 N_A_1290_126#_c_955_n N_VGND_c_2298_n 0.0299386f $X=6.59 $Y=0.83 $X2=0
+ $Y2=0
cc_871 N_A_1290_126#_c_958_n N_VGND_c_2298_n 0.0155369f $X=7.365 $Y=1.59 $X2=0
+ $Y2=0
cc_872 N_A_1290_126#_c_1011_n N_VGND_c_2298_n 0.0121548f $X=7.53 $Y=1.51 $X2=0
+ $Y2=0
cc_873 N_A_1290_126#_c_963_n N_VGND_c_2298_n 0.0323904f $X=7.637 $Y=1.125 $X2=0
+ $Y2=0
cc_874 N_A_1290_126#_M1020_g N_VGND_c_2302_n 2.22192e-19 $X=13.745 $Y=0.745
+ $X2=0 $Y2=0
cc_875 N_A_1290_126#_c_948_n N_VGND_c_2308_n 0.00625325f $X=8.715 $Y=1.345 $X2=0
+ $Y2=0
cc_876 N_A_1290_126#_c_949_n N_VGND_c_2308_n 0.0132569f $X=8.965 $Y=1.125 $X2=0
+ $Y2=0
cc_877 N_A_1290_126#_c_951_n N_VGND_c_2308_n 9.30698e-19 $X=13.727 $Y=1.352
+ $X2=0 $Y2=0
cc_878 N_A_1290_126#_M1020_g N_VGND_c_2308_n 0.0139437f $X=13.745 $Y=0.745 $X2=0
+ $Y2=0
cc_879 N_A_1290_126#_c_955_n N_VGND_c_2308_n 0.0180823f $X=6.59 $Y=0.83 $X2=0
+ $Y2=0
cc_880 N_A_1290_126#_c_963_n N_VGND_c_2308_n 0.00836502f $X=7.637 $Y=1.125 $X2=0
+ $Y2=0
cc_881 N_A_2014_537#_M1005_g N_RESET_B_c_1286_n 0.0354633f $X=10.455 $Y=0.84
+ $X2=0 $Y2=0
cc_882 N_A_2014_537#_c_1171_n N_RESET_B_M1013_g 0.0334589f $X=10.355 $Y=3.185
+ $X2=0 $Y2=0
cc_883 N_A_2014_537#_c_1170_n N_RESET_B_c_1305_n 0.019226f $X=10.355 $Y=2.685
+ $X2=0 $Y2=0
cc_884 N_A_2014_537#_c_1170_n N_RESET_B_c_1308_n 0.00852581f $X=10.355 $Y=2.685
+ $X2=0 $Y2=0
cc_885 N_A_2014_537#_c_1163_n N_RESET_B_c_1308_n 0.00539874f $X=10.455 $Y=1.965
+ $X2=0 $Y2=0
cc_886 N_A_2014_537#_c_1164_n N_RESET_B_c_1308_n 0.00382822f $X=12.315 $Y=1.36
+ $X2=0 $Y2=0
cc_887 N_A_2014_537#_c_1195_n N_RESET_B_c_1308_n 0.00871692f $X=10.39 $Y=1.44
+ $X2=0 $Y2=0
cc_888 N_A_2014_537#_c_1164_n N_RESET_B_c_1310_n 0.0110453f $X=12.315 $Y=1.36
+ $X2=0 $Y2=0
cc_889 N_A_2014_537#_c_1166_n N_RESET_B_c_1310_n 0.0350558f $X=13.4 $Y=1.91
+ $X2=0 $Y2=0
cc_890 N_A_2014_537#_c_1167_n N_RESET_B_c_1310_n 0.0102364f $X=12.645 $Y=1.91
+ $X2=0 $Y2=0
cc_891 N_A_2014_537#_c_1180_n N_RESET_B_c_1310_n 0.00364181f $X=13.4 $Y=2.61
+ $X2=0 $Y2=0
cc_892 N_A_2014_537#_c_1194_n N_RESET_B_c_1310_n 0.0149975f $X=13.485 $Y=2.525
+ $X2=0 $Y2=0
cc_893 N_A_2014_537#_c_1168_n N_RESET_B_c_1310_n 0.00585318f $X=12.48 $Y=1.36
+ $X2=0 $Y2=0
cc_894 N_A_2014_537#_c_1170_n N_RESET_B_c_1311_n 8.12568e-19 $X=10.355 $Y=2.685
+ $X2=0 $Y2=0
cc_895 N_A_2014_537#_c_1163_n N_RESET_B_c_1311_n 0.00173488f $X=10.455 $Y=1.965
+ $X2=0 $Y2=0
cc_896 N_A_2014_537#_c_1164_n N_RESET_B_c_1311_n 0.00189804f $X=12.315 $Y=1.36
+ $X2=0 $Y2=0
cc_897 N_A_2014_537#_c_1195_n N_RESET_B_c_1311_n 6.32988e-19 $X=10.39 $Y=1.44
+ $X2=0 $Y2=0
cc_898 N_A_2014_537#_c_1170_n N_RESET_B_M1008_g 0.0381711f $X=10.355 $Y=2.685
+ $X2=0 $Y2=0
cc_899 N_A_2014_537#_c_1164_n N_RESET_B_M1008_g 0.0276759f $X=12.315 $Y=1.36
+ $X2=0 $Y2=0
cc_900 N_A_2014_537#_c_1195_n N_RESET_B_M1008_g 0.00107695f $X=10.39 $Y=1.44
+ $X2=0 $Y2=0
cc_901 N_A_2014_537#_M1005_g N_RESET_B_M1008_g 0.10246f $X=10.455 $Y=0.84 $X2=0
+ $Y2=0
cc_902 N_A_2014_537#_c_1170_n N_RESET_B_c_1293_n 0.0040769f $X=10.355 $Y=2.685
+ $X2=0 $Y2=0
cc_903 N_A_2014_537#_c_1163_n N_RESET_B_c_1293_n 0.00677744f $X=10.455 $Y=1.965
+ $X2=0 $Y2=0
cc_904 N_A_2014_537#_c_1164_n N_RESET_B_c_1293_n 0.0397385f $X=12.315 $Y=1.36
+ $X2=0 $Y2=0
cc_905 N_A_2014_537#_c_1195_n N_RESET_B_c_1293_n 0.0231936f $X=10.39 $Y=1.44
+ $X2=0 $Y2=0
cc_906 N_A_2014_537#_M1005_g N_RESET_B_c_1293_n 0.00253678f $X=10.455 $Y=0.84
+ $X2=0 $Y2=0
cc_907 N_A_2014_537#_c_1164_n N_A_1816_659#_M1039_g 0.0325973f $X=12.315 $Y=1.36
+ $X2=0 $Y2=0
cc_908 N_A_2014_537#_c_1183_n N_A_1816_659#_M1039_g 0.0171279f $X=12.48 $Y=0.7
+ $X2=0 $Y2=0
cc_909 N_A_2014_537#_c_1165_n N_A_1816_659#_M1039_g 0.00933276f $X=12.56
+ $Y=1.825 $X2=0 $Y2=0
cc_910 N_A_2014_537#_c_1167_n N_A_1816_659#_M1039_g 0.00537403f $X=12.645
+ $Y=1.91 $X2=0 $Y2=0
cc_911 N_A_2014_537#_c_1168_n N_A_1816_659#_M1039_g 0.00295014f $X=12.48 $Y=1.36
+ $X2=0 $Y2=0
cc_912 N_A_2014_537#_c_1177_n N_A_1816_659#_M1003_g 0.00143963f $X=12.82 $Y=2.84
+ $X2=19.92 $Y2=0
cc_913 N_A_2014_537#_c_1171_n N_A_1816_659#_c_1507_n 0.00100653f $X=10.355
+ $Y=3.185 $X2=0 $Y2=0
cc_914 N_A_2014_537#_c_1171_n N_A_1816_659#_c_1510_n 0.0316858f $X=10.355
+ $Y=3.185 $X2=0 $Y2=0
cc_915 N_A_2014_537#_c_1170_n N_A_1816_659#_c_1511_n 7.3487e-19 $X=10.355
+ $Y=2.685 $X2=0 $Y2=0
cc_916 N_A_2014_537#_c_1171_n N_A_1816_659#_c_1512_n 3.3538e-19 $X=10.355
+ $Y=3.185 $X2=0 $Y2=0
cc_917 N_A_2014_537#_c_1166_n N_A_1816_659#_c_1517_n 2.25312e-19 $X=13.4 $Y=1.91
+ $X2=0 $Y2=0
cc_918 N_A_2014_537#_c_1167_n N_A_1816_659#_c_1517_n 0.00329357f $X=12.645
+ $Y=1.91 $X2=0 $Y2=0
cc_919 N_A_2014_537#_c_1181_n N_A_1816_659#_c_1517_n 0.00554711f $X=12.985
+ $Y=2.61 $X2=0 $Y2=0
cc_920 N_A_2014_537#_c_1168_n N_A_1816_659#_c_1517_n 0.00297302f $X=12.48
+ $Y=1.36 $X2=0 $Y2=0
cc_921 N_A_2014_537#_c_1166_n N_A_2624_107#_c_1723_n 0.00949277f $X=13.4 $Y=1.91
+ $X2=0 $Y2=0
cc_922 N_A_2014_537#_c_1166_n N_A_2624_107#_c_1725_n 0.00445434f $X=13.4 $Y=1.91
+ $X2=0 $Y2=0
cc_923 N_A_2014_537#_c_1177_n N_A_2624_107#_c_1736_n 0.0191448f $X=12.82 $Y=2.84
+ $X2=0 $Y2=0
cc_924 N_A_2014_537#_c_1166_n N_A_2624_107#_c_1739_n 0.0120328f $X=13.4 $Y=1.91
+ $X2=0 $Y2=0
cc_925 N_A_2014_537#_c_1180_n N_A_2624_107#_c_1739_n 0.0135105f $X=13.4 $Y=2.61
+ $X2=0 $Y2=0
cc_926 N_A_2014_537#_c_1194_n N_A_2624_107#_c_1739_n 0.0357275f $X=13.485
+ $Y=2.525 $X2=0 $Y2=0
cc_927 N_A_2014_537#_c_1177_n N_A_2624_107#_c_1757_n 0.00602838f $X=12.82
+ $Y=2.84 $X2=0 $Y2=0
cc_928 N_A_2014_537#_c_1180_n N_A_2624_107#_c_1757_n 0.00921598f $X=13.4 $Y=2.61
+ $X2=0 $Y2=0
cc_929 N_A_2014_537#_c_1171_n N_VPWR_c_1934_n 0.0392604f $X=10.355 $Y=3.185
+ $X2=0 $Y2=0
cc_930 N_A_2014_537#_c_1177_n N_VPWR_c_1937_n 0.0294728f $X=12.82 $Y=2.84 $X2=0
+ $Y2=0
cc_931 N_A_2014_537#_M1003_d N_VPWR_c_1949_n 0.00221032f $X=12.68 $Y=2.715 $X2=0
+ $Y2=0
cc_932 N_A_2014_537#_c_1171_n N_VPWR_c_1949_n 0.00188276f $X=10.355 $Y=3.185
+ $X2=0 $Y2=0
cc_933 N_A_2014_537#_c_1177_n N_VPWR_c_1949_n 0.0341333f $X=12.82 $Y=2.84 $X2=0
+ $Y2=0
cc_934 N_A_2014_537#_c_1164_n N_VGND_M1008_d 0.00213878f $X=12.315 $Y=1.36 $X2=0
+ $Y2=0
cc_935 N_A_2014_537#_M1005_g N_VGND_c_2300_n 0.00658188f $X=10.455 $Y=0.84 $X2=0
+ $Y2=0
cc_936 N_A_2014_537#_c_1183_n N_VGND_c_2308_n 0.0227545f $X=12.48 $Y=0.7 $X2=0
+ $Y2=0
cc_937 N_A_2014_537#_M1005_g N_VGND_c_2308_n 0.0120578f $X=10.455 $Y=0.84 $X2=0
+ $Y2=0
cc_938 N_RESET_B_c_1310_n N_A_1816_659#_M1039_g 0.00239513f $X=14.975 $Y=2.035
+ $X2=0 $Y2=0
cc_939 N_RESET_B_M1008_g N_A_1816_659#_M1039_g 0.0542007f $X=11.165 $Y=0.84
+ $X2=0 $Y2=0
cc_940 N_RESET_B_c_1293_n N_A_1816_659#_M1039_g 0.00137169f $X=11.08 $Y=1.71
+ $X2=0 $Y2=0
cc_941 N_RESET_B_c_1308_n N_A_1816_659#_c_1500_n 0.0242535f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_942 N_RESET_B_c_1305_n N_A_1816_659#_c_1510_n 0.0284013f $X=11.132 $Y=3.165
+ $X2=0 $Y2=0
cc_943 N_RESET_B_c_1305_n N_A_1816_659#_c_1511_n 0.0193504f $X=11.132 $Y=3.165
+ $X2=0 $Y2=0
cc_944 N_RESET_B_c_1310_n N_A_1816_659#_c_1511_n 0.004466f $X=14.975 $Y=2.035
+ $X2=0 $Y2=0
cc_945 N_RESET_B_M1013_g N_A_1816_659#_c_1512_n 0.0184292f $X=11.1 $Y=3.505
+ $X2=0 $Y2=0
cc_946 N_RESET_B_c_1305_n N_A_1816_659#_c_1512_n 0.00614737f $X=11.132 $Y=3.165
+ $X2=0 $Y2=0
cc_947 N_RESET_B_c_1310_n N_A_1816_659#_c_1515_n 0.00395745f $X=14.975 $Y=2.035
+ $X2=0 $Y2=0
cc_948 N_RESET_B_M1008_g N_A_1816_659#_c_1515_n 0.00331844f $X=11.165 $Y=0.84
+ $X2=0 $Y2=0
cc_949 N_RESET_B_c_1286_n N_A_1816_659#_c_1501_n 0.00142685f $X=10.915 $Y=0.215
+ $X2=0 $Y2=0
cc_950 N_RESET_B_c_1310_n N_A_1816_659#_c_1517_n 0.0174749f $X=14.975 $Y=2.035
+ $X2=0 $Y2=0
cc_951 N_RESET_B_M1008_g N_A_1816_659#_c_1517_n 0.0257179f $X=11.165 $Y=0.84
+ $X2=0 $Y2=0
cc_952 N_RESET_B_M1014_g N_A_2841_81#_c_1618_n 0.0140837f $X=15.24 $Y=0.745
+ $X2=0 $Y2=0
cc_953 RESET_B N_A_2841_81#_c_1620_n 0.00225566f $X=15.515 $Y=1.95 $X2=19.92
+ $Y2=0
cc_954 N_RESET_B_c_1310_n N_A_2841_81#_c_1620_n 0.00356366f $X=14.975 $Y=2.035
+ $X2=19.92 $Y2=0
cc_955 N_RESET_B_M1014_g N_A_2841_81#_c_1620_n 0.031824f $X=15.24 $Y=0.745
+ $X2=19.92 $Y2=0
cc_956 N_RESET_B_c_1289_n N_A_2841_81#_c_1625_n 0.033276f $X=15.24 $Y=1.765
+ $X2=19.92 $Y2=0
cc_957 RESET_B N_A_2841_81#_c_1625_n 0.0475999f $X=15.515 $Y=1.95 $X2=19.92
+ $Y2=0
cc_958 N_RESET_B_c_1310_n N_A_2841_81#_c_1625_n 0.0071781f $X=14.975 $Y=2.035
+ $X2=19.92 $Y2=0
cc_959 N_RESET_B_c_1312_n N_A_2841_81#_c_1625_n 0.00867358f $X=15.12 $Y=2.035
+ $X2=19.92 $Y2=0
cc_960 N_RESET_B_c_1289_n N_A_2841_81#_c_1626_n 0.0367199f $X=15.24 $Y=1.765
+ $X2=0 $Y2=0
cc_961 RESET_B N_A_2841_81#_c_1626_n 8.09846e-19 $X=15.515 $Y=1.95 $X2=0 $Y2=0
cc_962 N_RESET_B_c_1310_n N_A_2841_81#_c_1626_n 0.00558431f $X=14.975 $Y=2.035
+ $X2=0 $Y2=0
cc_963 N_RESET_B_c_1312_n N_A_2841_81#_c_1626_n 0.00267187f $X=15.12 $Y=2.035
+ $X2=0 $Y2=0
cc_964 N_RESET_B_c_1289_n N_A_2841_81#_c_1627_n 0.00569713f $X=15.24 $Y=1.765
+ $X2=0 $Y2=0
cc_965 N_RESET_B_c_1289_n N_A_2841_81#_c_1628_n 0.00449018f $X=15.24 $Y=1.765
+ $X2=0 $Y2=0
cc_966 RESET_B N_A_2841_81#_c_1628_n 0.00646391f $X=15.515 $Y=1.95 $X2=0 $Y2=0
cc_967 N_RESET_B_c_1289_n N_A_2841_81#_c_1629_n 4.10442e-19 $X=15.24 $Y=1.765
+ $X2=0 $Y2=0
cc_968 RESET_B N_A_2841_81#_c_1629_n 0.0103971f $X=15.515 $Y=1.95 $X2=0 $Y2=0
cc_969 N_RESET_B_M1014_g N_A_2841_81#_c_1622_n 0.00131544f $X=15.24 $Y=0.745
+ $X2=0 $Y2=0
cc_970 N_RESET_B_c_1289_n N_A_2841_81#_c_1624_n 0.036622f $X=15.24 $Y=1.765
+ $X2=0 $Y2=0
cc_971 RESET_B N_A_2841_81#_c_1624_n 8.60134e-19 $X=15.515 $Y=1.95 $X2=0 $Y2=0
cc_972 N_RESET_B_c_1310_n N_A_2841_81#_c_1624_n 0.0145783f $X=14.975 $Y=2.035
+ $X2=0 $Y2=0
cc_973 N_RESET_B_c_1312_n N_A_2841_81#_c_1624_n 0.0014283f $X=15.12 $Y=2.035
+ $X2=0 $Y2=0
cc_974 N_RESET_B_c_1301_n N_A_2841_81#_c_1632_n 0.0133211f $X=15.595 $Y=2.605
+ $X2=0 $Y2=0
cc_975 N_RESET_B_M1014_g N_A_2624_107#_c_1714_n 0.0522043f $X=15.24 $Y=0.745
+ $X2=0 $Y2=0
cc_976 N_RESET_B_c_1289_n N_A_2624_107#_M1021_g 0.0346484f $X=15.24 $Y=1.765
+ $X2=0 $Y2=0
cc_977 N_RESET_B_c_1289_n N_A_2624_107#_c_1719_n 0.0661433f $X=15.24 $Y=1.765
+ $X2=0 $Y2=0
cc_978 RESET_B N_A_2624_107#_c_1719_n 0.00969162f $X=15.515 $Y=1.95 $X2=0 $Y2=0
cc_979 N_RESET_B_c_1310_n N_A_2624_107#_c_1739_n 0.0217393f $X=14.975 $Y=2.035
+ $X2=0 $Y2=0
cc_980 RESET_B N_A_2624_107#_c_1726_n 0.0245582f $X=15.515 $Y=1.95 $X2=0 $Y2=0
cc_981 N_RESET_B_c_1310_n N_A_2624_107#_c_1726_n 0.0215882f $X=14.975 $Y=2.035
+ $X2=0 $Y2=0
cc_982 N_RESET_B_c_1312_n N_A_2624_107#_c_1726_n 0.00262536f $X=15.12 $Y=2.035
+ $X2=0 $Y2=0
cc_983 N_RESET_B_M1014_g N_A_2624_107#_c_1726_n 0.00265947f $X=15.24 $Y=0.745
+ $X2=0 $Y2=0
cc_984 RESET_B N_A_2624_107#_c_1727_n 0.0509576f $X=15.515 $Y=1.95 $X2=0 $Y2=0
cc_985 N_RESET_B_M1014_g N_A_2624_107#_c_1727_n 0.026036f $X=15.24 $Y=0.745
+ $X2=0 $Y2=0
cc_986 RESET_B N_A_2624_107#_c_1789_n 0.0184949f $X=15.515 $Y=1.95 $X2=0 $Y2=0
cc_987 N_RESET_B_M1014_g N_A_2624_107#_c_1789_n 0.00109305f $X=15.24 $Y=0.745
+ $X2=0 $Y2=0
cc_988 N_RESET_B_c_1302_n N_VPWR_c_1928_n 0.0317472f $X=5.292 $Y=3.165 $X2=0
+ $Y2=0
cc_989 N_RESET_B_c_1308_n N_VPWR_c_1931_n 0.00480479f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_990 N_RESET_B_M1013_g N_VPWR_c_1934_n 0.0128405f $X=11.1 $Y=3.505 $X2=0 $Y2=0
cc_991 N_RESET_B_M1013_g N_VPWR_c_1937_n 9.36931e-19 $X=11.1 $Y=3.505 $X2=0
+ $Y2=0
cc_992 N_RESET_B_c_1305_n N_VPWR_c_1937_n 5.62532e-19 $X=11.132 $Y=3.165 $X2=0
+ $Y2=0
cc_993 N_RESET_B_c_1301_n N_VPWR_c_1940_n 0.0424823f $X=15.595 $Y=2.605 $X2=0
+ $Y2=0
cc_994 N_RESET_B_c_1289_n N_VPWR_c_1943_n 5.95873e-19 $X=15.24 $Y=1.765 $X2=0
+ $Y2=0
cc_995 N_RESET_B_M1013_g N_VPWR_c_1949_n 0.0126713f $X=11.1 $Y=3.505 $X2=0 $Y2=0
cc_996 N_RESET_B_c_1301_n N_VPWR_c_1949_n 0.00394878f $X=15.595 $Y=2.605 $X2=0
+ $Y2=0
cc_997 N_RESET_B_c_1302_n N_VPWR_c_1949_n 0.00356272f $X=5.292 $Y=3.165 $X2=0
+ $Y2=0
cc_998 N_RESET_B_M1007_g N_A_339_655#_c_2080_n 0.003959f $X=5.42 $Y=0.84 $X2=0
+ $Y2=0
cc_999 N_RESET_B_c_1302_n N_A_339_655#_c_2091_n 0.00544217f $X=5.292 $Y=3.165
+ $X2=0 $Y2=0
cc_1000 N_RESET_B_M1007_g N_A_339_655#_c_2081_n 0.00220713f $X=5.42 $Y=0.84
+ $X2=0 $Y2=0
cc_1001 N_RESET_B_c_1302_n N_A_339_655#_c_2081_n 0.0203647f $X=5.292 $Y=3.165
+ $X2=0 $Y2=0
cc_1002 N_RESET_B_c_1309_n N_A_339_655#_c_2081_n 0.0012103f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_1003 N_RESET_B_c_1296_n N_A_339_655#_c_2081_n 0.030759f $X=5.4 $Y=1.46 $X2=0
+ $Y2=0
cc_1004 N_RESET_B_c_1297_n N_A_339_655#_c_2081_n 0.061214f $X=5.4 $Y=1.46 $X2=0
+ $Y2=0
cc_1005 N_RESET_B_c_1302_n N_A_339_655#_c_2095_n 0.0413937f $X=5.292 $Y=3.165
+ $X2=0 $Y2=0
cc_1006 N_RESET_B_c_1302_n N_A_339_655#_c_2159_n 0.00102421f $X=5.292 $Y=3.165
+ $X2=0 $Y2=0
cc_1007 N_RESET_B_c_1302_n N_A_339_655#_c_2099_n 3.85997e-19 $X=5.292 $Y=3.165
+ $X2=0 $Y2=0
cc_1008 N_RESET_B_c_1308_n N_A_339_655#_c_2101_n 0.0131146f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_1009 N_RESET_B_c_1308_n N_A_339_655#_c_2082_n 0.0229531f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_1010 N_RESET_B_c_1308_n N_A_339_655#_c_2083_n 0.00393752f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_1011 N_RESET_B_c_1308_n N_A_339_655#_c_2104_n 0.0129215f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_1012 N_RESET_B_c_1308_n N_A_339_655#_c_2084_n 0.0203876f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_1013 N_RESET_B_c_1302_n N_A_339_655#_c_2111_n 0.00418128f $X=5.292 $Y=3.165
+ $X2=0 $Y2=0
cc_1014 N_RESET_B_c_1286_n N_A_339_655#_c_2086_n 0.00171682f $X=10.915 $Y=0.215
+ $X2=0 $Y2=0
cc_1015 N_RESET_B_M1007_g N_VGND_c_2296_n 0.0464004f $X=5.42 $Y=0.84 $X2=0 $Y2=0
cc_1016 N_RESET_B_c_1286_n N_VGND_c_2296_n 0.00566423f $X=10.915 $Y=0.215 $X2=0
+ $Y2=0
cc_1017 N_RESET_B_c_1297_n N_VGND_c_2296_n 0.0190524f $X=5.4 $Y=1.46 $X2=0 $Y2=0
cc_1018 N_RESET_B_c_1286_n N_VGND_c_2298_n 0.0119775f $X=10.915 $Y=0.215 $X2=0
+ $Y2=0
cc_1019 N_RESET_B_c_1286_n N_VGND_c_2300_n 0.00108752f $X=10.915 $Y=0.215 $X2=0
+ $Y2=0
cc_1020 N_RESET_B_M1008_g N_VGND_c_2300_n 0.0392863f $X=11.165 $Y=0.84 $X2=0
+ $Y2=0
cc_1021 N_RESET_B_M1014_g N_VGND_c_2302_n 0.0409043f $X=15.24 $Y=0.745 $X2=0
+ $Y2=0
cc_1022 N_RESET_B_M1007_g N_VGND_c_2308_n 0.00966788f $X=5.42 $Y=0.84 $X2=0
+ $Y2=0
cc_1023 N_RESET_B_c_1286_n N_VGND_c_2308_n 0.0461268f $X=10.915 $Y=0.215 $X2=0
+ $Y2=0
cc_1024 N_RESET_B_c_1287_n N_VGND_c_2308_n 0.00222061f $X=5.67 $Y=0.215 $X2=0
+ $Y2=0
cc_1025 N_RESET_B_M1008_g N_VGND_c_2308_n 0.00248335f $X=11.165 $Y=0.84 $X2=0
+ $Y2=0
cc_1026 N_RESET_B_M1014_g N_VGND_c_2308_n 0.00330791f $X=15.24 $Y=0.745 $X2=0
+ $Y2=0
cc_1027 N_RESET_B_c_1296_n N_VGND_c_2308_n 0.00189555f $X=5.4 $Y=1.46 $X2=0
+ $Y2=0
cc_1028 N_RESET_B_c_1287_n N_noxref_25_c_2436_n 0.00746485f $X=5.67 $Y=0.215
+ $X2=0 $Y2=0
cc_1029 N_RESET_B_c_1296_n N_noxref_25_c_2436_n 8.45386e-19 $X=5.4 $Y=1.46 $X2=0
+ $Y2=0
cc_1030 N_A_1816_659#_c_1511_n N_VPWR_M1003_s 0.00251087f $X=11.55 $Y=3.075
+ $X2=0 $Y2=0
cc_1031 N_A_1816_659#_c_1507_n N_VPWR_c_1934_n 0.0111649f $X=9.22 $Y=3.505 $X2=0
+ $Y2=0
cc_1032 N_A_1816_659#_c_1510_n N_VPWR_c_1934_n 0.0662359f $X=11.325 $Y=2.99
+ $X2=0 $Y2=0
cc_1033 N_A_1816_659#_c_1512_n N_VPWR_c_1934_n 0.0124739f $X=11.49 $Y=3.505
+ $X2=0 $Y2=0
cc_1034 N_A_1816_659#_M1003_g N_VPWR_c_1937_n 0.0434267f $X=12.43 $Y=3.215 $X2=0
+ $Y2=0
cc_1035 N_A_1816_659#_c_1511_n N_VPWR_c_1937_n 0.00521298f $X=11.55 $Y=3.075
+ $X2=0 $Y2=0
cc_1036 N_A_1816_659#_c_1512_n N_VPWR_c_1937_n 0.0505877f $X=11.49 $Y=3.505
+ $X2=0 $Y2=0
cc_1037 N_A_1816_659#_c_1517_n N_VPWR_c_1937_n 0.00718846f $X=12.43 $Y=2.335
+ $X2=0 $Y2=0
cc_1038 N_A_1816_659#_M1017_d N_VPWR_c_1949_n 0.00221032f $X=9.08 $Y=3.295 $X2=0
+ $Y2=0
cc_1039 N_A_1816_659#_M1003_g N_VPWR_c_1949_n 0.00922274f $X=12.43 $Y=3.215
+ $X2=0 $Y2=0
cc_1040 N_A_1816_659#_c_1507_n N_VPWR_c_1949_n 0.037537f $X=9.22 $Y=3.505 $X2=0
+ $Y2=0
cc_1041 N_A_1816_659#_c_1510_n N_VPWR_c_1949_n 0.0381711f $X=11.325 $Y=2.99
+ $X2=0 $Y2=0
cc_1042 N_A_1816_659#_c_1511_n N_VPWR_c_1949_n 0.00637516f $X=11.55 $Y=3.075
+ $X2=0 $Y2=0
cc_1043 N_A_1816_659#_c_1512_n N_VPWR_c_1949_n 0.0502612f $X=11.49 $Y=3.505
+ $X2=0 $Y2=0
cc_1044 N_A_1816_659#_c_1507_n N_A_339_655#_c_2109_n 0.00768891f $X=9.22
+ $Y=3.505 $X2=0 $Y2=0
cc_1045 N_A_1816_659#_c_1500_n N_A_339_655#_c_2084_n 0.125363f $X=9.22 $Y=2.905
+ $X2=0 $Y2=0
cc_1046 N_A_1816_659#_c_1507_n N_A_339_655#_c_2084_n 0.0126204f $X=9.22 $Y=3.505
+ $X2=0 $Y2=0
cc_1047 N_A_1816_659#_c_1516_n N_A_339_655#_c_2084_n 0.0131377f $X=9.26 $Y=2.99
+ $X2=0 $Y2=0
cc_1048 N_A_1816_659#_c_1507_n N_A_339_655#_c_2112_n 0.00430337f $X=9.22
+ $Y=3.505 $X2=0 $Y2=0
cc_1049 N_A_1816_659#_c_1501_n N_A_339_655#_c_2086_n 0.0286496f $X=9.355 $Y=0.85
+ $X2=0 $Y2=0
cc_1050 N_A_1816_659#_M1039_g N_VGND_c_2300_n 0.00289672f $X=12.09 $Y=0.91 $X2=0
+ $Y2=0
cc_1051 N_A_1816_659#_M1039_g N_VGND_c_2308_n 0.0132824f $X=12.09 $Y=0.91 $X2=0
+ $Y2=0
cc_1052 N_A_1816_659#_c_1500_n N_VGND_c_2308_n 4.53261e-19 $X=9.22 $Y=2.905
+ $X2=0 $Y2=0
cc_1053 N_A_1816_659#_c_1501_n N_VGND_c_2308_n 0.0183697f $X=9.355 $Y=0.85 $X2=0
+ $Y2=0
cc_1054 N_A_2841_81#_c_1621_n N_A_2624_107#_c_1714_n 0.00567448f $X=16.46
+ $Y=1.835 $X2=0 $Y2=0
cc_1055 N_A_2841_81#_c_1622_n N_A_2624_107#_c_1714_n 0.0105762f $X=16.46
+ $Y=0.705 $X2=0 $Y2=0
cc_1056 N_A_2841_81#_c_1627_n N_A_2624_107#_M1021_g 0.0142654f $X=15.985
+ $Y=2.925 $X2=0 $Y2=0
cc_1057 N_A_2841_81#_c_1628_n N_A_2624_107#_M1021_g 0.0124288f $X=16.065 $Y=2.3
+ $X2=0 $Y2=0
cc_1058 N_A_2841_81#_c_1669_p N_A_2624_107#_M1021_g 0.0156678f $X=16.375 $Y=1.92
+ $X2=0 $Y2=0
cc_1059 N_A_2841_81#_c_1629_n N_A_2624_107#_M1021_g 0.00130737f $X=16.15 $Y=1.92
+ $X2=0 $Y2=0
cc_1060 N_A_2841_81#_c_1630_n N_A_2624_107#_M1021_g 0.00568935f $X=16.025
+ $Y=2.397 $X2=0 $Y2=0
cc_1061 N_A_2841_81#_c_1669_p N_A_2624_107#_M1032_g 4.9062e-19 $X=16.375 $Y=1.92
+ $X2=19.92 $Y2=0
cc_1062 N_A_2841_81#_c_1621_n N_A_2624_107#_c_1716_n 0.00323436f $X=16.46
+ $Y=1.835 $X2=0 $Y2=0
cc_1063 N_A_2841_81#_c_1622_n N_A_2624_107#_c_1716_n 5.99896e-19 $X=16.46
+ $Y=0.705 $X2=0 $Y2=0
cc_1064 N_A_2841_81#_c_1625_n N_A_2624_107#_c_1719_n 0.002228f $X=15.9 $Y=2.397
+ $X2=0 $Y2=0
cc_1065 N_A_2841_81#_c_1669_p N_A_2624_107#_c_1719_n 0.0158086f $X=16.375
+ $Y=1.92 $X2=0 $Y2=0
cc_1066 N_A_2841_81#_c_1629_n N_A_2624_107#_c_1719_n 0.00836545f $X=16.15
+ $Y=1.92 $X2=0 $Y2=0
cc_1067 N_A_2841_81#_c_1621_n N_A_2624_107#_c_1719_n 0.0498892f $X=16.46
+ $Y=1.835 $X2=0 $Y2=0
cc_1068 N_A_2841_81#_c_1630_n N_A_2624_107#_c_1719_n 0.00201974f $X=16.025
+ $Y=2.397 $X2=0 $Y2=0
cc_1069 N_A_2841_81#_c_1622_n N_A_2624_107#_c_1719_n 0.00263887f $X=16.46
+ $Y=0.705 $X2=0 $Y2=0
cc_1070 N_A_2841_81#_c_1620_n N_A_2624_107#_c_1739_n 2.44855e-19 $X=14.492
+ $Y=1.565 $X2=0 $Y2=0
cc_1071 N_A_2841_81#_c_1626_n N_A_2624_107#_c_1739_n 2.66042e-19 $X=14.965
+ $Y=2.39 $X2=0 $Y2=0
cc_1072 N_A_2841_81#_c_1632_n N_A_2624_107#_c_1752_n 0.00609327f $X=14.847
+ $Y=2.605 $X2=0 $Y2=0
cc_1073 N_A_2841_81#_c_1620_n N_A_2624_107#_c_1726_n 0.016627f $X=14.492
+ $Y=1.565 $X2=0 $Y2=0
cc_1074 N_A_2841_81#_c_1625_n N_A_2624_107#_c_1726_n 0.0140393f $X=15.9 $Y=2.397
+ $X2=0 $Y2=0
cc_1075 N_A_2841_81#_c_1626_n N_A_2624_107#_c_1726_n 0.0142687f $X=14.965
+ $Y=2.39 $X2=0 $Y2=0
cc_1076 N_A_2841_81#_c_1624_n N_A_2624_107#_c_1726_n 0.0220446f $X=14.847
+ $Y=2.225 $X2=0 $Y2=0
cc_1077 N_A_2841_81#_c_1632_n N_A_2624_107#_c_1726_n 0.00828918f $X=14.847
+ $Y=2.605 $X2=0 $Y2=0
cc_1078 N_A_2841_81#_c_1620_n N_A_2624_107#_c_1727_n 0.0126524f $X=14.492
+ $Y=1.565 $X2=0 $Y2=0
cc_1079 N_A_2841_81#_c_1620_n N_A_2624_107#_c_1756_n 0.00761268f $X=14.492
+ $Y=1.565 $X2=0 $Y2=0
cc_1080 N_A_2841_81#_c_1625_n N_A_2624_107#_c_1789_n 9.5793e-19 $X=15.9 $Y=2.397
+ $X2=0 $Y2=0
cc_1081 N_A_2841_81#_c_1669_p N_A_2624_107#_c_1789_n 0.00312583f $X=16.375
+ $Y=1.92 $X2=0 $Y2=0
cc_1082 N_A_2841_81#_c_1629_n N_A_2624_107#_c_1789_n 0.0135741f $X=16.15 $Y=1.92
+ $X2=0 $Y2=0
cc_1083 N_A_2841_81#_c_1621_n N_A_2624_107#_c_1789_n 0.0415047f $X=16.46
+ $Y=1.835 $X2=0 $Y2=0
cc_1084 N_A_2841_81#_c_1630_n N_A_2624_107#_c_1789_n 0.00254491f $X=16.025
+ $Y=2.397 $X2=0 $Y2=0
cc_1085 N_A_2841_81#_c_1622_n N_A_2624_107#_c_1789_n 0.00144656f $X=16.46
+ $Y=0.705 $X2=0 $Y2=0
cc_1086 N_A_2841_81#_c_1625_n N_VPWR_c_1940_n 0.0681252f $X=15.9 $Y=2.397 $X2=0
+ $Y2=0
cc_1087 N_A_2841_81#_c_1626_n N_VPWR_c_1940_n 0.00177185f $X=14.965 $Y=2.39
+ $X2=0 $Y2=0
cc_1088 N_A_2841_81#_c_1627_n N_VPWR_c_1940_n 0.0230119f $X=15.985 $Y=2.925
+ $X2=0 $Y2=0
cc_1089 N_A_2841_81#_c_1632_n N_VPWR_c_1940_n 0.0360048f $X=14.847 $Y=2.605
+ $X2=0 $Y2=0
cc_1090 N_A_2841_81#_c_1627_n N_VPWR_c_1943_n 0.0505544f $X=15.985 $Y=2.925
+ $X2=0 $Y2=0
cc_1091 N_A_2841_81#_c_1628_n N_VPWR_c_1943_n 0.00829577f $X=16.065 $Y=2.3 $X2=0
+ $Y2=0
cc_1092 N_A_2841_81#_c_1669_p N_VPWR_c_1943_n 0.0169065f $X=16.375 $Y=1.92 $X2=0
+ $Y2=0
cc_1093 N_A_2841_81#_c_1630_n N_VPWR_c_1943_n 0.0156881f $X=16.025 $Y=2.397
+ $X2=0 $Y2=0
cc_1094 N_A_2841_81#_c_1627_n N_VPWR_c_1949_n 0.012777f $X=15.985 $Y=2.925 $X2=0
+ $Y2=0
cc_1095 N_A_2841_81#_c_1632_n N_VPWR_c_1949_n 0.00739612f $X=14.847 $Y=2.605
+ $X2=0 $Y2=0
cc_1096 N_A_2841_81#_c_1618_n N_VGND_c_2302_n 0.0263601f $X=14.492 $Y=1.065
+ $X2=0 $Y2=0
cc_1097 N_A_2841_81#_c_1620_n N_VGND_c_2302_n 0.00186838f $X=14.492 $Y=1.565
+ $X2=0 $Y2=0
cc_1098 N_A_2841_81#_c_1621_n N_VGND_c_2304_n 0.0324396f $X=16.46 $Y=1.835 $X2=0
+ $Y2=0
cc_1099 N_A_2841_81#_c_1622_n N_VGND_c_2304_n 0.0301255f $X=16.46 $Y=0.705 $X2=0
+ $Y2=0
cc_1100 N_A_2841_81#_c_1618_n N_VGND_c_2308_n 0.010098f $X=14.492 $Y=1.065 $X2=0
+ $Y2=0
cc_1101 N_A_2841_81#_c_1621_n N_VGND_c_2308_n 5.69426e-19 $X=16.46 $Y=1.835
+ $X2=0 $Y2=0
cc_1102 N_A_2841_81#_c_1622_n N_VGND_c_2308_n 0.0259693f $X=16.46 $Y=0.705 $X2=0
+ $Y2=0
cc_1103 N_A_2624_107#_M1036_g N_A_3613_443#_M1022_g 0.0184541f $X=18.58 $Y=2.59
+ $X2=0 $Y2=0
cc_1104 N_A_2624_107#_M1009_g N_A_3613_443#_M1010_g 0.0225052f $X=18.61 $Y=0.915
+ $X2=0 $Y2=0
cc_1105 N_A_2624_107#_c_1716_n N_A_3613_443#_c_1879_n 0.00153377f $X=17.28
+ $Y=1.395 $X2=19.92 $Y2=0
cc_1106 N_A_2624_107#_c_1718_n N_A_3613_443#_c_1879_n 0.0170868f $X=18.33
+ $Y=1.657 $X2=19.92 $Y2=0
cc_1107 N_A_2624_107#_M1009_g N_A_3613_443#_c_1879_n 0.0188557f $X=18.61
+ $Y=0.915 $X2=19.92 $Y2=0
cc_1108 N_A_2624_107#_c_1722_n N_A_3613_443#_c_1879_n 0.0105785f $X=18.595
+ $Y=1.74 $X2=19.92 $Y2=0
cc_1109 N_A_2624_107#_M1032_g N_A_3613_443#_c_1885_n 0.00168144f $X=17.25 $Y=2.8
+ $X2=10.08 $Y2=0
cc_1110 N_A_2624_107#_M1036_g N_A_3613_443#_c_1885_n 0.0226028f $X=18.58 $Y=2.59
+ $X2=10.08 $Y2=0
cc_1111 N_A_2624_107#_c_1722_n N_A_3613_443#_c_1885_n 0.00667964f $X=18.595
+ $Y=1.74 $X2=10.08 $Y2=0
cc_1112 N_A_2624_107#_c_1722_n N_A_3613_443#_c_1880_n 0.0435396f $X=18.595
+ $Y=1.74 $X2=0 $Y2=0
cc_1113 N_A_2624_107#_c_1722_n N_A_3613_443#_c_1881_n 0.0229316f $X=18.595
+ $Y=1.74 $X2=0 $Y2=0
cc_1114 N_A_2624_107#_M1032_g N_A_3613_443#_c_1888_n 2.53022e-19 $X=17.25 $Y=2.8
+ $X2=0 $Y2=0
cc_1115 N_A_2624_107#_c_1718_n N_A_3613_443#_c_1888_n 0.0170156f $X=18.33
+ $Y=1.657 $X2=0 $Y2=0
cc_1116 N_A_2624_107#_c_1722_n N_A_3613_443#_c_1888_n 0.00452785f $X=18.595
+ $Y=1.74 $X2=0 $Y2=0
cc_1117 N_A_2624_107#_M1021_g N_VPWR_c_1940_n 5.28304e-19 $X=16.375 $Y=2.925
+ $X2=0 $Y2=0
cc_1118 N_A_2624_107#_c_1752_n N_VPWR_c_1940_n 0.0136768f $X=14.45 $Y=2.96 $X2=0
+ $Y2=0
cc_1119 N_A_2624_107#_c_1726_n N_VPWR_c_1940_n 0.0144514f $X=14.535 $Y=2.875
+ $X2=0 $Y2=0
cc_1120 N_A_2624_107#_M1021_g N_VPWR_c_1943_n 0.0756188f $X=16.375 $Y=2.925
+ $X2=0 $Y2=0
cc_1121 N_A_2624_107#_M1032_g N_VPWR_c_1943_n 0.0776455f $X=17.25 $Y=2.8 $X2=0
+ $Y2=0
cc_1122 N_A_2624_107#_c_1719_n N_VPWR_c_1943_n 0.00822545f $X=17.53 $Y=1.657
+ $X2=0 $Y2=0
cc_1123 N_A_2624_107#_M1036_g N_VPWR_c_1946_n 0.068332f $X=18.58 $Y=2.59 $X2=0
+ $Y2=0
cc_1124 N_A_2624_107#_c_1722_n N_VPWR_c_1946_n 9.10949e-19 $X=18.595 $Y=1.74
+ $X2=0 $Y2=0
cc_1125 N_A_2624_107#_M1021_g N_VPWR_c_1949_n 0.00645594f $X=16.375 $Y=2.925
+ $X2=0 $Y2=0
cc_1126 N_A_2624_107#_M1032_g N_VPWR_c_1949_n 0.0126141f $X=17.25 $Y=2.8 $X2=0
+ $Y2=0
cc_1127 N_A_2624_107#_M1036_g N_VPWR_c_1949_n 0.00584154f $X=18.58 $Y=2.59 $X2=0
+ $Y2=0
cc_1128 N_A_2624_107#_c_1736_n N_VPWR_c_1949_n 0.0487735f $X=13.6 $Y=3.59 $X2=0
+ $Y2=0
cc_1129 N_A_2624_107#_c_1752_n N_VPWR_c_1949_n 0.0271562f $X=14.45 $Y=2.96 $X2=0
+ $Y2=0
cc_1130 N_A_2624_107#_c_1757_n N_VPWR_c_1949_n 0.00682266f $X=13.6 $Y=2.96 $X2=0
+ $Y2=0
cc_1131 N_A_2624_107#_c_1752_n A_2871_543# 0.00314895f $X=14.45 $Y=2.96 $X2=0
+ $Y2=0
cc_1132 N_A_2624_107#_c_1726_n A_2871_543# 0.00193781f $X=14.535 $Y=2.875 $X2=0
+ $Y2=0
cc_1133 N_A_2624_107#_M1032_g N_Q_N_c_2263_n 0.0456337f $X=17.25 $Y=2.8 $X2=0
+ $Y2=0
cc_1134 N_A_2624_107#_c_1716_n N_Q_N_c_2263_n 0.0273659f $X=17.28 $Y=1.395 $X2=0
+ $Y2=0
cc_1135 N_A_2624_107#_c_1718_n N_Q_N_c_2263_n 0.034292f $X=18.33 $Y=1.657 $X2=0
+ $Y2=0
cc_1136 N_A_2624_107#_c_1719_n N_Q_N_c_2263_n 0.0302798f $X=17.53 $Y=1.657 $X2=0
+ $Y2=0
cc_1137 N_A_2624_107#_M1036_g N_Q_N_c_2263_n 0.00339068f $X=18.58 $Y=2.59 $X2=0
+ $Y2=0
cc_1138 N_A_2624_107#_M1009_g N_Q_N_c_2263_n 0.00440284f $X=18.61 $Y=0.915 $X2=0
+ $Y2=0
cc_1139 N_A_2624_107#_c_1722_n N_Q_N_c_2263_n 0.00261745f $X=18.595 $Y=1.74
+ $X2=0 $Y2=0
cc_1140 N_A_2624_107#_c_1714_n N_VGND_c_2302_n 0.00377624f $X=15.95 $Y=1.065
+ $X2=0 $Y2=0
cc_1141 N_A_2624_107#_c_1727_n N_VGND_c_2302_n 0.0497401f $X=15.865 $Y=1.16
+ $X2=0 $Y2=0
cc_1142 N_A_2624_107#_c_1756_n N_VGND_c_2302_n 0.0127568f $X=14.62 $Y=1.16 $X2=0
+ $Y2=0
cc_1143 N_A_2624_107#_c_1714_n N_VGND_c_2304_n 0.00244361f $X=15.95 $Y=1.065
+ $X2=0 $Y2=0
cc_1144 N_A_2624_107#_c_1716_n N_VGND_c_2304_n 0.0515359f $X=17.28 $Y=1.395
+ $X2=0 $Y2=0
cc_1145 N_A_2624_107#_c_1719_n N_VGND_c_2304_n 0.0109584f $X=17.53 $Y=1.657
+ $X2=0 $Y2=0
cc_1146 N_A_2624_107#_M1009_g N_VGND_c_2306_n 0.0547488f $X=18.61 $Y=0.915 $X2=0
+ $Y2=0
cc_1147 N_A_2624_107#_c_1722_n N_VGND_c_2306_n 0.00900332f $X=18.595 $Y=1.74
+ $X2=0 $Y2=0
cc_1148 N_A_2624_107#_M1028_d N_VGND_c_2308_n 0.00311352f $X=13.12 $Y=0.535
+ $X2=0 $Y2=0
cc_1149 N_A_2624_107#_c_1714_n N_VGND_c_2308_n 0.0184959f $X=15.95 $Y=1.065
+ $X2=0 $Y2=0
cc_1150 N_A_2624_107#_c_1716_n N_VGND_c_2308_n 0.013003f $X=17.28 $Y=1.395 $X2=0
+ $Y2=0
cc_1151 N_A_2624_107#_M1009_g N_VGND_c_2308_n 0.0120664f $X=18.61 $Y=0.915 $X2=0
+ $Y2=0
cc_1152 N_A_2624_107#_c_1724_n N_VGND_c_2308_n 0.0174005f $X=13.26 $Y=0.78 $X2=0
+ $Y2=0
cc_1153 N_A_2624_107#_c_1725_n N_VGND_c_2308_n 0.0156593f $X=13.75 $Y=1.21 $X2=0
+ $Y2=0
cc_1154 N_A_2624_107#_c_1727_n N_VGND_c_2308_n 0.0189547f $X=15.865 $Y=1.16
+ $X2=0 $Y2=0
cc_1155 N_A_2624_107#_c_1756_n N_VGND_c_2308_n 7.31377e-19 $X=14.62 $Y=1.16
+ $X2=0 $Y2=0
cc_1156 N_A_2624_107#_c_1789_n N_VGND_c_2308_n 0.0110291f $X=16.03 $Y=1.23 $X2=0
+ $Y2=0
cc_1157 N_A_3613_443#_M1022_g N_VPWR_c_1946_n 0.0703672f $X=19.475 $Y=2.965
+ $X2=0 $Y2=0
cc_1158 N_A_3613_443#_c_1885_n N_VPWR_c_1946_n 0.0614694f $X=18.19 $Y=2.36 $X2=0
+ $Y2=0
cc_1159 N_A_3613_443#_c_1880_n N_VPWR_c_1946_n 0.0722989f $X=19.355 $Y=1.82
+ $X2=0 $Y2=0
cc_1160 N_A_3613_443#_c_1881_n N_VPWR_c_1946_n 0.00155421f $X=19.355 $Y=1.82
+ $X2=0 $Y2=0
cc_1161 N_A_3613_443#_M1022_g N_VPWR_c_1949_n 0.0130327f $X=19.475 $Y=2.965
+ $X2=0 $Y2=0
cc_1162 N_A_3613_443#_c_1885_n N_VPWR_c_1949_n 0.0141253f $X=18.19 $Y=2.36 $X2=0
+ $Y2=0
cc_1163 N_A_3613_443#_c_1879_n N_Q_N_c_2263_n 0.0740405f $X=18.22 $Y=0.915 $X2=0
+ $Y2=0
cc_1164 N_A_3613_443#_c_1885_n N_Q_N_c_2263_n 0.0781004f $X=18.19 $Y=2.36 $X2=0
+ $Y2=0
cc_1165 N_A_3613_443#_c_1888_n N_Q_N_c_2263_n 0.0250019f $X=18.205 $Y=1.82 $X2=0
+ $Y2=0
cc_1166 N_A_3613_443#_M1022_g Q 0.0359985f $X=19.475 $Y=2.965 $X2=0 $Y2=0
cc_1167 N_A_3613_443#_M1010_g Q 0.0242689f $X=19.485 $Y=1.08 $X2=0 $Y2=0
cc_1168 N_A_3613_443#_c_1880_n Q 0.0250567f $X=19.355 $Y=1.82 $X2=0 $Y2=0
cc_1169 N_A_3613_443#_c_1881_n Q 0.0245002f $X=19.355 $Y=1.82 $X2=0 $Y2=0
cc_1170 N_A_3613_443#_M1010_g N_VGND_c_2306_n 0.0519816f $X=19.485 $Y=1.08 $X2=0
+ $Y2=0
cc_1171 N_A_3613_443#_c_1879_n N_VGND_c_2306_n 0.0602549f $X=18.22 $Y=0.915
+ $X2=0 $Y2=0
cc_1172 N_A_3613_443#_c_1880_n N_VGND_c_2306_n 0.0752622f $X=19.355 $Y=1.82
+ $X2=0 $Y2=0
cc_1173 N_A_3613_443#_c_1881_n N_VGND_c_2306_n 0.00180083f $X=19.355 $Y=1.82
+ $X2=0 $Y2=0
cc_1174 N_A_3613_443#_M1010_g N_VGND_c_2308_n 0.0124498f $X=19.485 $Y=1.08 $X2=0
+ $Y2=0
cc_1175 N_A_3613_443#_c_1879_n N_VGND_c_2308_n 0.015678f $X=18.22 $Y=0.915 $X2=0
+ $Y2=0
cc_1176 N_VPWR_c_1949_n N_A_339_655#_M1006_d 9.02611e-19 $X=19.37 $Y=3.59
+ $X2=-0.33 $Y2=1.885
cc_1177 N_VPWR_c_1925_n N_A_339_655#_c_2087_n 0.0558685f $X=3.33 $Y=3.51
+ $X2=19.92 $Y2=4.07
cc_1178 N_VPWR_c_1949_n N_A_339_655#_c_2087_n 0.0682774f $X=19.37 $Y=3.59
+ $X2=19.92 $Y2=4.07
cc_1179 N_VPWR_c_1925_n N_A_339_655#_c_2088_n 0.00991205f $X=3.33 $Y=3.51 $X2=0
+ $Y2=0
cc_1180 N_VPWR_c_1949_n N_A_339_655#_c_2088_n 0.0362681f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_1181 N_VPWR_c_1928_n N_A_339_655#_c_2091_n 0.0246641f $X=5.81 $Y=3.52
+ $X2=10.08 $Y2=4.07
cc_1182 N_VPWR_c_1949_n N_A_339_655#_c_2091_n 0.0326895f $X=19.37 $Y=3.59
+ $X2=10.08 $Y2=4.07
cc_1183 N_VPWR_M1012_d N_A_339_655#_c_2095_n 0.0100666f $X=5.5 $Y=3.275 $X2=0
+ $Y2=0
cc_1184 N_VPWR_c_1928_n N_A_339_655#_c_2095_n 0.0527425f $X=5.81 $Y=3.52 $X2=0
+ $Y2=0
cc_1185 N_VPWR_c_1949_n N_A_339_655#_c_2095_n 0.0131738f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_1186 N_VPWR_c_1928_n N_A_339_655#_c_2159_n 0.0174253f $X=5.81 $Y=3.52 $X2=0
+ $Y2=0
cc_1187 N_VPWR_c_1949_n N_A_339_655#_c_2159_n 0.0180853f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_1188 N_VPWR_c_1931_n N_A_339_655#_c_2096_n 0.00479486f $X=7.29 $Y=2.37 $X2=0
+ $Y2=0
cc_1189 N_VPWR_c_1949_n N_A_339_655#_c_2096_n 0.0289769f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_1190 N_VPWR_c_1928_n N_A_339_655#_c_2099_n 0.00742195f $X=5.81 $Y=3.52 $X2=0
+ $Y2=0
cc_1191 N_VPWR_c_1949_n N_A_339_655#_c_2099_n 0.00604449f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_1192 N_VPWR_c_1931_n N_A_339_655#_c_2101_n 0.101293f $X=7.29 $Y=2.37 $X2=0
+ $Y2=0
cc_1193 N_VPWR_c_1949_n N_A_339_655#_c_2101_n 0.0194693f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_1194 N_VPWR_c_1931_n N_A_339_655#_c_2082_n 0.0114292f $X=7.29 $Y=2.37 $X2=0
+ $Y2=0
cc_1195 N_VPWR_c_1931_n N_A_339_655#_c_2104_n 0.0452192f $X=7.29 $Y=2.37 $X2=0
+ $Y2=0
cc_1196 N_VPWR_c_1949_n N_A_339_655#_c_2105_n 0.0232787f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_1197 N_VPWR_c_1931_n N_A_339_655#_c_2107_n 0.0138528f $X=7.29 $Y=2.37 $X2=0
+ $Y2=0
cc_1198 N_VPWR_c_1949_n N_A_339_655#_c_2107_n 0.00778471f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_1199 N_VPWR_c_1949_n N_A_339_655#_c_2109_n 0.0134344f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_1200 N_VPWR_c_1949_n N_A_339_655#_c_2111_n 0.00737899f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_1201 N_VPWR_c_1949_n N_A_339_655#_c_2112_n 0.0355362f $X=19.37 $Y=3.59 $X2=0
+ $Y2=0
cc_1202 N_VPWR_c_1925_n A_496_655# 0.00454523f $X=3.33 $Y=3.51 $X2=0 $Y2=3.985
cc_1203 N_VPWR_c_1949_n A_496_655# 6.24922e-19 $X=19.37 $Y=3.59 $X2=0 $Y2=3.985
cc_1204 N_VPWR_c_1949_n A_794_655# 0.00201898f $X=19.37 $Y=3.59 $X2=0 $Y2=3.985
cc_1205 N_VPWR_c_1934_n A_1972_659# 0.00526711f $X=10.71 $Y=3.505 $X2=0
+ $Y2=3.985
cc_1206 N_VPWR_c_1949_n A_1972_659# 7.17924e-19 $X=19.37 $Y=3.59 $X2=0 $Y2=3.985
cc_1207 N_VPWR_c_1943_n N_Q_N_c_2263_n 0.104651f $X=16.86 $Y=2.27 $X2=10.08
+ $Y2=4.07
cc_1208 N_VPWR_c_1949_n N_Q_N_c_2263_n 0.0401825f $X=19.37 $Y=3.59 $X2=10.08
+ $Y2=4.07
cc_1209 N_VPWR_c_1946_n Q 0.0994363f $X=19.085 $Y=2.34 $X2=0 $Y2=0
cc_1210 N_VPWR_c_1949_n Q 0.0443798f $X=19.37 $Y=3.59 $X2=0 $Y2=0
cc_1211 N_A_339_655#_c_2080_n N_VGND_c_2296_n 0.00499024f $X=4.885 $Y=1.01 $X2=0
+ $Y2=0
cc_1212 N_A_339_655#_c_2080_n N_VGND_c_2308_n 0.0313265f $X=4.885 $Y=1.01 $X2=0
+ $Y2=0
cc_1213 N_A_339_655#_c_2084_n N_VGND_c_2308_n 4.53054e-19 $X=8.87 $Y=3.255 $X2=0
+ $Y2=0
cc_1214 N_A_339_655#_c_2085_n N_VGND_c_2308_n 0.0207071f $X=3.44 $Y=0.765 $X2=0
+ $Y2=0
cc_1215 N_A_339_655#_c_2086_n N_VGND_c_2308_n 0.0231953f $X=8.87 $Y=0.805 $X2=0
+ $Y2=0
cc_1216 N_A_339_655#_c_2080_n N_noxref_25_M1035_d 0.00412448f $X=4.885 $Y=1.01
+ $X2=0 $Y2=0
cc_1217 N_A_339_655#_c_2080_n N_noxref_25_c_2432_n 0.017636f $X=4.885 $Y=1.01
+ $X2=0.24 $Y2=0
cc_1218 N_A_339_655#_c_2085_n N_noxref_25_c_2432_n 0.0198708f $X=3.44 $Y=0.765
+ $X2=0.24 $Y2=0
cc_1219 N_A_339_655#_c_2080_n N_noxref_25_c_2436_n 0.0183528f $X=4.885 $Y=1.01
+ $X2=0 $Y2=0
cc_1220 N_A_339_655#_c_2080_n noxref_27 0.00153576f $X=4.885 $Y=1.01 $X2=0 $Y2=0
cc_1221 N_Q_N_c_2263_n N_VGND_c_2304_n 0.0580576f $X=17.67 $Y=0.68 $X2=0 $Y2=0
cc_1222 N_Q_N_c_2263_n N_VGND_c_2308_n 0.0390813f $X=17.67 $Y=0.68 $X2=0 $Y2=0
cc_1223 Q N_VGND_c_2306_n 0.0587777f $X=19.835 $Y=0.84 $X2=0 $Y2=0
cc_1224 Q N_VGND_c_2308_n 0.0147384f $X=19.835 $Y=0.84 $X2=0 $Y2=0
cc_1225 N_VGND_c_2308_n N_noxref_25_M1040_s 0.00254395f $X=19.4 $Y=0.48 $X2=0
+ $Y2=0
cc_1226 N_VGND_c_2308_n N_noxref_25_c_2431_n 0.025079f $X=19.4 $Y=0.48 $X2=0
+ $Y2=0
cc_1227 N_VGND_c_2308_n N_noxref_25_c_2432_n 0.0976472f $X=19.4 $Y=0.48 $X2=0.24
+ $Y2=0
cc_1228 N_VGND_c_2308_n N_noxref_25_c_2434_n 0.00701236f $X=19.4 $Y=0.48 $X2=0
+ $Y2=0
cc_1229 N_VGND_c_2296_n N_noxref_25_c_2436_n 0.0269499f $X=5.39 $Y=0.48 $X2=0
+ $Y2=0
cc_1230 N_VGND_c_2308_n N_noxref_25_c_2436_n 0.0305485f $X=19.4 $Y=0.48 $X2=0
+ $Y2=0
cc_1231 N_VGND_c_2308_n noxref_26 0.00875788f $X=19.4 $Y=0.48 $X2=0 $Y2=0
cc_1232 N_VGND_c_2308_n noxref_27 0.00212309f $X=19.4 $Y=0.48 $X2=0 $Y2=0
cc_1233 N_VGND_c_2300_n A_2141_126# 0.0024688f $X=11.64 $Y=0.66 $X2=0 $Y2=0
cc_1234 N_VGND_c_2308_n A_2799_107# 0.00442064f $X=19.4 $Y=0.48 $X2=0 $Y2=0
cc_1235 N_VGND_c_2308_n A_3098_107# 0.00262085f $X=19.4 $Y=0.48 $X2=0 $Y2=0
