* File: sky130_fd_sc_hvl__lsbufhv2hv_lh_1.spice
* Created: Fri Aug 28 09:36:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__lsbufhv2hv_lh_1.pex.spice"
.subckt sky130_fd_sc_hvl__lsbufhv2hv_lh_1  VNB VPB LOWHVPWR A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* LOWHVPWR	LOWHVPWR
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_M1011_g N_A_626_141#_M1011_s N_VNB_M1011_b NHV L=0.5
+ W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250001 A=0.375 P=2.5 MULT=1
MM1000 N_A_847_1221#_M1000_d N_A_626_141#_M1000_g N_VGND_M1000_s N_VNB_M1011_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 M=1 R=3
+ SA=250000 SB=250002 A=0.75 P=4 MULT=1
MM1006 N_A_935_141#_M1006_d N_A_626_141#_M1006_g N_VGND_M1011_d N_VNB_M1011_b
+ NHV L=0.5 W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1002 N_A_847_1221#_M1000_d N_A_626_141#_M1002_g N_VGND_M1002_s N_VNB_M1011_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001
+ SB=250002 A=0.75 P=4 MULT=1
MM1007 N_A_847_1221#_M1007_d N_A_626_141#_M1007_g N_VGND_M1002_s N_VNB_M1011_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002
+ SB=250001 A=0.75 P=4 MULT=1
MM1013 N_A_847_1221#_M1007_d N_A_626_141#_M1013_g N_VGND_M1013_s N_VNB_M1011_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.3975 PD=1.78 PS=3.53 NRD=0 NRS=0 M=1 R=3
+ SA=250002 SB=250000 A=0.75 P=4 MULT=1
MM1008 N_VGND_M1008_d N_A_935_141#_M1008_g N_A_1353_107#_M1008_s N_VNB_M1011_b
+ NHV L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 M=1 R=3
+ SA=250000 SB=250002 A=0.75 P=4 MULT=1
MM1010 N_VGND_M1010_d N_A_935_141#_M1010_g N_A_1353_107#_M1008_s N_VNB_M1011_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250001
+ SB=250002 A=0.75 P=4 MULT=1
MM1012 N_VGND_M1010_d N_A_935_141#_M1012_g N_A_1353_107#_M1012_s N_VNB_M1011_b
+ NHV L=0.5 W=1.5 AD=0.21 AS=0.21 PD=1.78 PS=1.78 NRD=0 NRS=0 M=1 R=3 SA=250002
+ SB=250001 A=0.75 P=4 MULT=1
MM1015 N_VGND_M1015_d N_A_935_141#_M1015_g N_A_1353_107#_M1012_s N_VNB_M1011_b
+ NHV L=0.5 W=1.5 AD=0.3975 AS=0.21 PD=3.53 PS=1.78 NRD=0 NRS=0 M=1 R=3
+ SA=250002 SB=250000 A=0.75 P=4 MULT=1
MM1004 N_X_M1004_d N_A_1353_107#_M1004_g N_VGND_M1004_s N_VNB_M1011_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5 SA=250000
+ SB=250000 A=0.375 P=2.5 MULT=1
MM1014 N_LOWHVPWR_M1014_d N_A_M1014_g N_A_626_141#_M1014_s N_LOWHVPWR_M1014_b
+ PHV L=0.5 W=0.75 AD=0.105 AS=0.19875 PD=1.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1009 N_A_935_141#_M1009_d N_A_626_141#_M1009_g N_LOWHVPWR_M1014_d
+ N_LOWHVPWR_M1014_b PHV L=0.5 W=0.75 AD=0.19875 AS=0.105 PD=2.03 PS=1.03 NRD=0
+ NRS=0 M=1 R=1.5 SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1003 N_VPWR_M1003_d N_A_847_1221#_M1003_g N_A_1353_107#_M1003_s N_VPB_M1003_b
+ PHV L=1 W=0.42 AD=0.2142 AS=0.2142 PD=1.99 PS=1.99 NRD=14.7643 NRS=14.7643 M=1
+ R=0.42 SA=500000 SB=500000 A=0.42 P=2.84 MULT=1
MM1005 N_VPWR_M1005_d N_A_1353_107#_M1005_g N_A_847_1221#_M1005_s N_VPB_M1003_b
+ PHV L=1 W=0.42 AD=0.125081 AS=0.2142 PD=0.95375 PS=1.99 NRD=110.417
+ NRS=14.7643 M=1 R=0.42 SA=500000 SB=500001 A=0.42 P=2.84 MULT=1
MM1001 N_X_M1001_d N_A_1353_107#_M1001_g N_VPWR_M1005_d N_VPB_M1003_b PHV L=0.5
+ W=1.5 AD=0.3975 AS=0.446719 PD=3.53 PS=3.40625 NRD=0 NRS=0 M=1 R=3 SA=250001
+ SB=250000 A=0.75 P=4 MULT=1
DX16_noxref N_VNB_M1011_b N_VPB_X16_noxref_D1 NWDIODE A=4.9381 P=11
DX17_noxref N_VNB_M1011_b N_LOWHVPWR_M1014_b NWDIODE A=5.681 P=9.54
DX18_noxref N_VNB_M1011_b N_VPB_M1003_b NWDIODE A=14.352 P=15.98
*
.include "sky130_fd_sc_hvl__lsbufhv2hv_lh_1.pxi.spice"
*
.ends
*
*
