* File: sky130_fd_sc_hvl__inv_16.pex.spice
* Created: Wed Sep  2 09:06:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__INV_16%VNB 5 7 11
r66 7 11 0.000530134 $w=1.344e-05 $l=5.7e-08 $layer=MET1_cond $X=6.72 $Y=0.057
+ $X2=6.72 $Y2=0
r67 5 11 0.664286 $w=1.7e-07 $l=2.38e-06 $layer=mcon $count=14 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r68 5 11 0.664286 $w=1.7e-07 $l=2.38e-06 $layer=mcon $count=14 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_16%VPB 4 6 14
r103 10 14 0.664286 $w=1.7e-07 $l=2.38e-06 $layer=mcon $count=14 $X=13.2 $Y=4.07
+ $X2=13.2 $Y2=4.07
r104 9 14 845.519 $w=1.68e-07 $l=1.296e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=13.2 $Y2=4.07
r105 9 10 0.664286 $w=1.7e-07 $l=2.38e-06 $layer=mcon $count=14 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r106 6 10 0.000530134 $w=1.344e-05 $l=5.7e-08 $layer=MET1_cond $X=6.72 $Y=4.013
+ $X2=6.72 $Y2=4.07
r107 4 14 13 $w=1.7e-07 $l=1.32424e-05 $layer=licon1_NTAP_notbjt $count=14 $X=0
+ $Y=3.985 $X2=13.2 $Y2=4.07
r108 4 9 13 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=14 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_16%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34
+ 36 38 41 43 45 48 50 52 55 57 59 62 64 66 69 71 73 76 78 80 83 85 87 90 92 94
+ 97 99 101 104 106 108 111 113 193 198 203 208 213 218 223 224 227 231 232 234
+ 235 238 239 241 242 245 246 248 249 251 254 255 257 258 261 262 264 265 268
+ 269 271
r364 249 251 0.0962407 $w=2.3e-07 $l=1.5e-07 $layer=MET1_cond $X=6.32 $Y=1.665
+ $X2=6.47 $Y2=1.665
r365 223 224 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.39 $Y=1.665
+ $X2=11.39 $Y2=1.665
r366 219 264 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=9.83 $Y=1.665
+ $X2=9.86 $Y2=1.665
r367 218 219 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.83 $Y=1.665
+ $X2=9.83 $Y2=1.665
r368 214 257 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=8.27 $Y=1.665
+ $X2=8.3 $Y2=1.665
r369 213 214 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.27 $Y=1.665
+ $X2=8.27 $Y2=1.665
r370 209 248 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=6.71 $Y=1.665
+ $X2=6.74 $Y2=1.665
r371 208 209 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.71 $Y=1.665
+ $X2=6.71 $Y2=1.665
r372 204 241 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=5.15 $Y=1.665
+ $X2=5.18 $Y2=1.665
r373 203 204 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.15 $Y=1.665
+ $X2=5.15 $Y2=1.665
r374 199 234 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=3.59 $Y=1.665
+ $X2=3.62 $Y2=1.665
r375 198 199 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.59 $Y=1.665
+ $X2=3.59 $Y2=1.665
r376 194 227 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=2.04 $Y=1.665
+ $X2=2.07 $Y2=1.665
r377 193 194 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.04 $Y=1.665
+ $X2=2.04 $Y2=1.665
r378 186 223 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.49
+ $Y=1.73 $X2=11.49 $Y2=1.73
r379 179 218 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.93
+ $Y=1.73 $X2=9.93 $Y2=1.73
r380 172 213 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.37
+ $Y=1.73 $X2=8.37 $Y2=1.73
r381 165 208 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.81
+ $Y=1.73 $X2=6.81 $Y2=1.73
r382 158 203 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.25
+ $Y=1.73 $X2=5.25 $Y2=1.73
r383 151 198 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.69
+ $Y=1.73 $X2=3.69 $Y2=1.73
r384 144 193 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.13
+ $Y=1.73 $X2=2.13 $Y2=1.73
r385 113 271 0.0372131 $w=2.3e-07 $l=5.8e-08 $layer=MET1_cond $X=10.942 $Y=1.665
+ $X2=11 $Y2=1.665
r386 113 268 0.0469141 $w=2.3e-07 $l=5.7e-08 $layer=MET1_cond $X=10.942 $Y=1.665
+ $X2=10.885 $Y2=1.665
r387 113 269 0.0475557 $w=2.3e-07 $l=5.8e-08 $layer=MET1_cond $X=9.917 $Y=1.665
+ $X2=9.975 $Y2=1.665
r388 113 264 0.0365714 $w=2.3e-07 $l=5.7e-08 $layer=MET1_cond $X=9.917 $Y=1.665
+ $X2=9.86 $Y2=1.665
r389 113 265 0.0372131 $w=2.3e-07 $l=5.8e-08 $layer=MET1_cond $X=9.382 $Y=1.665
+ $X2=9.44 $Y2=1.665
r390 113 261 0.0469141 $w=2.3e-07 $l=5.7e-08 $layer=MET1_cond $X=9.382 $Y=1.665
+ $X2=9.325 $Y2=1.665
r391 113 262 0.0475557 $w=2.3e-07 $l=5.8e-08 $layer=MET1_cond $X=8.357 $Y=1.665
+ $X2=8.415 $Y2=1.665
r392 113 257 0.0365714 $w=2.3e-07 $l=5.7e-08 $layer=MET1_cond $X=8.357 $Y=1.665
+ $X2=8.3 $Y2=1.665
r393 113 258 0.0372131 $w=2.3e-07 $l=5.8e-08 $layer=MET1_cond $X=7.822 $Y=1.665
+ $X2=7.88 $Y2=1.665
r394 113 254 0.0469141 $w=2.3e-07 $l=5.7e-08 $layer=MET1_cond $X=7.822 $Y=1.665
+ $X2=7.765 $Y2=1.665
r395 113 255 0.0475557 $w=2.3e-07 $l=5.8e-08 $layer=MET1_cond $X=6.797 $Y=1.665
+ $X2=6.855 $Y2=1.665
r396 113 248 0.0365714 $w=2.3e-07 $l=5.7e-08 $layer=MET1_cond $X=6.797 $Y=1.665
+ $X2=6.74 $Y2=1.665
r397 113 249 0.0372131 $w=2.3e-07 $l=5.8e-08 $layer=MET1_cond $X=6.262 $Y=1.665
+ $X2=6.32 $Y2=1.665
r398 113 245 0.0469141 $w=2.3e-07 $l=5.7e-08 $layer=MET1_cond $X=6.262 $Y=1.665
+ $X2=6.205 $Y2=1.665
r399 113 246 0.0475557 $w=2.3e-07 $l=5.8e-08 $layer=MET1_cond $X=5.237 $Y=1.665
+ $X2=5.295 $Y2=1.665
r400 113 241 0.0365714 $w=2.3e-07 $l=5.7e-08 $layer=MET1_cond $X=5.237 $Y=1.665
+ $X2=5.18 $Y2=1.665
r401 113 242 0.0372131 $w=2.3e-07 $l=5.8e-08 $layer=MET1_cond $X=4.702 $Y=1.665
+ $X2=4.76 $Y2=1.665
r402 113 238 0.0469141 $w=2.3e-07 $l=5.7e-08 $layer=MET1_cond $X=4.702 $Y=1.665
+ $X2=4.645 $Y2=1.665
r403 113 239 0.0475557 $w=2.3e-07 $l=5.8e-08 $layer=MET1_cond $X=3.677 $Y=1.665
+ $X2=3.735 $Y2=1.665
r404 113 234 0.0365714 $w=2.3e-07 $l=5.7e-08 $layer=MET1_cond $X=3.677 $Y=1.665
+ $X2=3.62 $Y2=1.665
r405 113 235 0.0372131 $w=2.3e-07 $l=5.8e-08 $layer=MET1_cond $X=3.142 $Y=1.665
+ $X2=3.2 $Y2=1.665
r406 113 231 0.0469141 $w=2.3e-07 $l=5.7e-08 $layer=MET1_cond $X=3.142 $Y=1.665
+ $X2=3.085 $Y2=1.665
r407 113 232 0.0475557 $w=2.3e-07 $l=5.8e-08 $layer=MET1_cond $X=2.127 $Y=1.665
+ $X2=2.185 $Y2=1.665
r408 113 227 0.0365714 $w=2.3e-07 $l=5.7e-08 $layer=MET1_cond $X=2.127 $Y=1.665
+ $X2=2.07 $Y2=1.665
r409 113 224 0.0789173 $w=2.3e-07 $l=1.23e-07 $layer=MET1_cond $X=11.267
+ $Y=1.665 $X2=11.39 $Y2=1.665
r410 113 271 0.171308 $w=2.3e-07 $l=2.67e-07 $layer=MET1_cond $X=11.267 $Y=1.665
+ $X2=11 $Y2=1.665
r411 113 268 0.438111 $w=1.7e-07 $l=4.55e-07 $layer=MET1_cond $X=10.43 $Y=1.665
+ $X2=10.885 $Y2=1.665
r412 113 269 0.438111 $w=1.7e-07 $l=4.55e-07 $layer=MET1_cond $X=10.43 $Y=1.665
+ $X2=9.975 $Y2=1.665
r413 113 219 0.115489 $w=2.3e-07 $l=1.8e-07 $layer=MET1_cond $X=9.65 $Y=1.665
+ $X2=9.83 $Y2=1.665
r414 113 265 0.134737 $w=2.3e-07 $l=2.1e-07 $layer=MET1_cond $X=9.65 $Y=1.665
+ $X2=9.44 $Y2=1.665
r415 113 261 0.438111 $w=1.7e-07 $l=4.55e-07 $layer=MET1_cond $X=8.87 $Y=1.665
+ $X2=9.325 $Y2=1.665
r416 113 262 0.438111 $w=1.7e-07 $l=4.55e-07 $layer=MET1_cond $X=8.87 $Y=1.665
+ $X2=8.415 $Y2=1.665
r417 113 214 0.115489 $w=2.3e-07 $l=1.8e-07 $layer=MET1_cond $X=8.09 $Y=1.665
+ $X2=8.27 $Y2=1.665
r418 113 258 0.134737 $w=2.3e-07 $l=2.1e-07 $layer=MET1_cond $X=8.09 $Y=1.665
+ $X2=7.88 $Y2=1.665
r419 113 254 0.438111 $w=1.7e-07 $l=4.55e-07 $layer=MET1_cond $X=7.31 $Y=1.665
+ $X2=7.765 $Y2=1.665
r420 113 255 0.438111 $w=1.7e-07 $l=4.55e-07 $layer=MET1_cond $X=7.31 $Y=1.665
+ $X2=6.855 $Y2=1.665
r421 113 209 0.115489 $w=2.3e-07 $l=1.8e-07 $layer=MET1_cond $X=6.53 $Y=1.665
+ $X2=6.71 $Y2=1.665
r422 113 251 0.0384963 $w=2.3e-07 $l=6e-08 $layer=MET1_cond $X=6.53 $Y=1.665
+ $X2=6.47 $Y2=1.665
r423 113 245 0.438111 $w=1.7e-07 $l=4.55e-07 $layer=MET1_cond $X=5.75 $Y=1.665
+ $X2=6.205 $Y2=1.665
r424 113 246 0.438111 $w=1.7e-07 $l=4.55e-07 $layer=MET1_cond $X=5.75 $Y=1.665
+ $X2=5.295 $Y2=1.665
r425 113 204 0.115489 $w=2.3e-07 $l=1.8e-07 $layer=MET1_cond $X=4.97 $Y=1.665
+ $X2=5.15 $Y2=1.665
r426 113 242 0.134737 $w=2.3e-07 $l=2.1e-07 $layer=MET1_cond $X=4.97 $Y=1.665
+ $X2=4.76 $Y2=1.665
r427 113 238 0.438111 $w=1.7e-07 $l=4.55e-07 $layer=MET1_cond $X=4.19 $Y=1.665
+ $X2=4.645 $Y2=1.665
r428 113 239 0.438111 $w=1.7e-07 $l=4.55e-07 $layer=MET1_cond $X=4.19 $Y=1.665
+ $X2=3.735 $Y2=1.665
r429 113 199 0.115489 $w=2.3e-07 $l=1.8e-07 $layer=MET1_cond $X=3.41 $Y=1.665
+ $X2=3.59 $Y2=1.665
r430 113 235 0.134737 $w=2.3e-07 $l=2.1e-07 $layer=MET1_cond $X=3.41 $Y=1.665
+ $X2=3.2 $Y2=1.665
r431 113 231 0.433297 $w=1.7e-07 $l=4.5e-07 $layer=MET1_cond $X=2.635 $Y=1.665
+ $X2=3.085 $Y2=1.665
r432 113 232 0.433297 $w=1.7e-07 $l=4.5e-07 $layer=MET1_cond $X=2.635 $Y=1.665
+ $X2=2.185 $Y2=1.665
r433 113 194 0.152702 $w=2.3e-07 $l=2.38e-07 $layer=MET1_cond $X=1.802 $Y=1.665
+ $X2=2.04 $Y2=1.665
r434 109 111 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=12.38 $Y=2.005
+ $X2=12.38 $Y2=2.965
r435 106 109 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=12.375 $Y=1.785
+ $X2=12.38 $Y2=1.785
r436 106 108 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=12.375 $Y=1.565
+ $X2=12.375 $Y2=1.08
r437 102 106 85.0911 $w=4.39e-07 $l=7.75e-07 $layer=POLY_cond $X=11.6 $Y=1.785
+ $X2=12.375 $Y2=1.785
r438 102 104 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=11.6 $Y=2.005
+ $X2=11.6 $Y2=2.965
r439 99 102 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=11.595 $Y=1.785
+ $X2=11.6 $Y2=1.785
r440 99 186 11.5285 $w=4.39e-07 $l=1.05e-07 $layer=POLY_cond $X=11.595 $Y=1.785
+ $X2=11.49 $Y2=1.785
r441 99 101 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.595 $Y=1.565
+ $X2=11.595 $Y2=1.08
r442 95 186 73.5626 $w=4.39e-07 $l=6.7e-07 $layer=POLY_cond $X=10.82 $Y=1.785
+ $X2=11.49 $Y2=1.785
r443 95 97 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=10.82 $Y=2.005
+ $X2=10.82 $Y2=2.965
r444 92 95 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=10.815 $Y=1.785
+ $X2=10.82 $Y2=1.785
r445 92 94 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=10.815 $Y=1.565
+ $X2=10.815 $Y2=1.08
r446 88 92 85.0911 $w=4.39e-07 $l=7.75e-07 $layer=POLY_cond $X=10.04 $Y=1.785
+ $X2=10.815 $Y2=1.785
r447 88 90 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=10.04 $Y=2.005
+ $X2=10.04 $Y2=2.965
r448 85 88 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=10.035 $Y=1.785
+ $X2=10.04 $Y2=1.785
r449 85 179 11.5285 $w=4.39e-07 $l=1.05e-07 $layer=POLY_cond $X=10.035 $Y=1.785
+ $X2=9.93 $Y2=1.785
r450 85 87 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=10.035 $Y=1.565
+ $X2=10.035 $Y2=1.08
r451 81 179 73.5626 $w=4.39e-07 $l=6.7e-07 $layer=POLY_cond $X=9.26 $Y=1.785
+ $X2=9.93 $Y2=1.785
r452 81 83 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=9.26 $Y=2.005
+ $X2=9.26 $Y2=2.965
r453 78 81 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=9.255 $Y=1.785
+ $X2=9.26 $Y2=1.785
r454 78 80 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.255 $Y=1.565
+ $X2=9.255 $Y2=1.08
r455 74 78 85.0911 $w=4.39e-07 $l=7.75e-07 $layer=POLY_cond $X=8.48 $Y=1.785
+ $X2=9.255 $Y2=1.785
r456 74 76 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=8.48 $Y=2.005
+ $X2=8.48 $Y2=2.965
r457 71 74 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=8.475 $Y=1.785
+ $X2=8.48 $Y2=1.785
r458 71 172 11.5285 $w=4.39e-07 $l=1.05e-07 $layer=POLY_cond $X=8.475 $Y=1.785
+ $X2=8.37 $Y2=1.785
r459 71 73 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=8.475 $Y=1.565
+ $X2=8.475 $Y2=1.08
r460 67 172 73.5626 $w=4.39e-07 $l=6.7e-07 $layer=POLY_cond $X=7.7 $Y=1.785
+ $X2=8.37 $Y2=1.785
r461 67 69 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=7.7 $Y=2.005 $X2=7.7
+ $Y2=2.965
r462 64 67 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=7.695 $Y=1.785
+ $X2=7.7 $Y2=1.785
r463 64 66 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.695 $Y=1.565
+ $X2=7.695 $Y2=1.08
r464 60 64 85.0911 $w=4.39e-07 $l=7.75e-07 $layer=POLY_cond $X=6.92 $Y=1.785
+ $X2=7.695 $Y2=1.785
r465 60 62 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=6.92 $Y=2.005
+ $X2=6.92 $Y2=2.965
r466 57 60 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=6.915 $Y=1.785
+ $X2=6.92 $Y2=1.785
r467 57 165 11.5285 $w=4.39e-07 $l=1.05e-07 $layer=POLY_cond $X=6.915 $Y=1.785
+ $X2=6.81 $Y2=1.785
r468 57 59 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.915 $Y=1.565
+ $X2=6.915 $Y2=1.08
r469 53 165 73.5626 $w=4.39e-07 $l=6.7e-07 $layer=POLY_cond $X=6.14 $Y=1.785
+ $X2=6.81 $Y2=1.785
r470 53 55 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=6.14 $Y=2.005
+ $X2=6.14 $Y2=2.965
r471 50 53 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=6.135 $Y=1.785
+ $X2=6.14 $Y2=1.785
r472 50 52 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=6.135 $Y=1.565
+ $X2=6.135 $Y2=1.08
r473 46 50 85.0911 $w=4.39e-07 $l=7.75e-07 $layer=POLY_cond $X=5.36 $Y=1.785
+ $X2=6.135 $Y2=1.785
r474 46 48 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=5.36 $Y=2.005
+ $X2=5.36 $Y2=2.965
r475 43 46 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=5.355 $Y=1.785
+ $X2=5.36 $Y2=1.785
r476 43 158 11.5285 $w=4.39e-07 $l=1.05e-07 $layer=POLY_cond $X=5.355 $Y=1.785
+ $X2=5.25 $Y2=1.785
r477 43 45 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=5.355 $Y=1.565
+ $X2=5.355 $Y2=1.08
r478 39 158 73.5626 $w=4.39e-07 $l=6.7e-07 $layer=POLY_cond $X=4.58 $Y=1.785
+ $X2=5.25 $Y2=1.785
r479 39 41 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=4.58 $Y=2.005
+ $X2=4.58 $Y2=2.965
r480 36 39 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=4.575 $Y=1.785
+ $X2=4.58 $Y2=1.785
r481 36 38 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=4.575 $Y=1.565
+ $X2=4.575 $Y2=1.08
r482 32 36 85.0911 $w=4.39e-07 $l=7.75e-07 $layer=POLY_cond $X=3.8 $Y=1.785
+ $X2=4.575 $Y2=1.785
r483 32 34 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=3.8 $Y=2.005 $X2=3.8
+ $Y2=2.965
r484 29 32 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=3.795 $Y=1.785
+ $X2=3.8 $Y2=1.785
r485 29 151 11.5285 $w=4.39e-07 $l=1.05e-07 $layer=POLY_cond $X=3.795 $Y=1.785
+ $X2=3.69 $Y2=1.785
r486 29 31 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.795 $Y=1.565
+ $X2=3.795 $Y2=1.08
r487 25 151 73.5626 $w=4.39e-07 $l=6.7e-07 $layer=POLY_cond $X=3.02 $Y=1.785
+ $X2=3.69 $Y2=1.785
r488 25 27 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=3.02 $Y=2.005
+ $X2=3.02 $Y2=2.965
r489 22 25 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=3.015 $Y=1.785
+ $X2=3.02 $Y2=1.785
r490 22 24 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.015 $Y=1.565
+ $X2=3.015 $Y2=1.08
r491 18 22 85.0911 $w=4.39e-07 $l=7.75e-07 $layer=POLY_cond $X=2.24 $Y=1.785
+ $X2=3.015 $Y2=1.785
r492 18 20 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=2.24 $Y=2.005
+ $X2=2.24 $Y2=2.965
r493 15 18 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=2.235 $Y=1.785
+ $X2=2.24 $Y2=1.785
r494 15 144 11.5285 $w=4.39e-07 $l=1.05e-07 $layer=POLY_cond $X=2.235 $Y=1.785
+ $X2=2.13 $Y2=1.785
r495 15 17 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.235 $Y=1.565
+ $X2=2.235 $Y2=1.08
r496 11 144 73.5626 $w=4.39e-07 $l=6.7e-07 $layer=POLY_cond $X=1.46 $Y=1.785
+ $X2=2.13 $Y2=1.785
r497 11 13 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.46 $Y=2.005
+ $X2=1.46 $Y2=2.965
r498 8 11 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=1.455 $Y=1.785
+ $X2=1.46 $Y2=1.785
r499 8 10 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.455 $Y=1.565
+ $X2=1.455 $Y2=1.08
r500 4 8 85.0911 $w=4.39e-07 $l=7.75e-07 $layer=POLY_cond $X=0.68 $Y=1.785
+ $X2=1.455 $Y2=1.785
r501 4 6 102.726 $w=5e-07 $l=9.6e-07 $layer=POLY_cond $X=0.68 $Y=2.005 $X2=0.68
+ $Y2=2.965
r502 1 4 0.548975 $w=4.39e-07 $l=5e-09 $layer=POLY_cond $X=0.675 $Y=1.785
+ $X2=0.68 $Y2=1.785
r503 1 3 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.675 $Y=1.565
+ $X2=0.675 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_16%VPWR 1 2 3 4 5 6 7 8 9 28 31 40 51 62 73 84
+ 95 106 117 121
r159 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.81 $Y=3.56
+ $X2=12.81 $Y2=3.56
r160 117 120 23.3381 $w=6.13e-07 $l=1.2e-06 $layer=LI1_cond $X=12.627 $Y=2.36
+ $X2=12.627 $Y2=3.56
r161 112 121 0.477962 $w=3.7e-07 $l=1.245e-06 $layer=MET1_cond $X=11.565 $Y=3.63
+ $X2=12.81 $Y2=3.63
r162 110 112 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.845 $Y=3.63
+ $X2=11.565 $Y2=3.63
r163 109 114 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=11.205 $Y=3.56
+ $X2=11.205 $Y2=3.59
r164 109 112 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.565 $Y=3.56
+ $X2=11.565 $Y2=3.56
r165 109 110 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.845 $Y=3.56
+ $X2=10.845 $Y2=3.56
r166 106 109 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=11.205 $Y=2.34
+ $X2=11.205 $Y2=3.56
r167 101 110 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=10.005 $Y=3.63
+ $X2=10.845 $Y2=3.63
r168 99 101 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=9.285 $Y=3.63
+ $X2=10.005 $Y2=3.63
r169 98 103 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=9.645 $Y=3.56
+ $X2=9.645 $Y2=3.59
r170 98 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.005 $Y=3.56
+ $X2=10.005 $Y2=3.56
r171 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.285 $Y=3.56
+ $X2=9.285 $Y2=3.56
r172 95 98 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=9.645 $Y=2.34
+ $X2=9.645 $Y2=3.56
r173 90 99 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=8.445 $Y=3.63
+ $X2=9.285 $Y2=3.63
r174 88 90 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.725 $Y=3.63
+ $X2=8.445 $Y2=3.63
r175 87 92 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=8.085 $Y=3.56
+ $X2=8.085 $Y2=3.59
r176 87 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.445 $Y=3.56
+ $X2=8.445 $Y2=3.56
r177 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.725 $Y=3.56
+ $X2=7.725 $Y2=3.56
r178 84 87 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=8.085 $Y=2.34
+ $X2=8.085 $Y2=3.56
r179 79 88 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=6.885 $Y=3.63
+ $X2=7.725 $Y2=3.63
r180 76 81 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=6.525 $Y=3.56
+ $X2=6.525 $Y2=3.59
r181 76 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.885 $Y=3.56
+ $X2=6.885 $Y2=3.56
r182 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.165 $Y=3.56
+ $X2=6.165 $Y2=3.56
r183 73 76 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=6.525 $Y=2.34
+ $X2=6.525 $Y2=3.56
r184 68 77 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=5.325 $Y=3.63
+ $X2=6.165 $Y2=3.63
r185 66 68 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=4.605 $Y=3.63
+ $X2=5.325 $Y2=3.63
r186 65 70 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=4.965 $Y=3.56
+ $X2=4.965 $Y2=3.59
r187 65 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.325 $Y=3.56
+ $X2=5.325 $Y2=3.56
r188 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.605 $Y=3.56
+ $X2=4.605 $Y2=3.56
r189 62 65 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=4.965 $Y=2.34
+ $X2=4.965 $Y2=3.56
r190 57 66 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=3.765 $Y=3.63
+ $X2=4.605 $Y2=3.63
r191 55 57 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.045 $Y=3.63
+ $X2=3.765 $Y2=3.63
r192 54 59 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=3.405 $Y=3.56
+ $X2=3.405 $Y2=3.59
r193 54 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.765 $Y=3.56
+ $X2=3.765 $Y2=3.56
r194 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.045 $Y=3.56
+ $X2=3.045 $Y2=3.56
r195 51 54 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=3.405 $Y=2.34
+ $X2=3.405 $Y2=3.56
r196 46 55 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=2.205 $Y=3.63
+ $X2=3.045 $Y2=3.63
r197 44 46 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.485 $Y=3.63
+ $X2=2.205 $Y2=3.63
r198 43 48 0.411236 $w=8.88e-07 $l=3e-08 $layer=LI1_cond $X=1.845 $Y=3.56
+ $X2=1.845 $Y2=3.59
r199 43 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.205 $Y=3.56
+ $X2=2.205 $Y2=3.56
r200 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.485 $Y=3.56
+ $X2=1.485 $Y2=3.56
r201 40 43 16.7236 $w=8.88e-07 $l=1.22e-06 $layer=LI1_cond $X=1.845 $Y=2.34
+ $X2=1.845 $Y2=3.56
r202 35 44 0.351273 $w=3.7e-07 $l=9.15e-07 $layer=MET1_cond $X=0.57 $Y=3.63
+ $X2=1.485 $Y2=3.63
r203 34 37 0.225675 $w=5.28e-07 $l=1e-08 $layer=LI1_cond $X=0.39 $Y=3.56
+ $X2=0.39 $Y2=3.57
r204 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.57 $Y=3.56
+ $X2=0.57 $Y2=3.56
r205 31 34 27.081 $w=5.28e-07 $l=1.2e-06 $layer=LI1_cond $X=0.39 $Y=2.36
+ $X2=0.39 $Y2=3.56
r206 28 79 0.0633444 $w=3.7e-07 $l=1.65e-07 $layer=MET1_cond $X=6.72 $Y=3.63
+ $X2=6.885 $Y2=3.63
r207 28 77 0.213068 $w=3.7e-07 $l=5.55e-07 $layer=MET1_cond $X=6.72 $Y=3.63
+ $X2=6.165 $Y2=3.63
r208 9 120 300 $w=1.7e-07 $l=1.42328e-06 $layer=licon1_PDIFF $count=2 $X=12.63
+ $Y=2.215 $X2=12.77 $Y2=3.57
r209 9 117 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=12.63
+ $Y=2.215 $X2=12.77 $Y2=2.36
r210 8 114 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=11.07
+ $Y=2.215 $X2=11.21 $Y2=3.59
r211 8 106 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=11.07
+ $Y=2.215 $X2=11.21 $Y2=2.34
r212 7 103 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=9.51
+ $Y=2.215 $X2=9.65 $Y2=3.59
r213 7 95 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=9.51
+ $Y=2.215 $X2=9.65 $Y2=2.34
r214 6 92 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=7.95
+ $Y=2.215 $X2=8.09 $Y2=3.59
r215 6 84 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=7.95
+ $Y=2.215 $X2=8.09 $Y2=2.34
r216 5 81 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=6.39
+ $Y=2.215 $X2=6.53 $Y2=3.59
r217 5 73 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=6.39
+ $Y=2.215 $X2=6.53 $Y2=2.34
r218 4 70 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=4.83
+ $Y=2.215 $X2=4.97 $Y2=3.59
r219 4 62 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.83
+ $Y=2.215 $X2=4.97 $Y2=2.34
r220 3 59 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=3.27
+ $Y=2.215 $X2=3.41 $Y2=3.59
r221 3 51 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=3.27
+ $Y=2.215 $X2=3.41 $Y2=2.34
r222 2 48 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.71
+ $Y=2.215 $X2=1.85 $Y2=3.59
r223 2 40 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.71
+ $Y=2.215 $X2=1.85 $Y2=2.34
r224 1 37 300 $w=1.7e-07 $l=1.41612e-06 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=2.215 $X2=0.29 $Y2=3.57
r225 1 31 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=2.215 $X2=0.29 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 49
+ 66 76 86 96 106 116 126 136 145 146 148 149 151 152 154 155 158 159 161 162
+ 164 165
r202 139 143 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=11.985 $Y=2.34
+ $X2=11.985 $Y2=3.59
r203 136 139 48.1931 $w=3.28e-07 $l=1.38e-06 $layer=LI1_cond $X=11.985 $Y=0.96
+ $X2=11.985 $Y2=2.34
r204 129 133 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=10.425 $Y=2.34
+ $X2=10.425 $Y2=3.59
r205 126 129 48.1931 $w=3.28e-07 $l=1.38e-06 $layer=LI1_cond $X=10.425 $Y=0.96
+ $X2=10.425 $Y2=2.34
r206 119 123 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=8.865 $Y=2.34
+ $X2=8.865 $Y2=3.59
r207 116 119 48.1931 $w=3.28e-07 $l=1.38e-06 $layer=LI1_cond $X=8.865 $Y=0.96
+ $X2=8.865 $Y2=2.34
r208 109 113 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=7.305 $Y=2.34
+ $X2=7.305 $Y2=3.59
r209 106 109 48.1931 $w=3.28e-07 $l=1.38e-06 $layer=LI1_cond $X=7.305 $Y=0.96
+ $X2=7.305 $Y2=2.34
r210 99 103 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=5.745 $Y=2.34
+ $X2=5.745 $Y2=3.59
r211 96 99 48.1931 $w=3.28e-07 $l=1.38e-06 $layer=LI1_cond $X=5.745 $Y=0.96
+ $X2=5.745 $Y2=2.34
r212 89 93 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=4.185 $Y=2.34
+ $X2=4.185 $Y2=3.59
r213 86 89 48.1931 $w=3.28e-07 $l=1.38e-06 $layer=LI1_cond $X=4.185 $Y=0.96
+ $X2=4.185 $Y2=2.34
r214 79 83 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=2.625 $Y=2.34
+ $X2=2.625 $Y2=3.59
r215 76 79 48.1931 $w=3.28e-07 $l=1.38e-06 $layer=LI1_cond $X=2.625 $Y=0.96
+ $X2=2.625 $Y2=2.34
r216 69 73 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=1.065 $Y=2.34
+ $X2=1.065 $Y2=3.59
r217 66 69 48.1931 $w=3.28e-07 $l=1.38e-06 $layer=LI1_cond $X=1.065 $Y=0.96
+ $X2=1.065 $Y2=2.34
r218 49 164 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.99 $Y=2.405
+ $X2=11.845 $Y2=2.405
r219 49 165 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.43 $Y=2.405
+ $X2=10.575 $Y2=2.405
r220 49 161 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.43 $Y=2.405
+ $X2=10.285 $Y2=2.405
r221 49 162 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.87 $Y=2.405
+ $X2=9.015 $Y2=2.405
r222 49 158 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.87 $Y=2.405
+ $X2=8.725 $Y2=2.405
r223 49 159 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.31 $Y=2.405
+ $X2=7.455 $Y2=2.405
r224 49 154 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.31 $Y=2.405
+ $X2=7.165 $Y2=2.405
r225 49 155 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.75 $Y=2.405
+ $X2=5.895 $Y2=2.405
r226 49 151 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.75 $Y=2.405
+ $X2=5.605 $Y2=2.405
r227 49 152 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.19 $Y=2.405
+ $X2=4.335 $Y2=2.405
r228 49 148 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.19 $Y=2.405
+ $X2=4.045 $Y2=2.405
r229 49 149 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.63 $Y=2.405
+ $X2=2.775 $Y2=2.405
r230 49 145 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.63 $Y=2.405
+ $X2=2.485 $Y2=2.405
r231 49 146 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.07 $Y=2.405
+ $X2=1.215 $Y2=2.405
r232 49 164 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=11.21 $Y=2.405
+ $X2=11.845 $Y2=2.405
r233 49 165 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=11.21 $Y=2.405
+ $X2=10.575 $Y2=2.405
r234 49 161 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=9.65 $Y=2.405
+ $X2=10.285 $Y2=2.405
r235 49 162 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=9.65 $Y=2.405
+ $X2=9.015 $Y2=2.405
r236 49 158 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=8.09 $Y=2.405
+ $X2=8.725 $Y2=2.405
r237 49 159 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=8.09 $Y=2.405
+ $X2=7.455 $Y2=2.405
r238 49 154 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=6.53 $Y=2.405
+ $X2=7.165 $Y2=2.405
r239 49 155 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=6.53 $Y=2.405
+ $X2=5.895 $Y2=2.405
r240 49 151 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=4.97 $Y=2.405
+ $X2=5.605 $Y2=2.405
r241 49 152 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=4.97 $Y=2.405
+ $X2=4.335 $Y2=2.405
r242 49 148 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=3.41 $Y=2.405
+ $X2=4.045 $Y2=2.405
r243 49 149 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=3.41 $Y=2.405
+ $X2=2.775 $Y2=2.405
r244 49 145 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=1.85 $Y=2.405
+ $X2=2.485 $Y2=2.405
r245 49 146 0.61143 $w=1.7e-07 $l=6.35e-07 $layer=MET1_cond $X=1.85 $Y=2.405
+ $X2=1.215 $Y2=2.405
r246 49 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.99 $Y=2.405
+ $X2=11.99 $Y2=2.405
r247 49 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.43 $Y=2.405
+ $X2=10.43 $Y2=2.405
r248 49 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.87 $Y=2.405
+ $X2=8.87 $Y2=2.405
r249 49 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.31 $Y=2.405
+ $X2=7.31 $Y2=2.405
r250 49 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.405
+ $X2=5.75 $Y2=2.405
r251 49 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.19 $Y=2.405
+ $X2=4.19 $Y2=2.405
r252 49 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.63 $Y=2.405
+ $X2=2.63 $Y2=2.405
r253 49 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.07 $Y=2.405
+ $X2=1.07 $Y2=2.405
r254 16 143 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=11.85
+ $Y=2.215 $X2=11.99 $Y2=3.59
r255 16 139 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=11.85
+ $Y=2.215 $X2=11.99 $Y2=2.34
r256 15 133 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=10.29
+ $Y=2.215 $X2=10.43 $Y2=3.59
r257 15 129 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=10.29
+ $Y=2.215 $X2=10.43 $Y2=2.34
r258 14 123 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=8.73
+ $Y=2.215 $X2=8.87 $Y2=3.59
r259 14 119 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=8.73
+ $Y=2.215 $X2=8.87 $Y2=2.34
r260 13 113 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=7.17
+ $Y=2.215 $X2=7.31 $Y2=3.59
r261 13 109 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=7.17
+ $Y=2.215 $X2=7.31 $Y2=2.34
r262 12 103 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=5.61
+ $Y=2.215 $X2=5.75 $Y2=3.59
r263 12 99 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=5.61
+ $Y=2.215 $X2=5.75 $Y2=2.34
r264 11 93 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=4.05
+ $Y=2.215 $X2=4.19 $Y2=3.59
r265 11 89 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.05
+ $Y=2.215 $X2=4.19 $Y2=2.34
r266 10 83 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.49
+ $Y=2.215 $X2=2.63 $Y2=3.59
r267 10 79 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.49
+ $Y=2.215 $X2=2.63 $Y2=2.34
r268 9 73 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=0.93
+ $Y=2.215 $X2=1.07 $Y2=3.59
r269 9 69 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.93
+ $Y=2.215 $X2=1.07 $Y2=2.34
r270 8 136 91 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=2 $X=11.845
+ $Y=0.705 $X2=11.985 $Y2=0.96
r271 7 126 91 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=2 $X=10.285
+ $Y=0.705 $X2=10.425 $Y2=0.96
r272 6 116 91 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=2 $X=8.725
+ $Y=0.705 $X2=8.865 $Y2=0.96
r273 5 106 91 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=2 $X=7.165
+ $Y=0.705 $X2=7.305 $Y2=0.96
r274 4 96 91 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=2 $X=5.605
+ $Y=0.705 $X2=5.745 $Y2=0.96
r275 3 86 91 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=2 $X=4.045
+ $Y=0.705 $X2=4.185 $Y2=0.96
r276 2 76 91 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=2 $X=2.485
+ $Y=0.705 $X2=2.625 $Y2=0.96
r277 1 66 91 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=2 $X=0.925
+ $Y=0.705 $X2=1.065 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_16%VGND 1 2 3 4 5 6 7 8 9 28 31 38 47 56 65 74
+ 83 92 101 102
r124 101 105 8.46007 $w=6.13e-07 $l=4.35e-07 $layer=LI1_cond $X=12.627 $Y=0.51
+ $X2=12.627 $Y2=0.945
r125 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.81 $Y=0.51
+ $X2=12.81 $Y2=0.51
r126 96 102 0.477962 $w=3.7e-07 $l=1.245e-06 $layer=MET1_cond $X=11.565 $Y=0.44
+ $X2=12.81 $Y2=0.44
r127 93 96 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.845 $Y=0.44
+ $X2=11.565 $Y2=0.44
r128 92 98 5.96292 $w=8.88e-07 $l=4.35e-07 $layer=LI1_cond $X=11.205 $Y=0.51
+ $X2=11.205 $Y2=0.945
r129 92 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.565 $Y=0.51
+ $X2=11.565 $Y2=0.51
r130 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.845 $Y=0.51
+ $X2=10.845 $Y2=0.51
r131 87 93 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=10.005 $Y=0.44
+ $X2=10.845 $Y2=0.44
r132 84 87 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=9.285 $Y=0.44
+ $X2=10.005 $Y2=0.44
r133 83 89 5.96292 $w=8.88e-07 $l=4.35e-07 $layer=LI1_cond $X=9.645 $Y=0.51
+ $X2=9.645 $Y2=0.945
r134 83 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.005 $Y=0.51
+ $X2=10.005 $Y2=0.51
r135 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.285 $Y=0.51
+ $X2=9.285 $Y2=0.51
r136 78 84 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=8.445 $Y=0.44
+ $X2=9.285 $Y2=0.44
r137 75 78 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=7.725 $Y=0.44
+ $X2=8.445 $Y2=0.44
r138 74 80 5.96292 $w=8.88e-07 $l=4.35e-07 $layer=LI1_cond $X=8.085 $Y=0.51
+ $X2=8.085 $Y2=0.945
r139 74 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.445 $Y=0.51
+ $X2=8.445 $Y2=0.51
r140 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.725 $Y=0.51
+ $X2=7.725 $Y2=0.51
r141 69 75 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=6.885 $Y=0.44
+ $X2=7.725 $Y2=0.44
r142 65 71 5.96292 $w=8.88e-07 $l=4.35e-07 $layer=LI1_cond $X=6.525 $Y=0.51
+ $X2=6.525 $Y2=0.945
r143 65 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.885 $Y=0.51
+ $X2=6.885 $Y2=0.51
r144 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.165 $Y=0.51
+ $X2=6.165 $Y2=0.51
r145 60 66 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=5.325 $Y=0.44
+ $X2=6.165 $Y2=0.44
r146 57 60 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=4.605 $Y=0.44
+ $X2=5.325 $Y2=0.44
r147 56 62 5.96292 $w=8.88e-07 $l=4.35e-07 $layer=LI1_cond $X=4.965 $Y=0.51
+ $X2=4.965 $Y2=0.945
r148 56 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.325 $Y=0.51
+ $X2=5.325 $Y2=0.51
r149 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.605 $Y=0.51
+ $X2=4.605 $Y2=0.51
r150 51 57 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=3.765 $Y=0.44
+ $X2=4.605 $Y2=0.44
r151 48 51 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.045 $Y=0.44
+ $X2=3.765 $Y2=0.44
r152 47 53 5.96292 $w=8.88e-07 $l=4.35e-07 $layer=LI1_cond $X=3.405 $Y=0.51
+ $X2=3.405 $Y2=0.945
r153 47 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.765 $Y=0.51
+ $X2=3.765 $Y2=0.51
r154 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.045 $Y=0.51
+ $X2=3.045 $Y2=0.51
r155 42 48 0.322481 $w=3.7e-07 $l=8.4e-07 $layer=MET1_cond $X=2.205 $Y=0.44
+ $X2=3.045 $Y2=0.44
r156 39 42 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.485 $Y=0.44
+ $X2=2.205 $Y2=0.44
r157 38 44 5.96292 $w=8.88e-07 $l=4.35e-07 $layer=LI1_cond $X=1.845 $Y=0.51
+ $X2=1.845 $Y2=0.945
r158 38 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.205 $Y=0.51
+ $X2=2.205 $Y2=0.51
r159 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.485 $Y=0.51
+ $X2=1.485 $Y2=0.51
r160 32 39 0.362791 $w=3.7e-07 $l=9.45e-07 $layer=MET1_cond $X=0.54 $Y=0.44
+ $X2=1.485 $Y2=0.44
r161 31 35 9.72512 $w=5.33e-07 $l=4.35e-07 $layer=LI1_cond $X=0.362 $Y=0.51
+ $X2=0.362 $Y2=0.945
r162 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.54 $Y=0.51
+ $X2=0.54 $Y2=0.51
r163 28 69 0.0633444 $w=3.7e-07 $l=1.65e-07 $layer=MET1_cond $X=6.72 $Y=0.44
+ $X2=6.885 $Y2=0.44
r164 28 66 0.213068 $w=3.7e-07 $l=5.55e-07 $layer=MET1_cond $X=6.72 $Y=0.44
+ $X2=6.165 $Y2=0.44
r165 9 105 91 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=2 $X=12.625
+ $Y=0.705 $X2=12.765 $Y2=0.945
r166 8 98 91 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=2 $X=11.065
+ $Y=0.705 $X2=11.205 $Y2=0.945
r167 7 89 91 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=2 $X=9.505
+ $Y=0.705 $X2=9.645 $Y2=0.945
r168 6 80 91 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=2 $X=7.945
+ $Y=0.705 $X2=8.085 $Y2=0.945
r169 5 71 91 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=2 $X=6.385
+ $Y=0.705 $X2=6.525 $Y2=0.945
r170 4 62 91 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=2 $X=4.825
+ $Y=0.705 $X2=4.965 $Y2=0.945
r171 3 53 91 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=2 $X=3.265
+ $Y=0.705 $X2=3.405 $Y2=0.945
r172 2 44 91 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=2 $X=1.705
+ $Y=0.705 $X2=1.845 $Y2=0.945
r173 1 35 91 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.705 $X2=0.285 $Y2=0.945
.ends

