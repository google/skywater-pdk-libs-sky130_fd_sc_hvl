* File: sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3.pxi.spice
* Created: Fri Aug 28 09:37:12 2020
* 
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%VNB N_VNB_M1018_b VNB VNB
+ N_VNB_c_10_p N_VNB_c_6_p VNB VNB
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%VNB
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%VPB N_VPB_M1005_b N_VPB_c_333_p
+ VPB N_VPB_c_373_p N_VPB_c_313_p N_VPB_c_335_p VPB
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%VPB
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%LVPWR N_LVPWR_M1006_s
+ N_LVPWR_M1003_s N_LVPWR_M1013_s N_LVPWR_M1026_s N_LVPWR_M1025_s
+ N_LVPWR_M1038_s N_LVPWR_M1031_s N_LVPWR_M1044_s N_LVPWR_M1006_b
+ N_LVPWR_c_453_p N_LVPWR_c_398_n N_LVPWR_c_431_p N_LVPWR_c_399_n
+ N_LVPWR_c_400_n N_LVPWR_c_401_n N_LVPWR_c_402_n N_LVPWR_c_457_p
+ N_LVPWR_c_435_p N_LVPWR_c_403_n N_LVPWR_c_404_n N_LVPWR_c_405_n
+ N_LVPWR_c_463_p N_LVPWR_c_444_p N_LVPWR_c_406_n N_LVPWR_c_471_p
+ N_LVPWR_c_579_p N_LVPWR_c_566_p N_LVPWR_c_464_p LVPWR N_LVPWR_c_396_n LVPWR
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%LVPWR
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%VGND N_VGND_M1000_s
+ N_VGND_M1008_d N_VGND_M1004_d N_VGND_M1047_d N_VGND_M1012_d N_VGND_M1010_d
+ N_VGND_M1040_d N_VGND_M1029_d N_VGND_M1041_d N_VGND_M1002_d N_VGND_M1045_d
+ N_VGND_M1007_d N_VGND_M1018_d N_VGND_M1019_d N_VGND_M1009_d N_VGND_M1033_d
+ N_VGND_M1016_d N_VGND_M1024_d N_VGND_M1046_d N_VGND_M1000_g N_VGND_c_590_n
+ N_VGND_c_591_n N_VGND_c_593_n N_VGND_c_594_n N_VGND_c_595_n N_VGND_c_597_n
+ N_VGND_c_598_n N_VGND_c_599_n N_VGND_c_600_n N_VGND_c_602_n N_VGND_c_603_n
+ N_VGND_c_604_n N_VGND_c_605_n N_VGND_c_606_n N_VGND_c_607_n N_VGND_c_608_n
+ N_VGND_c_609_n N_VGND_c_610_n N_VGND_c_612_n N_VGND_c_613_n N_VGND_c_615_n
+ N_VGND_c_616_n N_VGND_c_618_n N_VGND_c_620_n N_VGND_c_621_n N_VGND_c_622_n
+ N_VGND_c_624_n N_VGND_c_626_n N_VGND_c_628_n N_VGND_c_629_n N_VGND_c_630_n
+ N_VGND_c_632_n N_VGND_c_633_n N_VGND_c_635_n N_VGND_c_637_n N_VGND_c_638_n
+ N_VGND_c_639_n N_VGND_c_640_n N_VGND_c_642_n N_VGND_c_644_n N_VGND_c_646_n
+ N_VGND_c_648_n N_VGND_c_650_n N_VGND_c_652_n N_VGND_c_654_n N_VGND_c_656_n
+ N_VGND_c_658_n N_VGND_c_660_n N_VGND_c_662_n N_VGND_c_664_n N_VGND_c_666_n
+ N_VGND_c_668_n N_VGND_c_670_n N_VGND_c_672_n VGND VGND N_VGND_c_674_n
+ N_VGND_c_676_n N_VGND_c_678_n N_VGND_c_680_n N_VGND_c_682_n VGND VGND
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%VGND
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_262_107# N_A_262_107#_M1012_s
+ N_A_262_107#_M1034_s N_A_262_107#_M39_noxref_s N_A_262_107#_M40_noxref_d
+ N_A_262_107#_M1008_g N_A_262_107#_M1005_g N_A_262_107#_c_842_n
+ N_A_262_107#_M1030_g N_A_262_107#_M1011_g N_A_262_107#_c_845_n
+ N_A_262_107#_M1047_g N_A_262_107#_M1036_g N_A_262_107#_c_848_n
+ N_A_262_107#_c_849_n N_A_262_107#_c_850_n N_A_262_107#_c_851_n
+ N_A_262_107#_c_852_n N_A_262_107#_c_868_n N_A_262_107#_c_853_n
+ N_A_262_107#_c_854_n N_A_262_107#_c_871_n N_A_262_107#_c_855_n
+ N_A_262_107#_c_874_n PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_262_107#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_840_107# N_A_840_107#_M1001_s
+ N_A_840_107#_M1032_s N_A_840_107#_M1002_s N_A_840_107#_M1043_d
+ N_A_840_107#_M1012_g N_A_840_107#_M39_noxref_g N_A_840_107#_c_968_n
+ N_A_840_107#_M1034_g N_A_840_107#_M40_noxref_g N_A_840_107#_c_971_n
+ N_A_840_107#_c_988_n N_A_840_107#_c_990_n N_A_840_107#_c_991_n
+ N_A_840_107#_M1022_g N_A_840_107#_c_972_n N_A_840_107#_c_973_n
+ N_A_840_107#_c_996_n N_A_840_107#_c_997_n N_A_840_107#_c_974_n
+ N_A_840_107#_c_975_n N_A_840_107#_c_976_n N_A_840_107#_c_977_n
+ N_A_840_107#_c_978_n N_A_840_107#_c_979_n N_A_840_107#_c_980_n
+ N_A_840_107#_c_1001_n N_A_840_107#_c_1002_n N_A_840_107#_c_1003_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_840_107#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_362_1243#
+ N_A_362_1243#_M1000_d N_A_362_1243#_M1004_s N_A_362_1243#_M1023_s
+ N_A_362_1243#_M1022_s N_A_362_1243#_M1043_g N_A_362_1243#_c_1134_n
+ N_A_362_1243#_c_1123_n N_A_362_1243#_c_1124_n N_A_362_1243#_c_1125_n
+ N_A_362_1243#_c_1126_n N_A_362_1243#_c_1127_n N_A_362_1243#_c_1128_n
+ N_A_362_1243#_c_1129_n N_A_362_1243#_c_1138_n N_A_362_1243#_c_1144_n
+ N_A_362_1243#_c_1139_n N_A_362_1243#_c_1130_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_362_1243#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_2092_381#
+ N_A_2092_381#_M1045_s N_A_2092_381#_M1020_s N_A_2092_381#_M43_noxref_g
+ N_A_2092_381#_c_1220_n N_A_2092_381#_c_1221_n N_A_2092_381#_M44_noxref_g
+ N_A_2092_381#_c_1224_n N_A_2092_381#_M45_noxref_g N_A_2092_381#_c_1227_n
+ N_A_2092_381#_M46_noxref_g N_A_2092_381#_M1002_g N_A_2092_381#_c_1230_n
+ N_A_2092_381#_c_1231_n N_A_2092_381#_c_1232_n N_A_2092_381#_c_1233_n
+ N_A_2092_381#_c_1216_n N_A_2092_381#_c_1235_n N_A_2092_381#_c_1217_n
+ N_A_2092_381#_c_1237_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_2092_381#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_1472_1171#
+ N_A_1472_1171#_M1007_s N_A_1472_1171#_M1014_s N_A_1472_1171#_M1003_d
+ N_A_1472_1171#_M1035_d N_A_1472_1171#_M1001_g N_A_1472_1171#_c_1312_n
+ N_A_1472_1171#_c_1313_n N_A_1472_1171#_M1029_g N_A_1472_1171#_c_1315_n
+ N_A_1472_1171#_c_1316_n N_A_1472_1171#_c_1317_n N_A_1472_1171#_c_1318_n
+ N_A_1472_1171#_M1032_g N_A_1472_1171#_c_1320_n N_A_1472_1171#_M1041_g
+ N_A_1472_1171#_c_1322_n N_A_1472_1171#_c_1323_n N_A_1472_1171#_c_1335_n
+ N_A_1472_1171#_c_1324_n N_A_1472_1171#_c_1325_n N_A_1472_1171#_c_1326_n
+ N_A_1472_1171#_c_1338_n N_A_1472_1171#_c_1339_n N_A_1472_1171#_c_1374_n
+ N_A_1472_1171#_c_1327_n N_A_1472_1171#_c_1344_n N_A_1472_1171#_c_1347_n
+ N_A_1472_1171#_c_1378_n N_A_1472_1171#_c_1328_n N_A_1472_1171#_c_1353_n
+ N_A_1472_1171#_c_1329_n N_A_1472_1171#_c_1330_n N_A_1472_1171#_c_1428_p
+ N_A_1472_1171#_c_1331_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_1472_1171#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%SLEEP_B N_SLEEP_B_M1020_g
+ N_SLEEP_B_M1045_g N_SLEEP_B_c_1468_n SLEEP_B N_SLEEP_B_c_1469_n
+ N_SLEEP_B_c_1470_n PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%SLEEP_B
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_3617_1198#
+ N_A_3617_1198#_M1024_s N_A_3617_1198#_M1031_d N_A_3617_1198#_M1018_g
+ N_A_3617_1198#_c_1508_n N_A_3617_1198#_M1006_g N_A_3617_1198#_M1019_g
+ N_A_3617_1198#_c_1511_n N_A_3617_1198#_M1013_g N_A_3617_1198#_M1027_g
+ N_A_3617_1198#_c_1514_n N_A_3617_1198#_M1015_g N_A_3617_1198#_c_1517_n
+ N_A_3617_1198#_M1025_g N_A_3617_1198#_M1033_g N_A_3617_1198#_c_1500_n
+ N_A_3617_1198#_c_1501_n N_A_3617_1198#_c_1502_n N_A_3617_1198#_c_1503_n
+ N_A_3617_1198#_c_1504_n N_A_3617_1198#_c_1505_n N_A_3617_1198#_c_1506_n
+ N_A_3617_1198#_c_1507_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_3617_1198#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_528_1171#
+ N_A_528_1171#_M1018_s N_A_528_1171#_M1027_s N_A_528_1171#_M1006_d
+ N_A_528_1171#_M1015_d N_A_528_1171#_M1004_g N_A_528_1171#_c_1613_n
+ N_A_528_1171#_c_1614_n N_A_528_1171#_M1010_g N_A_528_1171#_c_1616_n
+ N_A_528_1171#_M1023_g N_A_528_1171#_c_1618_n N_A_528_1171#_M1040_g
+ N_A_528_1171#_c_1620_n N_A_528_1171#_c_1646_n N_A_528_1171#_c_1647_n
+ N_A_528_1171#_c_1621_n N_A_528_1171#_c_1622_n N_A_528_1171#_c_1623_n
+ N_A_528_1171#_c_1624_n N_A_528_1171#_c_1625_n N_A_528_1171#_c_1626_n
+ N_A_528_1171#_M1007_g N_A_528_1171#_c_1655_n N_A_528_1171#_M1003_g
+ N_A_528_1171#_c_1659_n N_A_528_1171#_M1026_g N_A_528_1171#_M1009_g
+ N_A_528_1171#_c_1663_n N_A_528_1171#_M1035_g N_A_528_1171#_M1014_g
+ N_A_528_1171#_c_1667_n N_A_528_1171#_M1038_g N_A_528_1171#_M1016_g
+ N_A_528_1171#_c_1631_n N_A_528_1171#_c_1632_n N_A_528_1171#_c_1633_n
+ N_A_528_1171#_c_1634_n N_A_528_1171#_c_1635_n N_A_528_1171#_c_1636_n
+ N_A_528_1171#_c_1637_n N_A_528_1171#_c_1638_n N_A_528_1171#_c_1639_n
+ N_A_528_1171#_c_1682_n N_A_528_1171#_c_1640_n N_A_528_1171#_c_1641_n
+ N_A_528_1171#_c_1684_n N_A_528_1171#_c_1736_n N_A_528_1171#_c_1642_n
+ N_A_528_1171#_c_1688_n N_A_528_1171#_c_1690_n N_A_528_1171#_c_1691_n
+ N_A_528_1171#_c_1741_n N_A_528_1171#_c_1696_n N_A_528_1171#_c_1847_n
+ N_A_528_1171#_c_1643_n N_A_528_1171#_c_1644_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_528_1171#
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A N_A_c_1874_n N_A_c_1867_n
+ N_A_c_1876_n N_A_M1031_g N_A_M1024_g N_A_c_1869_n N_A_c_1870_n N_A_M1046_g
+ N_A_c_1883_n N_A_M1044_g N_A_c_1872_n A
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%X N_X_M1008_s N_X_M1030_s
+ N_X_M1005_s N_X_M1011_s N_X_c_1920_n N_X_c_1921_n N_X_c_1922_n N_X_c_1927_n
+ N_X_c_1958_n X PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%X
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%VPWR N_VPWR_M1005_d
+ N_VPWR_M1036_d N_VPWR_M39_noxref_d N_VPWR_M43_noxref_s N_VPWR_M44_noxref_d
+ N_VPWR_M46_noxref_d N_VPWR_M1020_d N_VPWR_c_1988_n N_VPWR_c_1990_n
+ N_VPWR_c_1992_n N_VPWR_c_1993_n N_VPWR_c_1994_n N_VPWR_c_1995_n
+ N_VPWR_c_1997_n N_VPWR_c_1998_n N_VPWR_c_1999_n N_VPWR_c_2000_n
+ N_VPWR_c_2001_n N_VPWR_c_2002_n N_VPWR_c_2003_n N_VPWR_c_2004_n
+ N_VPWR_c_2006_n N_VPWR_c_2007_n VPWR VPWR N_VPWR_c_2008_n N_VPWR_c_2009_n
+ N_VPWR_c_2117_n N_VPWR_c_2010_n N_VPWR_c_2118_n N_VPWR_c_2011_n
+ N_VPWR_c_2013_n N_VPWR_c_2015_n N_VPWR_c_2016_n N_VPWR_c_1981_n
+ N_VPWR_c_1982_n VPWR VPWR PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%VPWR
x_PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_1410_571#
+ N_A_1410_571#_M1022_d N_A_1410_571#_M43_noxref_d N_A_1410_571#_M45_noxref_d
+ N_A_1410_571#_c_2253_n N_A_1410_571#_c_2254_n N_A_1410_571#_c_2245_n
+ N_A_1410_571#_c_2246_n N_A_1410_571#_c_2247_n N_A_1410_571#_c_2257_n
+ N_A_1410_571#_c_2248_n N_A_1410_571#_c_2260_n N_A_1410_571#_c_2262_n
+ N_A_1410_571#_c_2263_n N_A_1410_571#_c_2249_n
+ PM_SKY130_FD_SC_HVL__LSBUFLV2HV_CLKISO_HLKG_3%A_1410_571#
cc_1 N_VNB_M1018_b VPB 0.114982f $X=-0.33 $Y=-0.265 $X2=0 $Y2=3.955
cc_2 N_VNB_M1018_b N_LVPWR_c_396_n 0.274064f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_3 N_VNB_M1018_b N_VGND_M1000_g 0.0542433f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_4 N_VNB_M1018_b N_VGND_c_590_n 0.0197738f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_5 N_VNB_M1018_b N_VGND_c_591_n 0.0431432f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_6 N_VNB_c_6_p N_VGND_c_591_n 6.57436e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_7 N_VNB_M1018_b N_VGND_c_593_n 0.00438934f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_8 N_VNB_M1018_b N_VGND_c_594_n 0.0697054f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_9 N_VNB_M1018_b N_VGND_c_595_n 0.0221881f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_10 N_VNB_c_10_p N_VGND_c_595_n 7.75064e-19 $X=24.72 $Y=0 $X2=0 $Y2=0
cc_11 N_VNB_M1018_b N_VGND_c_597_n 0.00578741f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_12 N_VNB_M1018_b N_VGND_c_598_n 0.0126108f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_13 N_VNB_M1018_b N_VGND_c_599_n 0.0216684f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_14 N_VNB_M1018_b N_VGND_c_600_n 0.0221881f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_15 N_VNB_c_10_p N_VGND_c_600_n 7.75064e-19 $X=24.72 $Y=0 $X2=0 $Y2=0
cc_16 N_VNB_M1018_b N_VGND_c_602_n 0.00590474f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_17 N_VNB_M1018_b N_VGND_c_603_n 0.00582151f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_18 N_VNB_M1018_b N_VGND_c_604_n 0.0195211f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_19 N_VNB_M1018_b N_VGND_c_605_n 0.0211102f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_20 N_VNB_M1018_b N_VGND_c_606_n 0.0195211f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_21 N_VNB_M1018_b N_VGND_c_607_n 0.0237351f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_22 N_VNB_M1018_b N_VGND_c_608_n 0.0597712f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_23 N_VNB_M1018_b N_VGND_c_609_n 0.0446987f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_24 N_VNB_M1018_b N_VGND_c_610_n 0.0204756f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_25 N_VNB_c_10_p N_VGND_c_610_n 8.95109e-19 $X=24.72 $Y=0 $X2=0 $Y2=0
cc_26 N_VNB_M1018_b N_VGND_c_612_n 0.0165579f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_27 N_VNB_M1018_b N_VGND_c_613_n 0.0191184f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_28 N_VNB_c_6_p N_VGND_c_613_n 8.95109e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_29 N_VNB_M1018_b N_VGND_c_615_n 0.0237061f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_30 N_VNB_M1018_b N_VGND_c_616_n 0.0353151f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_31 N_VNB_c_10_p N_VGND_c_616_n 0.00165372f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_32 N_VNB_M1018_b N_VGND_c_618_n 0.0348222f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_33 N_VNB_c_6_p N_VGND_c_618_n 0.00159855f $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_34 N_VNB_M1018_b N_VGND_c_620_n 0.0016092f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_35 N_VNB_M1018_b N_VGND_c_621_n 0.0016092f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_36 N_VNB_M1018_b N_VGND_c_622_n 0.0353151f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_37 N_VNB_c_6_p N_VGND_c_622_n 0.00165372f $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_38 N_VNB_M1018_b N_VGND_c_624_n 0.0348222f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_39 N_VNB_c_10_p N_VGND_c_624_n 0.00159855f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_40 N_VNB_M1018_b N_VGND_c_626_n 0.0191184f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_41 N_VNB_c_10_p N_VGND_c_626_n 8.95109e-19 $X=24.72 $Y=0 $X2=0 $Y2=0
cc_42 N_VNB_M1018_b N_VGND_c_628_n 0.0237061f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_43 N_VNB_M1018_b N_VGND_c_629_n 0.0123561f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_44 N_VNB_M1018_b N_VGND_c_630_n 0.0151705f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_45 N_VNB_c_6_p N_VGND_c_630_n 6.46887e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_46 N_VNB_M1018_b N_VGND_c_632_n 0.0113571f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_47 N_VNB_M1018_b N_VGND_c_633_n 0.0414003f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_48 N_VNB_c_6_p N_VGND_c_633_n 0.00190198f $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_49 N_VNB_M1018_b N_VGND_c_635_n 0.0162337f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_50 N_VNB_c_6_p N_VGND_c_635_n 6.78113e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_51 N_VNB_M1018_b N_VGND_c_637_n 0.0366696f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_52 N_VNB_M1018_b N_VGND_c_638_n 0.0134401f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_53 N_VNB_M1018_b N_VGND_c_639_n 0.00184939f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_54 N_VNB_M1018_b N_VGND_c_640_n 0.07514f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_55 N_VNB_c_6_p N_VGND_c_640_n 0.00323351f $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_56 N_VNB_M1018_b N_VGND_c_642_n 0.0134069f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_57 N_VNB_c_6_p N_VGND_c_642_n 6.57436e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_58 N_VNB_M1018_b N_VGND_c_644_n 0.1563f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_59 N_VNB_c_6_p N_VGND_c_644_n 0.00649835f $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_60 N_VNB_M1018_b N_VGND_c_646_n 0.0134069f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_61 N_VNB_c_6_p N_VGND_c_646_n 6.57436e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_62 N_VNB_M1018_b N_VGND_c_648_n 0.154118f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_63 N_VNB_c_6_p N_VGND_c_648_n 0.00640849f $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_64 N_VNB_M1018_b N_VGND_c_650_n 0.0134069f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_65 N_VNB_c_6_p N_VGND_c_650_n 6.57436e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_66 N_VNB_M1018_b N_VGND_c_652_n 0.154118f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_67 N_VNB_c_6_p N_VGND_c_652_n 0.00640849f $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_68 N_VNB_M1018_b N_VGND_c_654_n 0.0134069f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_69 N_VNB_c_6_p N_VGND_c_654_n 6.57436e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_70 N_VNB_M1018_b N_VGND_c_656_n 0.154118f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_71 N_VNB_c_6_p N_VGND_c_656_n 0.00640849f $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_72 N_VNB_M1018_b N_VGND_c_658_n 0.0134069f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_73 N_VNB_c_6_p N_VGND_c_658_n 6.57436e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_74 N_VNB_M1018_b N_VGND_c_660_n 0.0933458f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_75 N_VNB_c_6_p N_VGND_c_660_n 0.00384754f $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_76 N_VNB_M1018_b N_VGND_c_662_n 0.0134069f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_77 N_VNB_c_6_p N_VGND_c_662_n 6.57436e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_78 N_VNB_M1018_b N_VGND_c_664_n 0.0970044f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_79 N_VNB_c_6_p N_VGND_c_664_n 0.0039808f $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_80 N_VNB_M1018_b N_VGND_c_666_n 0.0161406f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_81 N_VNB_c_6_p N_VGND_c_666_n 8.95109e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_82 N_VNB_M1018_b N_VGND_c_668_n 0.0161406f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_83 N_VNB_c_10_p N_VGND_c_668_n 8.95109e-19 $X=24.72 $Y=0 $X2=0 $Y2=0
cc_84 N_VNB_M1018_b N_VGND_c_670_n 0.0174978f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_85 N_VNB_c_6_p N_VGND_c_670_n 8.95109e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_86 N_VNB_M1018_b N_VGND_c_672_n 0.0132559f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_87 N_VNB_c_6_p N_VGND_c_672_n 6.78113e-19 $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_88 N_VNB_M1018_b N_VGND_c_674_n 0.0360591f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_89 N_VNB_c_10_p N_VGND_c_674_n 0.00122924f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_90 N_VNB_M1018_b N_VGND_c_676_n 0.0360591f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_91 N_VNB_c_10_p N_VGND_c_676_n 0.00122924f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_92 N_VNB_M1018_b N_VGND_c_678_n 0.0588705f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_93 N_VNB_c_10_p N_VGND_c_678_n 0.00201575f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_94 N_VNB_M1018_b N_VGND_c_680_n 1.00005f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_95 N_VNB_c_10_p N_VGND_c_680_n 2.66844f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_96 N_VNB_M1018_b N_VGND_c_682_n 0.879115f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_97 N_VNB_c_6_p N_VGND_c_682_n 2.66841f $X=24.72 $Y=8.14 $X2=0 $Y2=0
cc_98 N_VNB_M1018_b N_A_262_107#_M1008_g 0.0644744f $X=-0.33 $Y=-0.265 $X2=0.36
+ $Y2=4.07
cc_99 N_VNB_c_10_p N_A_262_107#_M1008_g 0.00201121f $X=24.72 $Y=0 $X2=0.36
+ $Y2=4.07
cc_100 N_VNB_M1018_b N_A_262_107#_c_842_n 0.00773022f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_101 N_VNB_M1018_b N_A_262_107#_M1030_g 0.054067f $X=-0.33 $Y=-0.265 $X2=9.71
+ $Y2=4.07
cc_102 N_VNB_c_10_p N_A_262_107#_M1030_g 6.63698e-19 $X=24.72 $Y=0 $X2=9.71
+ $Y2=4.07
cc_103 N_VNB_M1018_b N_A_262_107#_c_845_n 0.00773022f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_104 N_VNB_M1018_b N_A_262_107#_M1047_g 0.053801f $X=-0.33 $Y=-0.265 $X2=9.71
+ $Y2=4.07
cc_105 N_VNB_c_10_p N_A_262_107#_M1047_g 6.63698e-19 $X=24.72 $Y=0 $X2=9.71
+ $Y2=4.07
cc_106 N_VNB_M1018_b N_A_262_107#_c_848_n 0.0134646f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_107 N_VNB_M1018_b N_A_262_107#_c_849_n 0.00875564f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_108 N_VNB_M1018_b N_A_262_107#_c_850_n 0.0107791f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_109 N_VNB_M1018_b N_A_262_107#_c_851_n 0.0354319f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_110 N_VNB_M1018_b N_A_262_107#_c_852_n 0.0119607f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_111 N_VNB_M1018_b N_A_262_107#_c_853_n 0.00102836f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_112 N_VNB_M1018_b N_A_262_107#_c_854_n 0.0183692f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_113 N_VNB_M1018_b N_A_262_107#_c_855_n 0.00118464f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_114 N_VNB_M1018_b N_A_840_107#_M1012_g 0.0596315f $X=-0.33 $Y=-0.265 $X2=0.36
+ $Y2=4.07
cc_115 N_VNB_c_10_p N_A_840_107#_M1012_g 0.00138773f $X=24.72 $Y=0 $X2=0.36
+ $Y2=4.07
cc_116 N_VNB_M1018_b N_A_840_107#_c_968_n 0.00788262f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_117 N_VNB_M1018_b N_A_840_107#_M1034_g 0.0598997f $X=-0.33 $Y=-0.265 $X2=9.71
+ $Y2=4.07
cc_118 N_VNB_c_10_p N_A_840_107#_M1034_g 0.00138773f $X=24.72 $Y=0 $X2=9.71
+ $Y2=4.07
cc_119 N_VNB_M1018_b N_A_840_107#_c_971_n 0.0511748f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_120 N_VNB_M1018_b N_A_840_107#_c_972_n 0.0136727f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_121 N_VNB_M1018_b N_A_840_107#_c_973_n 0.00981693f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_122 N_VNB_M1018_b N_A_840_107#_c_974_n 4.11818e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_123 N_VNB_M1018_b N_A_840_107#_c_975_n 0.00296628f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_124 N_VNB_M1018_b N_A_840_107#_c_976_n 0.0584349f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_125 N_VNB_M1018_b N_A_840_107#_c_977_n 0.00973381f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_126 N_VNB_M1018_b N_A_840_107#_c_978_n 0.00296628f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_127 N_VNB_M1018_b N_A_840_107#_c_979_n 0.0445768f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_128 N_VNB_M1018_b N_A_840_107#_c_980_n 0.0121968f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_129 N_VNB_M1018_b N_A_362_1243#_c_1123_n 0.0102797f $X=-0.33 $Y=-0.265
+ $X2=0.24 $Y2=4.07
cc_130 N_VNB_M1018_b N_A_362_1243#_c_1124_n 0.0388133f $X=-0.33 $Y=-0.265
+ $X2=9.71 $Y2=4.07
cc_131 N_VNB_M1018_b N_A_362_1243#_c_1125_n 0.0107502f $X=-0.33 $Y=-0.265
+ $X2=9.71 $Y2=4.07
cc_132 N_VNB_M1018_b N_A_362_1243#_c_1126_n 0.00296628f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_133 N_VNB_M1018_b N_A_362_1243#_c_1127_n 0.075507f $X=-0.33 $Y=-0.265 $X2=0.6
+ $Y2=4.07
cc_134 N_VNB_M1018_b N_A_362_1243#_c_1128_n 0.00296628f $X=-0.33 $Y=-0.265
+ $X2=0.6 $Y2=4.07
cc_135 N_VNB_M1018_b N_A_362_1243#_c_1129_n 4.11818e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_136 N_VNB_M1018_b N_A_362_1243#_c_1130_n 0.00682709f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_137 N_VNB_M1018_b N_A_2092_381#_M1002_g 0.0951986f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_138 N_VNB_M1018_b N_A_2092_381#_c_1216_n 0.0184295f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_139 N_VNB_M1018_b N_A_2092_381#_c_1217_n 0.0136621f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_140 N_VNB_M1018_b N_A_1472_1171#_M1001_g 0.0662291f $X=-0.33 $Y=-0.265
+ $X2=0.36 $Y2=4.07
cc_141 N_VNB_M1018_b N_A_1472_1171#_c_1312_n 0.0129209f $X=-0.33 $Y=-0.265
+ $X2=0.24 $Y2=4.07
cc_142 N_VNB_M1018_b N_A_1472_1171#_c_1313_n 0.035712f $X=-0.33 $Y=-0.265
+ $X2=0.24 $Y2=4.07
cc_143 N_VNB_M1018_b N_A_1472_1171#_M1029_g 0.0654137f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_144 N_VNB_M1018_b N_A_1472_1171#_c_1315_n 0.0462271f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_145 N_VNB_M1018_b N_A_1472_1171#_c_1316_n 0.32507f $X=-0.33 $Y=-0.265
+ $X2=9.71 $Y2=4.07
cc_146 N_VNB_M1018_b N_A_1472_1171#_c_1317_n 0.0118354f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_147 N_VNB_M1018_b N_A_1472_1171#_c_1318_n 0.0161013f $X=-0.33 $Y=-0.265
+ $X2=0.445 $Y2=4.07
cc_148 N_VNB_M1018_b N_A_1472_1171#_M1032_g 0.0654137f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_149 N_VNB_M1018_b N_A_1472_1171#_c_1320_n 0.0476809f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_150 N_VNB_M1018_b N_A_1472_1171#_M1041_g 0.0720582f $X=-0.33 $Y=-0.265
+ $X2=10.215 $Y2=4.07
cc_151 N_VNB_M1018_b N_A_1472_1171#_c_1322_n 0.0390805f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_152 N_VNB_M1018_b N_A_1472_1171#_c_1323_n 0.0418462f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_153 N_VNB_M1018_b N_A_1472_1171#_c_1324_n 0.0218673f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_154 N_VNB_M1018_b N_A_1472_1171#_c_1325_n 0.169779f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_155 N_VNB_M1018_b N_A_1472_1171#_c_1326_n 0.0011811f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_156 N_VNB_M1018_b N_A_1472_1171#_c_1327_n 0.0035469f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_157 N_VNB_M1018_b N_A_1472_1171#_c_1328_n 0.0108018f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_158 N_VNB_M1018_b N_A_1472_1171#_c_1329_n 0.0239872f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_159 N_VNB_M1018_b N_A_1472_1171#_c_1330_n 0.00189252f $X=-0.33 $Y=-0.265
+ $X2=0 $Y2=0
cc_160 N_VNB_M1018_b N_A_1472_1171#_c_1331_n 0.00127131f $X=-0.33 $Y=-0.265
+ $X2=0 $Y2=0
cc_161 N_VNB_M1018_b N_SLEEP_B_M1045_g 0.0742506f $X=-0.33 $Y=-0.265 $X2=-0.33
+ $Y2=1.885
cc_162 N_VNB_M1018_b N_SLEEP_B_c_1468_n 0.00935176f $X=-0.33 $Y=-0.265 $X2=0.445
+ $Y2=4.875
cc_163 N_VNB_M1018_b N_SLEEP_B_c_1469_n 0.0203608f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_164 N_VNB_M1018_b N_SLEEP_B_c_1470_n 0.00483784f $X=-0.33 $Y=-0.265 $X2=0.36
+ $Y2=4.07
cc_165 N_VNB_M1018_b N_A_3617_1198#_M1018_g 0.0261472f $X=-0.33 $Y=-0.265
+ $X2=0.445 $Y2=4.155
cc_166 N_VNB_M1018_b N_A_3617_1198#_M1019_g 0.0238903f $X=-0.33 $Y=-0.265
+ $X2=0.24 $Y2=4.07
cc_167 N_VNB_M1018_b N_A_3617_1198#_M1027_g 0.0238184f $X=-0.33 $Y=-0.265
+ $X2=9.71 $Y2=4.07
cc_168 N_VNB_M1018_b N_A_3617_1198#_M1033_g 0.031461f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_169 N_VNB_M1018_b N_A_3617_1198#_c_1500_n 0.00128362f $X=-0.33 $Y=-0.265
+ $X2=9.71 $Y2=4.07
cc_170 N_VNB_M1018_b N_A_3617_1198#_c_1501_n 0.022427f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_171 N_VNB_M1018_b N_A_3617_1198#_c_1502_n 5.85262e-19 $X=-0.33 $Y=-0.265
+ $X2=0 $Y2=0
cc_172 N_VNB_M1018_b N_A_3617_1198#_c_1503_n 8.20237e-19 $X=-0.33 $Y=-0.265
+ $X2=0 $Y2=0
cc_173 N_VNB_M1018_b N_A_3617_1198#_c_1504_n 0.00485792f $X=-0.33 $Y=-0.265
+ $X2=0 $Y2=0
cc_174 N_VNB_M1018_b N_A_3617_1198#_c_1505_n 7.07123e-19 $X=-0.33 $Y=-0.265
+ $X2=0 $Y2=0
cc_175 N_VNB_M1018_b N_A_3617_1198#_c_1506_n 0.00162535f $X=-0.33 $Y=-0.265
+ $X2=0 $Y2=0
cc_176 N_VNB_M1018_b N_A_3617_1198#_c_1507_n 0.0763371f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_177 N_VNB_M1018_b N_A_528_1171#_M1004_g 0.0692617f $X=-0.33 $Y=-0.265
+ $X2=0.36 $Y2=4.07
cc_178 N_VNB_M1018_b N_A_528_1171#_c_1613_n 0.0166478f $X=-0.33 $Y=-0.265
+ $X2=0.24 $Y2=4.07
cc_179 N_VNB_M1018_b N_A_528_1171#_c_1614_n 0.0437638f $X=-0.33 $Y=-0.265
+ $X2=0.24 $Y2=4.07
cc_180 N_VNB_M1018_b N_A_528_1171#_M1010_g 0.0654137f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_181 N_VNB_M1018_b N_A_528_1171#_c_1616_n 0.0161013f $X=-0.33 $Y=-0.265
+ $X2=9.71 $Y2=4.07
cc_182 N_VNB_M1018_b N_A_528_1171#_M1023_g 0.0654137f $X=-0.33 $Y=-0.265
+ $X2=0.445 $Y2=4.07
cc_183 N_VNB_M1018_b N_A_528_1171#_c_1618_n 0.0150914f $X=-0.33 $Y=-0.265
+ $X2=0.6 $Y2=4.07
cc_184 N_VNB_M1018_b N_A_528_1171#_M1040_g 0.0662291f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_185 N_VNB_M1018_b N_A_528_1171#_c_1620_n 0.00947027f $X=-0.33 $Y=-0.265
+ $X2=10.215 $Y2=4.07
cc_186 N_VNB_M1018_b N_A_528_1171#_c_1621_n 0.081416f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_187 N_VNB_M1018_b N_A_528_1171#_c_1622_n 0.698906f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_188 N_VNB_M1018_b N_A_528_1171#_c_1623_n 0.0236434f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_189 N_VNB_M1018_b N_A_528_1171#_c_1624_n 0.0513906f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_190 N_VNB_M1018_b N_A_528_1171#_c_1625_n 0.0212642f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_191 N_VNB_M1018_b N_A_528_1171#_c_1626_n 0.0153985f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_192 N_VNB_M1018_b N_A_528_1171#_M1007_g 0.0257667f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_193 N_VNB_M1018_b N_A_528_1171#_M1009_g 0.0238184f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_194 N_VNB_M1018_b N_A_528_1171#_M1014_g 0.0238903f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_195 N_VNB_M1018_b N_A_528_1171#_M1016_g 0.0261472f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_196 N_VNB_M1018_b N_A_528_1171#_c_1631_n 0.0447883f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_197 N_VNB_M1018_b N_A_528_1171#_c_1632_n 0.0447883f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_198 N_VNB_M1018_b N_A_528_1171#_c_1633_n 0.0419712f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_199 N_VNB_M1018_b N_A_528_1171#_c_1634_n 0.173529f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_200 N_VNB_M1018_b N_A_528_1171#_c_1635_n 0.0212025f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_201 N_VNB_M1018_b N_A_528_1171#_c_1636_n 0.00132306f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_202 N_VNB_M1018_b N_A_528_1171#_c_1637_n 0.00110578f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_203 N_VNB_M1018_b N_A_528_1171#_c_1638_n 0.0197102f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_204 N_VNB_M1018_b N_A_528_1171#_c_1639_n 0.0239872f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_205 N_VNB_M1018_b N_A_528_1171#_c_1640_n 0.00344971f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_206 N_VNB_M1018_b N_A_528_1171#_c_1641_n 0.00735212f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_207 N_VNB_M1018_b N_A_528_1171#_c_1642_n 0.00636659f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_208 N_VNB_M1018_b N_A_528_1171#_c_1643_n 0.00127131f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_209 N_VNB_M1018_b N_A_528_1171#_c_1644_n 0.0675185f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_210 N_VNB_M1018_b N_A_c_1867_n 0.0126875f $X=-0.33 $Y=-0.265 $X2=9.135
+ $Y2=3.985
cc_211 N_VNB_M1018_b N_A_M1024_g 0.0260771f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_212 N_VNB_M1018_b N_A_c_1869_n 0.00970685f $X=-0.33 $Y=-0.265 $X2=0.445
+ $Y2=4.875
cc_213 N_VNB_M1018_b N_A_c_1870_n 0.0575202f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_214 N_VNB_M1018_b N_A_M1046_g 0.0267421f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_215 N_VNB_M1018_b N_A_c_1872_n 0.00957891f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_216 N_VNB_M1018_b A 0.00655144f $X=-0.33 $Y=-0.265 $X2=0.24 $Y2=4.07
cc_217 N_VNB_M1018_b N_X_c_1920_n 0.0193153f $X=-0.33 $Y=-0.265 $X2=0.36
+ $Y2=4.07
cc_218 N_VNB_M1018_b N_X_c_1921_n 0.00637968f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_219 N_VNB_M1018_b N_X_c_1922_n 0.0114852f $X=-0.33 $Y=-0.265 $X2=9.71
+ $Y2=4.07
cc_220 N_VNB_M1018_b X 0.00758039f $X=-0.33 $Y=-0.265 $X2=0.6 $Y2=4.07
cc_221 N_VNB_M1018_b N_VPWR_c_1981_n 0.14065f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_222 N_VNB_M1018_b N_VPWR_c_1982_n 0.296931f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_223 N_VNB_M1018_b N_A_1410_571#_c_2245_n 0.0156926f $X=-0.33 $Y=-0.265
+ $X2=0.24 $Y2=4.07
cc_224 N_VNB_M1018_b N_A_1410_571#_c_2246_n 0.0950661f $X=-0.33 $Y=-0.265
+ $X2=0.24 $Y2=4.07
cc_225 N_VNB_M1018_b N_A_1410_571#_c_2247_n 0.0201989f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_226 N_VNB_M1018_b N_A_1410_571#_c_2248_n 0.0266458f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_227 N_VNB_M1018_b N_A_1410_571#_c_2249_n 0.00334172f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_228 VPB N_LVPWR_M1006_b 0.0298079f $X=0 $Y=3.955 $X2=0.24 $Y2=8.14
cc_229 VPB N_LVPWR_c_398_n 0.0731761f $X=0 $Y=3.955 $X2=24.72 $Y2=8.14
cc_230 VPB N_LVPWR_c_399_n 6.33813e-19 $X=0 $Y=3.955 $X2=24.72 $Y2=0
cc_231 VPB N_LVPWR_c_400_n 2.53444e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_232 VPB N_LVPWR_c_401_n 6.33813e-19 $X=0 $Y=3.955 $X2=0.24 $Y2=8.14
cc_233 VPB N_LVPWR_c_402_n 2.12267e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_234 VPB N_LVPWR_c_403_n 6.33457e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_235 VPB N_LVPWR_c_404_n 6.07368e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_236 VPB N_LVPWR_c_405_n 0.0476201f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_237 VPB N_LVPWR_c_406_n 0.00571296f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_238 N_VPB_M1005_b N_LVPWR_c_396_n 0.272057f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_239 N_VPB_M1005_b N_A_262_107#_M1005_g 0.0581844f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_240 VPB N_A_262_107#_M1005_g 0.0119381f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_241 N_VPB_M1005_b N_A_262_107#_c_842_n 0.00389472f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_242 N_VPB_M1005_b N_A_262_107#_M1011_g 0.0504539f $X=-0.33 $Y=1.885 $X2=0.24
+ $Y2=8.14
cc_243 VPB N_A_262_107#_M1011_g 0.0119381f $X=0 $Y=3.955 $X2=0.24 $Y2=8.14
cc_244 N_VPB_M1005_b N_A_262_107#_c_845_n 0.00389472f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_245 N_VPB_M1005_b N_A_262_107#_M1036_g 0.0499732f $X=-0.33 $Y=1.885 $X2=0.24
+ $Y2=0
cc_246 VPB N_A_262_107#_M1036_g 0.0119381f $X=0 $Y=3.955 $X2=0.24 $Y2=0
cc_247 N_VPB_M1005_b N_A_262_107#_c_848_n 0.00285612f $X=-0.33 $Y=1.885
+ $X2=10.215 $Y2=0
cc_248 N_VPB_M1005_b N_A_262_107#_c_849_n 0.00185726f $X=-0.33 $Y=1.885
+ $X2=10.215 $Y2=0
cc_249 N_VPB_M1005_b N_A_262_107#_c_850_n 0.0103511f $X=-0.33 $Y=1.885 $X2=12.48
+ $Y2=0
cc_250 N_VPB_M1005_b N_A_262_107#_c_851_n 0.0215782f $X=-0.33 $Y=1.885 $X2=0.24
+ $Y2=8.14
cc_251 N_VPB_M1005_b N_A_262_107#_c_868_n 0.00644265f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_252 VPB N_A_262_107#_c_868_n 0.00139266f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_253 N_VPB_M1005_b N_A_262_107#_c_853_n 0.00637968f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_254 N_VPB_M1005_b N_A_262_107#_c_871_n 0.00626133f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_255 VPB N_A_262_107#_c_871_n 0.00139266f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_256 N_VPB_M1005_b N_A_262_107#_c_855_n 8.48061e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_257 N_VPB_M1005_b N_A_262_107#_c_874_n 3.44689e-19 $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_258 VPB N_A_840_107#_M1043_d 7.10164e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_259 N_VPB_M1005_b N_A_840_107#_M39_noxref_g 0.0597635f $X=-0.33 $Y=1.885
+ $X2=0 $Y2=0
cc_260 VPB N_A_840_107#_M39_noxref_g 0.014036f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_261 N_VPB_M1005_b N_A_840_107#_c_968_n 0.00330464f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_262 N_VPB_M1005_b N_A_840_107#_M40_noxref_g 0.0573124f $X=-0.33 $Y=1.885
+ $X2=0.24 $Y2=8.14
cc_263 VPB N_A_840_107#_M40_noxref_g 0.0121759f $X=0 $Y=3.955 $X2=0.24 $Y2=8.14
cc_264 N_VPB_M1005_b N_A_840_107#_c_971_n 0.0110228f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_265 N_VPB_M1005_b N_A_840_107#_c_988_n 0.193027f $X=-0.33 $Y=1.885 $X2=24.72
+ $Y2=8.14
cc_266 VPB N_A_840_107#_c_988_n 0.0105961f $X=0 $Y=3.955 $X2=24.72 $Y2=8.14
cc_267 N_VPB_M1005_b N_A_840_107#_c_990_n 0.034671f $X=-0.33 $Y=1.885 $X2=24.72
+ $Y2=8.14
cc_268 N_VPB_M1005_b N_A_840_107#_c_991_n 0.0314051f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_269 N_VPB_M1005_b N_A_840_107#_M1022_g 0.0811596f $X=-0.33 $Y=1.885 $X2=0.24
+ $Y2=0
cc_270 VPB N_A_840_107#_M1022_g 0.0124384f $X=0 $Y=3.955 $X2=0.24 $Y2=0
cc_271 N_VPB_M1005_b N_A_840_107#_c_972_n 0.001105f $X=-0.33 $Y=1.885 $X2=10.215
+ $Y2=0
cc_272 N_VPB_M1005_b N_A_840_107#_c_973_n 7.95968e-19 $X=-0.33 $Y=1.885
+ $X2=10.215 $Y2=0
cc_273 N_VPB_M1005_b N_A_840_107#_c_996_n 0.0307062f $X=-0.33 $Y=1.885 $X2=24.72
+ $Y2=0
cc_274 N_VPB_M1005_b N_A_840_107#_c_997_n 0.0305807f $X=-0.33 $Y=1.885
+ $X2=10.215 $Y2=8.14
cc_275 VPB N_A_840_107#_c_997_n 0.023895f $X=0 $Y=3.955 $X2=10.215 $Y2=8.14
cc_276 N_VPB_M1005_b N_A_840_107#_c_974_n 0.0155181f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_277 N_VPB_M1005_b N_A_840_107#_c_979_n 0.00195276f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_278 N_VPB_M1005_b N_A_840_107#_c_1001_n 0.00379158f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_279 N_VPB_M1005_b N_A_840_107#_c_1002_n 0.0821097f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_280 N_VPB_M1005_b N_A_840_107#_c_1003_n 0.00195276f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_281 VPB N_A_362_1243#_M1022_s 7.10164e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_282 N_VPB_M1005_b N_A_362_1243#_M1043_g 0.0547578f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_283 VPB N_A_362_1243#_M1043_g 0.0124384f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_284 N_VPB_M1005_b N_A_362_1243#_c_1134_n 0.15526f $X=-0.33 $Y=1.885 $X2=0.24
+ $Y2=0
cc_285 N_VPB_M1005_b N_A_362_1243#_c_1125_n 0.00372344f $X=-0.33 $Y=1.885
+ $X2=24.72 $Y2=0
cc_286 N_VPB_M1005_b N_A_362_1243#_c_1129_n 0.0608486f $X=-0.33 $Y=1.885
+ $X2=10.215 $Y2=0
cc_287 VPB N_A_362_1243#_c_1129_n 0.023895f $X=0 $Y=3.955 $X2=10.215 $Y2=0
cc_288 N_VPB_M1005_b N_A_362_1243#_c_1138_n 0.0121311f $X=-0.33 $Y=1.885
+ $X2=24.72 $Y2=0
cc_289 N_VPB_M1005_b N_A_362_1243#_c_1139_n 0.0076747f $X=-0.33 $Y=1.885
+ $X2=10.215 $Y2=8.14
cc_290 N_VPB_M1005_b N_A_2092_381#_M43_noxref_g 0.0686961f $X=-0.33 $Y=1.885
+ $X2=-0.33 $Y2=-0.265
cc_291 VPB N_A_2092_381#_M43_noxref_g 0.0119896f $X=0 $Y=3.955 $X2=-0.33
+ $Y2=-0.265
cc_292 N_VPB_M1005_b N_A_2092_381#_c_1220_n 0.0134555f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_293 N_VPB_M1005_b N_A_2092_381#_c_1221_n 0.0322899f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=8.025
cc_294 N_VPB_M1005_b N_A_2092_381#_M44_noxref_g 0.0552111f $X=-0.33 $Y=1.885
+ $X2=0 $Y2=0
cc_295 VPB N_A_2092_381#_M44_noxref_g 0.0119896f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_296 N_VPB_M1005_b N_A_2092_381#_c_1224_n 0.0150582f $X=-0.33 $Y=1.885
+ $X2=0.24 $Y2=0
cc_297 N_VPB_M1005_b N_A_2092_381#_M45_noxref_g 0.0552111f $X=-0.33 $Y=1.885
+ $X2=0 $Y2=0
cc_298 VPB N_A_2092_381#_M45_noxref_g 0.0119896f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_299 N_VPB_M1005_b N_A_2092_381#_c_1227_n 0.0162979f $X=-0.33 $Y=1.885
+ $X2=24.72 $Y2=0
cc_300 N_VPB_M1005_b N_A_2092_381#_M46_noxref_g 0.0634363f $X=-0.33 $Y=1.885
+ $X2=0 $Y2=0
cc_301 VPB N_A_2092_381#_M46_noxref_g 0.0119896f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_302 N_VPB_M1005_b N_A_2092_381#_c_1230_n 0.0201302f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_303 N_VPB_M1005_b N_A_2092_381#_c_1231_n 0.0243788f $X=-0.33 $Y=1.885
+ $X2=24.72 $Y2=8.14
cc_304 N_VPB_M1005_b N_A_2092_381#_c_1232_n 0.0241151f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_305 N_VPB_M1005_b N_A_2092_381#_c_1233_n 0.00924261f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_306 N_VPB_M1005_b N_A_2092_381#_c_1216_n 0.0564348f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_307 N_VPB_M1005_b N_A_2092_381#_c_1235_n 0.0140467f $X=-0.33 $Y=1.885
+ $X2=24.72 $Y2=0
cc_308 VPB N_A_2092_381#_c_1235_n 0.0079246f $X=0 $Y=3.955 $X2=24.72 $Y2=0
cc_309 N_VPB_M1005_b N_A_2092_381#_c_1237_n 0.00462492f $X=-0.33 $Y=1.885
+ $X2=12.48 $Y2=8.14
cc_310 N_VPB_M1005_b N_A_1472_1171#_c_1315_n 0.304781f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_311 VPB N_A_1472_1171#_c_1315_n 0.0108513f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_312 N_VPB_c_313_p N_A_1472_1171#_c_1315_n 0.00509221f $X=9.71 $Y=4.07 $X2=0
+ $Y2=0
cc_313 N_VPB_M1005_b N_A_1472_1171#_c_1335_n 0.0133586f $X=-0.33 $Y=1.885
+ $X2=24.72 $Y2=0
cc_314 N_VPB_M1005_b N_A_1472_1171#_c_1324_n 0.0812691f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_315 N_VPB_M1005_b N_SLEEP_B_M1020_g 0.0994468f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_316 VPB N_SLEEP_B_M1020_g 0.0106055f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_317 N_VPB_M1005_b N_SLEEP_B_c_1468_n 0.0159727f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_318 N_VPB_M1005_b N_SLEEP_B_c_1469_n 0.026842f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_319 N_VPB_M1005_b N_SLEEP_B_c_1470_n 0.0084967f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_320 N_VPB_M1005_b N_A_528_1171#_c_1620_n 0.0104579f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_321 N_VPB_M1005_b N_A_528_1171#_c_1646_n 0.0843457f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_322 N_VPB_M1005_b N_A_528_1171#_c_1647_n 0.0136449f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_323 N_VPB_M1005_b N_A_528_1171#_c_1621_n 0.206826f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_324 VPB N_A_528_1171#_c_1621_n 0.00916008f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_325 VPB N_A_528_1171#_c_1634_n 0.0237634f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_326 VPB N_X_M1005_s 7.10164e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_327 VPB N_X_M1011_s 9.03845e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_328 N_VPB_M1005_b N_X_c_1921_n 0.00637968f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_329 N_VPB_M1005_b N_X_c_1927_n 0.00592869f $X=-0.33 $Y=1.885 $X2=0.24
+ $Y2=8.14
cc_330 VPB N_X_c_1927_n 0.0221482f $X=0 $Y=3.955 $X2=0.24 $Y2=8.14
cc_331 N_VPB_M1005_b X 0.0159591f $X=-0.33 $Y=1.885 $X2=24.72 $Y2=8.14
cc_332 N_VPB_c_333_p X 0.025006f $X=0.445 $Y=4.875 $X2=24.72 $Y2=8.14
cc_333 VPB X 0.0213977f $X=0 $Y=3.955 $X2=24.72 $Y2=8.14
cc_334 N_VPB_c_335_p X 0.00500364f $X=0.6 $Y=4.07 $X2=24.72 $Y2=8.14
cc_335 VPB N_VPWR_M1005_d 5.79313e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_336 VPB N_VPWR_M1036_d 4.28188e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_337 VPB N_VPWR_M43_noxref_s 5.54125e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_338 VPB N_VPWR_M44_noxref_d 7.05251e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_339 VPB N_VPWR_M46_noxref_d 5.54125e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_340 N_VPB_M1005_b N_VPWR_c_1988_n 0.00267608f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_341 VPB N_VPWR_c_1988_n 0.0223893f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_342 N_VPB_M1005_b N_VPWR_c_1990_n 0.00204917f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_343 VPB N_VPWR_c_1990_n 0.0241379f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_344 VPB N_VPWR_c_1992_n 0.00146138f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_345 N_VPB_M1005_b N_VPWR_c_1993_n 0.00268475f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_346 N_VPB_M1005_b N_VPWR_c_1994_n 0.00273109f $X=-0.33 $Y=1.885 $X2=24.72
+ $Y2=0
cc_347 VPB N_VPWR_c_1995_n 0.0209049f $X=0 $Y=3.955 $X2=10.215 $Y2=8.14
cc_348 N_VPB_c_313_p N_VPWR_c_1995_n 0.00688562f $X=9.71 $Y=4.07 $X2=10.215
+ $Y2=8.14
cc_349 N_VPB_M1005_b N_VPWR_c_1997_n 0.00740878f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_350 N_VPB_M1005_b N_VPWR_c_1998_n 0.0120819f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_351 N_VPB_M1005_b N_VPWR_c_1999_n 0.00218996f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_352 VPB N_VPWR_c_2000_n 0.0219246f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_353 N_VPB_M1005_b N_VPWR_c_2001_n 0.0124759f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_354 N_VPB_M1005_b N_VPWR_c_2002_n 0.00377265f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_355 VPB N_VPWR_c_2003_n 0.023645f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_356 N_VPB_M1005_b N_VPWR_c_2004_n 0.00373058f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_357 VPB N_VPWR_c_2004_n 0.00836082f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_358 N_VPB_M1005_b N_VPWR_c_2006_n 0.00352682f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_359 N_VPB_M1005_b N_VPWR_c_2007_n 0.00260086f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_360 VPB N_VPWR_c_2008_n 0.00485676f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_361 VPB N_VPWR_c_2009_n 0.00485652f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_362 VPB N_VPWR_c_2010_n 0.00472006f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_363 N_VPB_M1005_b N_VPWR_c_2011_n 0.00874617f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_364 VPB N_VPWR_c_2011_n 0.00358511f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_365 N_VPB_M1005_b N_VPWR_c_2013_n 0.00874617f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_366 VPB N_VPWR_c_2013_n 0.00364598f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_367 VPB N_VPWR_c_2015_n 0.00478093f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_368 N_VPB_M1005_b N_VPWR_c_2016_n 0.00874617f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_369 VPB N_VPWR_c_2016_n 0.00364598f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_370 N_VPB_M1005_b N_VPWR_c_1981_n 0.119804f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_371 VPB N_VPWR_c_1981_n 2.5949f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_372 N_VPB_c_373_p N_VPWR_c_1981_n 0.00524668f $X=0.36 $Y=4.07 $X2=0 $Y2=0
cc_373 N_VPB_c_313_p N_VPWR_c_1981_n 0.00605652f $X=9.71 $Y=4.07 $X2=0 $Y2=0
cc_374 N_VPB_M1005_b N_VPWR_c_1982_n 0.322817f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_375 N_VPB_c_333_p N_VPWR_c_1982_n 0.036829f $X=0.445 $Y=4.875 $X2=0 $Y2=0
cc_376 VPB N_VPWR_c_1982_n 2.59205f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_377 N_VPB_c_373_p N_VPWR_c_1982_n 0.00275993f $X=0.36 $Y=4.07 $X2=0 $Y2=0
cc_378 N_VPB_c_313_p N_VPWR_c_1982_n 0.00605652f $X=9.71 $Y=4.07 $X2=0 $Y2=0
cc_379 N_VPB_c_335_p N_VPWR_c_1982_n 0.00127427f $X=0.6 $Y=4.07 $X2=0 $Y2=0
cc_380 VPB N_A_1410_571#_M1022_d 7.42444e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_381 VPB N_A_1410_571#_M43_noxref_d 9.03845e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_382 VPB N_A_1410_571#_M45_noxref_d 9.03845e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_383 VPB N_A_1410_571#_c_2253_n 0.0226784f $X=0 $Y=3.955 $X2=0 $Y2=8.025
cc_384 N_VPB_M1005_b N_A_1410_571#_c_2254_n 0.0041183f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_385 N_VPB_M1005_b N_A_1410_571#_c_2245_n 0.00436436f $X=-0.33 $Y=1.885
+ $X2=0.24 $Y2=0
cc_386 N_VPB_M1005_b N_A_1410_571#_c_2246_n 0.0430425f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_387 N_VPB_M1005_b N_A_1410_571#_c_2257_n 0.011256f $X=-0.33 $Y=1.885
+ $X2=24.72 $Y2=0
cc_388 VPB N_A_1410_571#_c_2257_n 0.022201f $X=0 $Y=3.955 $X2=24.72 $Y2=0
cc_389 N_VPB_M1005_b N_A_1410_571#_c_2248_n 0.0257274f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_390 N_VPB_M1005_b N_A_1410_571#_c_2260_n 0.011256f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_391 VPB N_A_1410_571#_c_2260_n 0.022201f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_392 N_VPB_M1005_b N_A_1410_571#_c_2262_n 0.00193709f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_393 N_VPB_M1005_b N_A_1410_571#_c_2263_n 0.0058983f $X=-0.33 $Y=1.885
+ $X2=10.215 $Y2=0
cc_394 N_VPB_M1005_b N_A_1410_571#_c_2249_n 8.13705e-19 $X=-0.33 $Y=1.885
+ $X2=12.48 $Y2=0
cc_395 N_LVPWR_c_396_n N_A_262_107#_M39_noxref_s 0.00214577f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_396 N_LVPWR_c_396_n N_A_262_107#_M40_noxref_d 0.00214577f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_397 N_LVPWR_c_396_n N_A_262_107#_M1005_g 0.0308092f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_398 N_LVPWR_c_396_n N_A_262_107#_M1011_g 0.0308092f $X=20.245 $Y=3.155
+ $X2=0.24 $Y2=8.14
cc_399 N_LVPWR_c_396_n N_A_262_107#_M1036_g 0.0308092f $X=20.245 $Y=3.155
+ $X2=0.24 $Y2=0
cc_400 N_LVPWR_c_396_n N_A_262_107#_c_868_n 0.0335159f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_401 N_LVPWR_c_396_n N_A_262_107#_c_871_n 0.0354358f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_402 N_LVPWR_c_396_n N_A_840_107#_M1043_d 0.00214577f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_403 N_LVPWR_c_396_n N_A_840_107#_M39_noxref_g 0.0308092f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_404 N_LVPWR_c_396_n N_A_840_107#_M40_noxref_g 0.0297368f $X=20.245 $Y=3.155
+ $X2=0.24 $Y2=8.14
cc_405 N_LVPWR_c_396_n N_A_840_107#_c_988_n 0.0181201f $X=20.245 $Y=3.155
+ $X2=24.72 $Y2=8.14
cc_406 N_LVPWR_c_396_n N_A_840_107#_M1022_g 0.0155174f $X=20.245 $Y=3.155
+ $X2=0.24 $Y2=0
cc_407 N_LVPWR_c_396_n N_A_840_107#_c_997_n 0.0356305f $X=20.245 $Y=3.155
+ $X2=10.215 $Y2=8.14
cc_408 N_LVPWR_c_396_n N_A_362_1243#_M1022_s 0.00136103f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_409 N_LVPWR_c_396_n N_A_362_1243#_M1043_g 0.0136213f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_410 N_LVPWR_c_396_n N_A_362_1243#_c_1134_n 0.00317928f $X=20.245 $Y=3.155
+ $X2=0.24 $Y2=0
cc_411 N_LVPWR_c_396_n N_A_362_1243#_c_1129_n 0.0302944f $X=20.245 $Y=3.155
+ $X2=10.215 $Y2=0
cc_412 N_LVPWR_c_396_n N_A_362_1243#_c_1144_n 0.0144491f $X=20.245 $Y=3.155
+ $X2=0.24 $Y2=8.14
cc_413 N_LVPWR_c_396_n N_A_2092_381#_M43_noxref_g 0.0303711f $X=20.245 $Y=3.155
+ $X2=-0.33 $Y2=-0.265
cc_414 N_LVPWR_c_396_n N_A_2092_381#_M44_noxref_g 0.0303711f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_415 N_LVPWR_c_396_n N_A_2092_381#_M45_noxref_g 0.0303711f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_416 N_LVPWR_c_396_n N_A_2092_381#_M46_noxref_g 0.0303711f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_417 N_LVPWR_c_396_n N_A_1472_1171#_c_1315_n 0.0196295f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_418 N_LVPWR_c_431_p N_A_1472_1171#_c_1338_n 0.0121024f $X=17.98 $Y=2.5
+ $X2=10.215 $Y2=8.14
cc_419 N_LVPWR_M1006_b N_A_1472_1171#_c_1339_n 0.00220879f $X=17.395 $Y=2.045
+ $X2=24.72 $Y2=8.14
cc_420 N_LVPWR_c_431_p N_A_1472_1171#_c_1339_n 0.05467f $X=17.98 $Y=2.5
+ $X2=24.72 $Y2=8.14
cc_421 N_LVPWR_c_401_n N_A_1472_1171#_c_1339_n 0.0235488f $X=18.795 $Y=3.62
+ $X2=24.72 $Y2=8.14
cc_422 N_LVPWR_c_435_p N_A_1472_1171#_c_1339_n 0.0424688f $X=18.88 $Y=2.84
+ $X2=24.72 $Y2=8.14
cc_423 N_LVPWR_c_396_n N_A_1472_1171#_c_1339_n 0.0370826f $X=20.245 $Y=3.155
+ $X2=24.72 $Y2=8.14
cc_424 N_LVPWR_M1026_s N_A_1472_1171#_c_1344_n 0.00370197f $X=18.73 $Y=2.225
+ $X2=0 $Y2=0
cc_425 N_LVPWR_c_435_p N_A_1472_1171#_c_1344_n 0.013264f $X=18.88 $Y=2.84 $X2=0
+ $Y2=0
cc_426 N_LVPWR_c_396_n N_A_1472_1171#_c_1344_n 0.0127011f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_427 N_LVPWR_M1006_b N_A_1472_1171#_c_1347_n 0.00220879f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_428 N_LVPWR_c_435_p N_A_1472_1171#_c_1347_n 0.0424688f $X=18.88 $Y=2.84 $X2=0
+ $Y2=0
cc_429 N_LVPWR_c_404_n N_A_1472_1171#_c_1347_n 0.0235488f $X=19.665 $Y=3.62
+ $X2=0 $Y2=0
cc_430 N_LVPWR_c_405_n N_A_1472_1171#_c_1347_n 0.0207642f $X=20.042 $Y=4.605
+ $X2=0 $Y2=0
cc_431 N_LVPWR_c_444_p N_A_1472_1171#_c_1347_n 0.0230985f $X=19.78 $Y=2.84 $X2=0
+ $Y2=0
cc_432 N_LVPWR_c_396_n N_A_1472_1171#_c_1347_n 0.0370688f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_433 N_LVPWR_M1038_s N_A_1472_1171#_c_1353_n 0.00452537f $X=19.63 $Y=2.225
+ $X2=0 $Y2=0
cc_434 N_LVPWR_M1006_b N_A_1472_1171#_c_1353_n 0.00714046f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_435 N_LVPWR_c_444_p N_A_1472_1171#_c_1353_n 0.0210982f $X=19.78 $Y=2.84 $X2=0
+ $Y2=0
cc_436 N_LVPWR_c_396_n N_A_1472_1171#_c_1353_n 0.0070151f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_437 N_LVPWR_M1038_s N_A_1472_1171#_c_1329_n 0.00194528f $X=19.63 $Y=2.225
+ $X2=0 $Y2=0
cc_438 N_LVPWR_M1006_b N_A_1472_1171#_c_1329_n 0.0129845f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_439 N_LVPWR_M1006_b N_A_3617_1198#_c_1508_n 0.0165822f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_440 N_LVPWR_c_453_p N_A_3617_1198#_c_1508_n 0.00697554f $X=17.95 $Y=4.94
+ $X2=0 $Y2=0
cc_441 N_LVPWR_c_399_n N_A_3617_1198#_c_1508_n 0.00525604f $X=18.765 $Y=4.52
+ $X2=0 $Y2=0
cc_442 N_LVPWR_M1006_b N_A_3617_1198#_c_1511_n 0.0153181f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_443 N_LVPWR_c_399_n N_A_3617_1198#_c_1511_n 0.00525604f $X=18.765 $Y=4.52
+ $X2=0 $Y2=0
cc_444 N_LVPWR_c_457_p N_A_3617_1198#_c_1511_n 0.00477471f $X=18.85 $Y=4.94
+ $X2=0 $Y2=0
cc_445 N_LVPWR_M1006_b N_A_3617_1198#_c_1514_n 0.0153204f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_446 N_LVPWR_c_457_p N_A_3617_1198#_c_1514_n 0.00477471f $X=18.85 $Y=4.94
+ $X2=0 $Y2=0
cc_447 N_LVPWR_c_403_n N_A_3617_1198#_c_1514_n 0.00525604f $X=19.665 $Y=4.52
+ $X2=0 $Y2=0
cc_448 N_LVPWR_M1006_b N_A_3617_1198#_c_1517_n 0.0178427f $X=17.395 $Y=2.045
+ $X2=0.24 $Y2=8.14
cc_449 N_LVPWR_c_403_n N_A_3617_1198#_c_1517_n 0.00525604f $X=19.665 $Y=4.52
+ $X2=0.24 $Y2=8.14
cc_450 N_LVPWR_c_463_p N_A_3617_1198#_c_1517_n 0.0080034f $X=19.75 $Y=4.94
+ $X2=0.24 $Y2=8.14
cc_451 N_LVPWR_c_464_p N_A_3617_1198#_c_1517_n 0.00274422f $X=19.75 $Y=5.64
+ $X2=0.24 $Y2=8.14
cc_452 N_LVPWR_M1006_b N_A_3617_1198#_c_1500_n 0.0113953f $X=17.395 $Y=2.045
+ $X2=24.72 $Y2=8.14
cc_453 N_LVPWR_c_464_p N_A_3617_1198#_c_1500_n 0.0242571f $X=19.75 $Y=5.64
+ $X2=24.72 $Y2=8.14
cc_454 N_LVPWR_c_464_p N_A_3617_1198#_c_1501_n 0.0276992f $X=19.75 $Y=5.64
+ $X2=12.48 $Y2=0
cc_455 N_LVPWR_M1006_b N_A_3617_1198#_c_1502_n 0.00378227f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_456 N_LVPWR_c_463_p N_A_3617_1198#_c_1502_n 0.0478139f $X=19.75 $Y=4.94 $X2=0
+ $Y2=0
cc_457 N_LVPWR_c_406_n N_A_3617_1198#_c_1502_n 0.0203363f $X=21.07 $Y=4.52 $X2=0
+ $Y2=0
cc_458 N_LVPWR_c_471_p N_A_3617_1198#_c_1502_n 0.0394212f $X=21.235 $Y=4.94
+ $X2=0 $Y2=0
cc_459 N_LVPWR_c_464_p N_A_3617_1198#_c_1502_n 0.0365766f $X=19.75 $Y=5.64 $X2=0
+ $Y2=0
cc_460 N_LVPWR_M1006_b N_A_3617_1198#_c_1504_n 0.00396f $X=17.395 $Y=2.045 $X2=0
+ $Y2=0
cc_461 N_LVPWR_M1006_b N_A_3617_1198#_c_1507_n 0.0481502f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_462 N_LVPWR_c_396_n N_A_528_1171#_c_1621_n 0.0175339f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_463 N_LVPWR_M1006_b N_A_528_1171#_c_1625_n 0.0137498f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_464 N_LVPWR_c_431_p N_A_528_1171#_c_1625_n 0.00152596f $X=17.98 $Y=2.5 $X2=0
+ $Y2=0
cc_465 N_LVPWR_M1006_b N_A_528_1171#_c_1626_n 0.00670308f $X=17.395 $Y=2.045
+ $X2=0.24 $Y2=8.14
cc_466 N_LVPWR_M1006_b N_A_528_1171#_c_1655_n 0.0181926f $X=17.395 $Y=2.045
+ $X2=24.72 $Y2=8.14
cc_467 N_LVPWR_c_431_p N_A_528_1171#_c_1655_n 0.00795889f $X=17.98 $Y=2.5
+ $X2=24.72 $Y2=8.14
cc_468 N_LVPWR_c_401_n N_A_528_1171#_c_1655_n 0.00525604f $X=18.795 $Y=3.62
+ $X2=24.72 $Y2=8.14
cc_469 N_LVPWR_c_396_n N_A_528_1171#_c_1655_n 0.00671336f $X=20.245 $Y=3.155
+ $X2=24.72 $Y2=8.14
cc_470 N_LVPWR_M1006_b N_A_528_1171#_c_1659_n 0.0153204f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_471 N_LVPWR_c_401_n N_A_528_1171#_c_1659_n 0.00525604f $X=18.795 $Y=3.62
+ $X2=0 $Y2=0
cc_472 N_LVPWR_c_435_p N_A_528_1171#_c_1659_n 0.00463487f $X=18.88 $Y=2.84 $X2=0
+ $Y2=0
cc_473 N_LVPWR_c_396_n N_A_528_1171#_c_1659_n 0.00272136f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_474 N_LVPWR_M1006_b N_A_528_1171#_c_1663_n 0.0153181f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_475 N_LVPWR_c_435_p N_A_528_1171#_c_1663_n 0.00463487f $X=18.88 $Y=2.84 $X2=0
+ $Y2=0
cc_476 N_LVPWR_c_404_n N_A_528_1171#_c_1663_n 0.00525604f $X=19.665 $Y=3.62
+ $X2=0 $Y2=0
cc_477 N_LVPWR_c_396_n N_A_528_1171#_c_1663_n 0.00272136f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_478 N_LVPWR_M1006_b N_A_528_1171#_c_1667_n 0.0165817f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_479 N_LVPWR_c_404_n N_A_528_1171#_c_1667_n 0.00525604f $X=19.665 $Y=3.62
+ $X2=0 $Y2=0
cc_480 N_LVPWR_c_405_n N_A_528_1171#_c_1667_n 0.00631272f $X=20.042 $Y=4.605
+ $X2=0 $Y2=0
cc_481 N_LVPWR_c_396_n N_A_528_1171#_c_1667_n 0.00269582f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_482 N_LVPWR_c_453_p N_A_528_1171#_c_1634_n 0.03606f $X=17.95 $Y=4.94 $X2=0
+ $Y2=0
cc_483 N_LVPWR_c_398_n N_A_528_1171#_c_1634_n 0.0109568f $X=19.665 $Y=4.07 $X2=0
+ $Y2=0
cc_484 N_LVPWR_c_431_p N_A_528_1171#_c_1634_n 0.0441987f $X=17.98 $Y=2.5 $X2=0
+ $Y2=0
cc_485 N_LVPWR_c_400_n N_A_528_1171#_c_1634_n 0.00509394f $X=18.035 $Y=4.52
+ $X2=0 $Y2=0
cc_486 N_LVPWR_c_402_n N_A_528_1171#_c_1634_n 0.00467594f $X=18.065 $Y=3.62
+ $X2=0 $Y2=0
cc_487 N_LVPWR_c_396_n N_A_528_1171#_c_1634_n 0.037739f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_488 N_LVPWR_M1006_b N_A_528_1171#_c_1636_n 0.0294012f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_489 N_LVPWR_c_431_p N_A_528_1171#_c_1636_n 0.0219559f $X=17.98 $Y=2.5 $X2=0
+ $Y2=0
cc_490 N_LVPWR_M1006_b N_A_528_1171#_c_1637_n 0.0311198f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_491 N_LVPWR_M1006_s N_A_528_1171#_c_1639_n 0.00105295f $X=17.805 $Y=4.795
+ $X2=0 $Y2=0
cc_492 N_LVPWR_M1006_b N_A_528_1171#_c_1639_n 0.0111759f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_493 N_LVPWR_M1006_s N_A_528_1171#_c_1682_n 0.00132101f $X=17.805 $Y=4.795
+ $X2=0 $Y2=0
cc_494 N_LVPWR_c_453_p N_A_528_1171#_c_1682_n 0.00110254f $X=17.95 $Y=4.94 $X2=0
+ $Y2=0
cc_495 N_LVPWR_M1006_b N_A_528_1171#_c_1684_n 0.00220879f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_496 N_LVPWR_c_453_p N_A_528_1171#_c_1684_n 0.0462948f $X=17.95 $Y=4.94 $X2=0
+ $Y2=0
cc_497 N_LVPWR_c_399_n N_A_528_1171#_c_1684_n 0.0235488f $X=18.765 $Y=4.52 $X2=0
+ $Y2=0
cc_498 N_LVPWR_c_457_p N_A_528_1171#_c_1684_n 0.0449718f $X=18.85 $Y=4.94 $X2=0
+ $Y2=0
cc_499 N_LVPWR_M1013_s N_A_528_1171#_c_1688_n 0.00408911f $X=18.7 $Y=4.795 $X2=0
+ $Y2=0
cc_500 N_LVPWR_c_457_p N_A_528_1171#_c_1688_n 0.0136682f $X=18.85 $Y=4.94 $X2=0
+ $Y2=0
cc_501 N_LVPWR_c_464_p N_A_528_1171#_c_1690_n 0.013092f $X=19.75 $Y=5.64 $X2=0
+ $Y2=0
cc_502 N_LVPWR_M1006_b N_A_528_1171#_c_1691_n 0.00220879f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_503 N_LVPWR_c_457_p N_A_528_1171#_c_1691_n 0.0449718f $X=18.85 $Y=4.94 $X2=0
+ $Y2=0
cc_504 N_LVPWR_c_403_n N_A_528_1171#_c_1691_n 0.0235488f $X=19.665 $Y=4.52 $X2=0
+ $Y2=0
cc_505 N_LVPWR_c_463_p N_A_528_1171#_c_1691_n 0.0473746f $X=19.75 $Y=4.94 $X2=0
+ $Y2=0
cc_506 N_LVPWR_c_464_p N_A_528_1171#_c_1691_n 0.0150435f $X=19.75 $Y=5.64 $X2=0
+ $Y2=0
cc_507 N_LVPWR_M1006_s N_A_528_1171#_c_1696_n 0.00443371f $X=17.805 $Y=4.795
+ $X2=0 $Y2=0
cc_508 N_LVPWR_M1006_b N_A_528_1171#_c_1696_n 2.62635e-19 $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_509 N_LVPWR_c_453_p N_A_528_1171#_c_1696_n 0.0207902f $X=17.95 $Y=4.94 $X2=0
+ $Y2=0
cc_510 N_LVPWR_M1006_b N_A_528_1171#_c_1644_n 0.0475794f $X=17.395 $Y=2.045
+ $X2=0 $Y2=0
cc_511 N_LVPWR_M1006_b N_A_c_1874_n 0.00673933f $X=17.395 $Y=2.045 $X2=0 $Y2=0
cc_512 N_LVPWR_M1006_b N_A_c_1867_n 8.58417e-19 $X=17.395 $Y=2.045 $X2=0 $Y2=0
cc_513 N_LVPWR_M1006_b N_A_c_1876_n 0.017409f $X=17.395 $Y=2.045 $X2=0 $Y2=0
cc_514 N_LVPWR_c_463_p N_A_c_1876_n 0.00685525f $X=19.75 $Y=4.94 $X2=0 $Y2=0
cc_515 N_LVPWR_c_406_n N_A_c_1876_n 0.0051848f $X=21.07 $Y=4.52 $X2=0 $Y2=0
cc_516 N_LVPWR_c_471_p N_A_c_1876_n 6.46346e-19 $X=21.235 $Y=4.94 $X2=0 $Y2=0
cc_517 N_LVPWR_c_464_p N_A_c_1876_n 0.00290686f $X=19.75 $Y=5.64 $X2=0 $Y2=0
cc_518 N_LVPWR_M1006_b N_A_c_1870_n 0.00802803f $X=17.395 $Y=2.045 $X2=0
+ $Y2=8.025
cc_519 N_LVPWR_c_471_p N_A_c_1870_n 0.00155503f $X=21.235 $Y=4.94 $X2=0
+ $Y2=8.025
cc_520 N_LVPWR_M1006_b N_A_c_1883_n 0.018729f $X=17.395 $Y=2.045 $X2=0.24 $Y2=0
cc_521 N_LVPWR_c_406_n N_A_c_1883_n 0.00489337f $X=21.07 $Y=4.52 $X2=0.24 $Y2=0
cc_522 N_LVPWR_c_471_p N_A_c_1883_n 0.0147417f $X=21.235 $Y=4.94 $X2=0.24 $Y2=0
cc_523 N_LVPWR_M1006_b A 0.00739755f $X=17.395 $Y=2.045 $X2=0 $Y2=0
cc_524 N_LVPWR_c_471_p A 0.026709f $X=21.235 $Y=4.94 $X2=0 $Y2=0
cc_525 N_LVPWR_c_396_n N_X_M1005_s 0.00214577f $X=20.245 $Y=3.155 $X2=0 $Y2=0
cc_526 N_LVPWR_c_396_n N_X_M1011_s 0.00273098f $X=20.245 $Y=3.155 $X2=0 $Y2=0
cc_527 N_LVPWR_c_396_n N_X_c_1927_n 0.0355586f $X=20.245 $Y=3.155 $X2=0.24
+ $Y2=8.14
cc_528 N_LVPWR_c_396_n X 0.0377231f $X=20.245 $Y=3.155 $X2=24.72 $Y2=8.14
cc_529 N_LVPWR_c_396_n N_VPWR_M1005_d 0.0022433f $X=20.245 $Y=3.155 $X2=0 $Y2=0
cc_530 N_LVPWR_c_396_n N_VPWR_M1036_d 0.00165809f $X=20.245 $Y=3.155 $X2=0 $Y2=0
cc_531 N_LVPWR_c_396_n N_VPWR_M39_noxref_d 0.00216162f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_532 N_LVPWR_c_396_n N_VPWR_M43_noxref_s 0.0019895f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_533 N_LVPWR_c_396_n N_VPWR_M44_noxref_d 0.00253209f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_534 N_LVPWR_c_396_n N_VPWR_M46_noxref_d 0.0019895f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_535 N_LVPWR_c_396_n N_VPWR_c_1988_n 0.0365879f $X=20.245 $Y=3.155 $X2=0 $Y2=0
cc_536 N_LVPWR_c_396_n N_VPWR_c_1990_n 0.0345436f $X=20.245 $Y=3.155 $X2=0 $Y2=0
cc_537 N_LVPWR_c_396_n N_VPWR_c_1993_n 0.0365879f $X=20.245 $Y=3.155 $X2=0 $Y2=0
cc_538 N_LVPWR_c_396_n N_VPWR_c_1994_n 0.0374775f $X=20.245 $Y=3.155 $X2=24.72
+ $Y2=0
cc_539 N_LVPWR_c_396_n N_VPWR_c_1999_n 0.0353458f $X=20.245 $Y=3.155 $X2=0 $Y2=0
cc_540 N_LVPWR_c_396_n N_VPWR_c_2002_n 0.0374775f $X=20.245 $Y=3.155 $X2=0 $Y2=0
cc_541 N_LVPWR_c_396_n N_VPWR_c_2008_n 0.00480463f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_542 N_LVPWR_c_396_n N_VPWR_c_2013_n 0.00368087f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_543 N_LVPWR_c_396_n N_VPWR_c_2015_n 0.00481449f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_544 N_LVPWR_c_396_n N_VPWR_c_2016_n 0.00368087f $X=20.245 $Y=3.155 $X2=0
+ $Y2=0
cc_545 N_LVPWR_M1006_b N_VPWR_c_1981_n 0.0487138f $X=17.395 $Y=2.045 $X2=0 $Y2=0
cc_546 N_LVPWR_c_398_n N_VPWR_c_1981_n 0.0150761f $X=19.665 $Y=4.07 $X2=0 $Y2=0
cc_547 N_LVPWR_c_431_p N_VPWR_c_1981_n 0.0106548f $X=17.98 $Y=2.5 $X2=0 $Y2=0
cc_548 N_LVPWR_c_401_n N_VPWR_c_1981_n 0.029248f $X=18.795 $Y=3.62 $X2=0 $Y2=0
cc_549 N_LVPWR_c_402_n N_VPWR_c_1981_n 0.00982503f $X=18.065 $Y=3.62 $X2=0 $Y2=0
cc_550 N_LVPWR_c_435_p N_VPWR_c_1981_n 0.00997577f $X=18.88 $Y=2.84 $X2=0 $Y2=0
cc_551 N_LVPWR_c_404_n N_VPWR_c_1981_n 0.027788f $X=19.665 $Y=3.62 $X2=0 $Y2=0
cc_552 N_LVPWR_c_405_n N_VPWR_c_1981_n 0.0701049f $X=20.042 $Y=4.605 $X2=0 $Y2=0
cc_553 N_LVPWR_c_566_p N_VPWR_c_1981_n 0.00432131f $X=18.88 $Y=3.62 $X2=0 $Y2=0
cc_554 N_LVPWR_c_396_n N_VPWR_c_1981_n 2.60464f $X=20.245 $Y=3.155 $X2=0 $Y2=0
cc_555 N_LVPWR_M1006_b N_VPWR_c_1982_n 0.0704607f $X=17.395 $Y=2.045 $X2=0 $Y2=0
cc_556 N_LVPWR_c_453_p N_VPWR_c_1982_n 0.0215789f $X=17.95 $Y=4.94 $X2=0 $Y2=0
cc_557 N_LVPWR_c_398_n N_VPWR_c_1982_n 0.0145956f $X=19.665 $Y=4.07 $X2=0 $Y2=0
cc_558 N_LVPWR_c_399_n N_VPWR_c_1982_n 0.029248f $X=18.765 $Y=4.52 $X2=0 $Y2=0
cc_559 N_LVPWR_c_400_n N_VPWR_c_1982_n 0.00986368f $X=18.035 $Y=4.52 $X2=0 $Y2=0
cc_560 N_LVPWR_c_457_p N_VPWR_c_1982_n 0.0174306f $X=18.85 $Y=4.94 $X2=0 $Y2=0
cc_561 N_LVPWR_c_403_n N_VPWR_c_1982_n 0.029248f $X=19.665 $Y=4.52 $X2=0 $Y2=0
cc_562 N_LVPWR_c_405_n N_VPWR_c_1982_n 0.0401349f $X=20.042 $Y=4.605 $X2=0 $Y2=0
cc_563 N_LVPWR_c_463_p N_VPWR_c_1982_n 0.056449f $X=19.75 $Y=4.94 $X2=0 $Y2=0
cc_564 N_LVPWR_c_406_n N_VPWR_c_1982_n 0.0584025f $X=21.07 $Y=4.52 $X2=0 $Y2=0
cc_565 N_LVPWR_c_471_p N_VPWR_c_1982_n 0.0275033f $X=21.235 $Y=4.94 $X2=0 $Y2=0
cc_566 N_LVPWR_c_579_p N_VPWR_c_1982_n 0.00433346f $X=18.85 $Y=4.52 $X2=0 $Y2=0
cc_567 N_LVPWR_c_396_n N_A_1410_571#_M1022_d 8.01616e-19 $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_568 N_LVPWR_c_396_n N_A_1410_571#_M43_noxref_d 0.00273098f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_569 N_LVPWR_c_396_n N_A_1410_571#_M45_noxref_d 0.00273098f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_570 N_LVPWR_c_396_n N_A_1410_571#_c_2253_n 0.0204136f $X=20.245 $Y=3.155
+ $X2=0 $Y2=8.025
cc_571 N_LVPWR_c_396_n N_A_1410_571#_c_2254_n 0.00101656f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_572 N_LVPWR_c_396_n N_A_1410_571#_c_2257_n 0.0356241f $X=20.245 $Y=3.155
+ $X2=24.72 $Y2=0
cc_573 N_LVPWR_c_396_n N_A_1410_571#_c_2260_n 0.0356241f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_574 N_LVPWR_c_396_n N_A_1410_571#_c_2262_n 0.0123567f $X=20.245 $Y=3.155
+ $X2=0 $Y2=0
cc_575 N_LVPWR_c_396_n N_A_1410_571#_c_2263_n 0.0125804f $X=20.245 $Y=3.155
+ $X2=10.215 $Y2=0
cc_576 N_VGND_c_597_n N_A_262_107#_M1008_g 0.00289338f $X=1.95 $Y=0.81 $X2=0
+ $Y2=0
cc_577 N_VGND_c_680_n N_A_262_107#_M1008_g 0.0323575f $X=19.825 $Y=0.51 $X2=0
+ $Y2=0
cc_578 N_VGND_M1000_g N_A_262_107#_M1005_g 0.0179771f $X=1.56 $Y=6.425 $X2=0
+ $Y2=0
cc_579 N_VGND_c_597_n N_A_262_107#_c_842_n 7.39577e-19 $X=1.95 $Y=0.81 $X2=0
+ $Y2=0
cc_580 N_VGND_c_597_n N_A_262_107#_M1030_g 0.00289338f $X=1.95 $Y=0.81 $X2=0
+ $Y2=0
cc_581 N_VGND_c_674_n N_A_262_107#_M1030_g 0.0126165f $X=2.31 $Y=0.37 $X2=0
+ $Y2=0
cc_582 N_VGND_c_680_n N_A_262_107#_M1030_g 0.0306279f $X=19.825 $Y=0.51 $X2=0
+ $Y2=0
cc_583 N_VGND_c_602_n N_A_262_107#_M1047_g 0.00510247f $X=3.51 $Y=0.81 $X2=24.72
+ $Y2=8.14
cc_584 N_VGND_c_676_n N_A_262_107#_M1047_g 0.0126165f $X=3.395 $Y=0.37 $X2=24.72
+ $Y2=8.14
cc_585 N_VGND_c_680_n N_A_262_107#_M1047_g 0.0315672f $X=19.825 $Y=0.51
+ $X2=24.72 $Y2=8.14
cc_586 N_VGND_c_602_n N_A_262_107#_c_850_n 0.0148068f $X=3.51 $Y=0.81 $X2=12.48
+ $Y2=0
cc_587 N_VGND_c_602_n N_A_262_107#_c_851_n 0.0050964f $X=3.51 $Y=0.81 $X2=0.24
+ $Y2=8.14
cc_588 N_VGND_c_602_n N_A_262_107#_c_852_n 0.0475789f $X=3.51 $Y=0.81 $X2=12.48
+ $Y2=8.14
cc_589 N_VGND_c_603_n N_A_262_107#_c_852_n 6.48091e-19 $X=4.84 $Y=0.81 $X2=12.48
+ $Y2=8.14
cc_590 N_VGND_c_680_n N_A_262_107#_c_852_n 0.00998275f $X=19.825 $Y=0.51
+ $X2=12.48 $Y2=8.14
cc_591 N_VGND_c_603_n N_A_262_107#_c_853_n 0.0110199f $X=4.84 $Y=0.81 $X2=0
+ $Y2=0
cc_592 N_VGND_c_603_n N_A_262_107#_c_854_n 6.48091e-19 $X=4.84 $Y=0.81 $X2=0
+ $Y2=0
cc_593 N_VGND_c_680_n N_A_262_107#_c_854_n 0.00998275f $X=19.825 $Y=0.51 $X2=0
+ $Y2=0
cc_594 N_VGND_c_602_n N_A_840_107#_M1012_g 0.00392115f $X=3.51 $Y=0.81 $X2=0
+ $Y2=0
cc_595 N_VGND_c_603_n N_A_840_107#_M1012_g 0.00289338f $X=4.84 $Y=0.81 $X2=0
+ $Y2=0
cc_596 N_VGND_c_678_n N_A_840_107#_M1012_g 0.00583748f $X=5.02 $Y=0.37 $X2=0
+ $Y2=0
cc_597 N_VGND_c_680_n N_A_840_107#_M1012_g 0.0319624f $X=19.825 $Y=0.51 $X2=0
+ $Y2=0
cc_598 N_VGND_c_603_n N_A_840_107#_c_968_n 0.00203706f $X=4.84 $Y=0.81 $X2=0
+ $Y2=0
cc_599 N_VGND_c_603_n N_A_840_107#_M1034_g 0.00289338f $X=4.84 $Y=0.81 $X2=0
+ $Y2=0
cc_600 N_VGND_c_678_n N_A_840_107#_M1034_g 0.00583748f $X=5.02 $Y=0.37 $X2=0
+ $Y2=0
cc_601 N_VGND_c_680_n N_A_840_107#_M1034_g 0.0319624f $X=19.825 $Y=0.51 $X2=0
+ $Y2=0
cc_602 N_VGND_c_652_n N_A_840_107#_c_975_n 0.00620865f $X=9.47 $Y=7.685 $X2=0
+ $Y2=0
cc_603 N_VGND_c_682_n N_A_840_107#_c_975_n 0.00641183f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_604 N_VGND_c_606_n N_A_840_107#_c_976_n 0.0147574f $X=9.58 $Y=6.36 $X2=0
+ $Y2=0
cc_605 N_VGND_c_656_n N_A_840_107#_c_978_n 0.00620865f $X=11.83 $Y=7.685 $X2=0
+ $Y2=0
cc_606 N_VGND_c_682_n N_A_840_107#_c_978_n 0.00641183f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_607 N_VGND_c_607_n N_A_840_107#_c_979_n 0.0156327f $X=11.94 $Y=6.36 $X2=0
+ $Y2=0
cc_608 N_VGND_c_607_n N_A_840_107#_c_980_n 0.0111833f $X=11.94 $Y=6.36 $X2=0
+ $Y2=0
cc_609 N_VGND_c_608_n N_A_840_107#_c_980_n 6.41575e-19 $X=13.445 $Y=6.36 $X2=0
+ $Y2=0
cc_610 N_VGND_M1000_g N_A_362_1243#_c_1123_n 0.00589085f $X=1.56 $Y=6.425 $X2=0
+ $Y2=0
cc_611 N_VGND_c_590_n N_A_362_1243#_c_1123_n 6.41575e-19 $X=1.17 $Y=6.36 $X2=0
+ $Y2=0
cc_612 N_VGND_c_598_n N_A_362_1243#_c_1123_n 0.0169795f $X=2.5 $Y=6.36 $X2=0
+ $Y2=0
cc_613 N_VGND_c_598_n N_A_362_1243#_c_1124_n 0.0159914f $X=2.5 $Y=6.36 $X2=24.72
+ $Y2=0
cc_614 N_VGND_c_644_n N_A_362_1243#_c_1126_n 0.00620865f $X=4.75 $Y=7.685 $X2=0
+ $Y2=0
cc_615 N_VGND_c_682_n N_A_362_1243#_c_1126_n 0.00641183f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_616 N_VGND_c_604_n N_A_362_1243#_c_1127_n 0.0147574f $X=4.86 $Y=6.36 $X2=0
+ $Y2=0
cc_617 N_VGND_c_648_n N_A_362_1243#_c_1128_n 0.00620865f $X=7.11 $Y=7.685
+ $X2=24.72 $Y2=8.14
cc_618 N_VGND_c_682_n N_A_362_1243#_c_1128_n 0.00641183f $X=21.265 $Y=7.63
+ $X2=24.72 $Y2=8.14
cc_619 N_VGND_c_608_n N_A_2092_381#_M1002_g 0.00888967f $X=13.445 $Y=6.36 $X2=0
+ $Y2=0
cc_620 N_VGND_c_608_n N_A_2092_381#_c_1233_n 0.00905009f $X=13.445 $Y=6.36 $X2=0
+ $Y2=0
cc_621 N_VGND_c_608_n N_A_2092_381#_c_1216_n 0.00427281f $X=13.445 $Y=6.36 $X2=0
+ $Y2=0
cc_622 N_VGND_c_608_n N_A_2092_381#_c_1217_n 0.0314858f $X=13.445 $Y=6.36
+ $X2=10.215 $Y2=8.14
cc_623 N_VGND_c_609_n N_A_2092_381#_c_1217_n 6.41575e-19 $X=14.775 $Y=6.36
+ $X2=10.215 $Y2=8.14
cc_624 N_VGND_c_605_n N_A_1472_1171#_M1001_g 0.00495835f $X=7.22 $Y=6.36 $X2=0
+ $Y2=0
cc_625 N_VGND_c_652_n N_A_1472_1171#_M1001_g 0.0333719f $X=9.47 $Y=7.685 $X2=0
+ $Y2=0
cc_626 N_VGND_c_682_n N_A_1472_1171#_M1001_g 0.0288803f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_627 N_VGND_c_606_n N_A_1472_1171#_M1029_g 0.00495835f $X=9.58 $Y=6.36 $X2=0
+ $Y2=0
cc_628 N_VGND_c_652_n N_A_1472_1171#_M1029_g 0.0333719f $X=9.47 $Y=7.685 $X2=0
+ $Y2=0
cc_629 N_VGND_c_682_n N_A_1472_1171#_M1029_g 0.0288803f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_630 N_VGND_c_606_n N_A_1472_1171#_c_1318_n 0.00227604f $X=9.58 $Y=6.36 $X2=0
+ $Y2=0
cc_631 N_VGND_c_606_n N_A_1472_1171#_M1032_g 0.00495835f $X=9.58 $Y=6.36 $X2=0
+ $Y2=0
cc_632 N_VGND_c_656_n N_A_1472_1171#_M1032_g 0.0333719f $X=11.83 $Y=7.685 $X2=0
+ $Y2=0
cc_633 N_VGND_c_682_n N_A_1472_1171#_M1032_g 0.0288803f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_634 N_VGND_c_607_n N_A_1472_1171#_M1041_g 0.00888603f $X=11.94 $Y=6.36 $X2=0
+ $Y2=0
cc_635 N_VGND_c_656_n N_A_1472_1171#_M1041_g 0.0333719f $X=11.83 $Y=7.685 $X2=0
+ $Y2=0
cc_636 N_VGND_c_682_n N_A_1472_1171#_M1041_g 0.0288803f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_637 N_VGND_M1007_d N_A_1472_1171#_c_1325_n 0.00350673f $X=17.8 $Y=0.755 $X2=0
+ $Y2=0
cc_638 N_VGND_c_612_n N_A_1472_1171#_c_1325_n 0.0229947f $X=17.945 $Y=0.9 $X2=0
+ $Y2=0
cc_639 N_VGND_c_616_n N_A_1472_1171#_c_1374_n 0.0163928f $X=18.71 $Y=0.51 $X2=0
+ $Y2=0
cc_640 N_VGND_c_680_n N_A_1472_1171#_c_1374_n 0.0076335f $X=19.825 $Y=0.51 $X2=0
+ $Y2=0
cc_641 N_VGND_M1009_d N_A_1472_1171#_c_1327_n 0.00229612f $X=18.735 $Y=0.755
+ $X2=0 $Y2=0
cc_642 N_VGND_c_621_n N_A_1472_1171#_c_1327_n 0.0194017f $X=18.875 $Y=0.98 $X2=0
+ $Y2=0
cc_643 N_VGND_c_624_n N_A_1472_1171#_c_1378_n 0.012069f $X=19.62 $Y=0.51 $X2=0
+ $Y2=0
cc_644 N_VGND_c_680_n N_A_1472_1171#_c_1378_n 0.00516602f $X=19.825 $Y=0.51
+ $X2=0 $Y2=0
cc_645 N_VGND_M1016_d N_A_1472_1171#_c_1328_n 0.00309016f $X=19.645 $Y=0.755
+ $X2=0 $Y2=0
cc_646 N_VGND_c_628_n N_A_1472_1171#_c_1328_n 0.0232152f $X=19.785 $Y=0.98 $X2=0
+ $Y2=0
cc_647 N_VGND_c_608_n N_SLEEP_B_M1045_g 0.00703514f $X=13.445 $Y=6.36 $X2=0
+ $Y2=0
cc_648 N_VGND_c_609_n N_SLEEP_B_M1045_g 0.00863053f $X=14.775 $Y=6.36 $X2=0
+ $Y2=0
cc_649 N_VGND_c_664_n N_SLEEP_B_M1045_g 0.0129076f $X=14.665 $Y=7.685 $X2=0
+ $Y2=0
cc_650 N_VGND_c_682_n N_SLEEP_B_M1045_g 0.0136096f $X=21.265 $Y=7.63 $X2=0 $Y2=0
cc_651 N_VGND_c_609_n N_SLEEP_B_c_1469_n 0.00465036f $X=14.775 $Y=6.36 $X2=0
+ $Y2=0
cc_652 N_VGND_c_609_n N_SLEEP_B_c_1470_n 0.0114872f $X=14.775 $Y=6.36 $X2=0
+ $Y2=0
cc_653 N_VGND_c_613_n N_A_3617_1198#_M1018_g 4.54744e-19 $X=17.945 $Y=7.515
+ $X2=-0.33 $Y2=-0.265
cc_654 N_VGND_c_615_n N_A_3617_1198#_M1018_g 0.0121142f $X=17.945 $Y=7.16
+ $X2=-0.33 $Y2=-0.265
cc_655 N_VGND_c_618_n N_A_3617_1198#_M1018_g 0.00512208f $X=18.69 $Y=7.63
+ $X2=-0.33 $Y2=-0.265
cc_656 N_VGND_c_682_n N_A_3617_1198#_M1018_g 0.00435847f $X=21.265 $Y=7.63
+ $X2=-0.33 $Y2=-0.265
cc_657 N_VGND_c_615_n N_A_3617_1198#_M1019_g 5.73449e-19 $X=17.945 $Y=7.16
+ $X2=0.24 $Y2=0
cc_658 N_VGND_c_618_n N_A_3617_1198#_M1019_g 0.00616943f $X=18.69 $Y=7.63
+ $X2=0.24 $Y2=0
cc_659 N_VGND_c_620_n N_A_3617_1198#_M1019_g 0.00233719f $X=18.855 $Y=7.16
+ $X2=0.24 $Y2=0
cc_660 N_VGND_c_682_n N_A_3617_1198#_M1019_g 0.00523016f $X=21.265 $Y=7.63
+ $X2=0.24 $Y2=0
cc_661 N_VGND_c_620_n N_A_3617_1198#_M1027_g 0.010436f $X=18.855 $Y=7.16
+ $X2=24.72 $Y2=0
cc_662 N_VGND_c_622_n N_A_3617_1198#_M1027_g 0.00512208f $X=19.62 $Y=7.63
+ $X2=24.72 $Y2=0
cc_663 N_VGND_c_666_n N_A_3617_1198#_M1027_g 4.54744e-19 $X=18.855 $Y=7.63
+ $X2=24.72 $Y2=0
cc_664 N_VGND_c_682_n N_A_3617_1198#_M1027_g 0.00435847f $X=21.265 $Y=7.63
+ $X2=24.72 $Y2=0
cc_665 N_VGND_c_620_n N_A_3617_1198#_M1033_g 5.66437e-19 $X=18.855 $Y=7.16 $X2=0
+ $Y2=0
cc_666 N_VGND_c_622_n N_A_3617_1198#_M1033_g 0.00616943f $X=19.62 $Y=7.63 $X2=0
+ $Y2=0
cc_667 N_VGND_c_629_n N_A_3617_1198#_M1033_g 0.00565513f $X=19.785 $Y=6.79 $X2=0
+ $Y2=0
cc_668 N_VGND_c_682_n N_A_3617_1198#_M1033_g 0.00523016f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_669 N_VGND_c_629_n N_A_3617_1198#_c_1500_n 0.0245688f $X=19.785 $Y=6.79
+ $X2=24.72 $Y2=8.14
cc_670 N_VGND_c_632_n N_A_3617_1198#_c_1501_n 0.0177842f $X=20.35 $Y=6.79
+ $X2=12.48 $Y2=0
cc_671 N_VGND_c_632_n N_A_3617_1198#_c_1503_n 0.0264979f $X=20.35 $Y=6.79 $X2=0
+ $Y2=0
cc_672 N_VGND_c_633_n N_A_3617_1198#_c_1503_n 0.0193811f $X=21.125 $Y=7.63 $X2=0
+ $Y2=0
cc_673 N_VGND_c_637_n N_A_3617_1198#_c_1503_n 0.0264979f $X=21.21 $Y=6.79 $X2=0
+ $Y2=0
cc_674 N_VGND_c_682_n N_A_3617_1198#_c_1503_n 0.00987443f $X=21.265 $Y=7.63
+ $X2=0 $Y2=0
cc_675 N_VGND_c_598_n N_A_528_1171#_M1004_g 9.46322e-19 $X=2.5 $Y=6.36 $X2=0
+ $Y2=0
cc_676 N_VGND_c_599_n N_A_528_1171#_M1004_g 0.00786538f $X=2.47 $Y=7.57 $X2=0
+ $Y2=0
cc_677 N_VGND_c_644_n N_A_528_1171#_M1004_g 0.0333719f $X=4.75 $Y=7.685 $X2=0
+ $Y2=0
cc_678 N_VGND_c_682_n N_A_528_1171#_M1004_g 0.0288803f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_679 N_VGND_c_604_n N_A_528_1171#_M1010_g 0.00495835f $X=4.86 $Y=6.36 $X2=0
+ $Y2=0
cc_680 N_VGND_c_644_n N_A_528_1171#_M1010_g 0.0333719f $X=4.75 $Y=7.685 $X2=0
+ $Y2=0
cc_681 N_VGND_c_682_n N_A_528_1171#_M1010_g 0.0288803f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_682 N_VGND_c_604_n N_A_528_1171#_c_1616_n 0.00227604f $X=4.86 $Y=6.36
+ $X2=24.72 $Y2=0
cc_683 N_VGND_c_604_n N_A_528_1171#_M1023_g 0.00495835f $X=4.86 $Y=6.36 $X2=0
+ $Y2=0
cc_684 N_VGND_c_648_n N_A_528_1171#_M1023_g 0.0333719f $X=7.11 $Y=7.685 $X2=0
+ $Y2=0
cc_685 N_VGND_c_682_n N_A_528_1171#_M1023_g 0.0288803f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_686 N_VGND_c_605_n N_A_528_1171#_M1040_g 0.00495835f $X=7.22 $Y=6.36 $X2=0
+ $Y2=0
cc_687 N_VGND_c_648_n N_A_528_1171#_M1040_g 0.0333719f $X=7.11 $Y=7.685 $X2=0
+ $Y2=0
cc_688 N_VGND_c_682_n N_A_528_1171#_M1040_g 0.0288803f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_689 N_VGND_c_605_n N_A_528_1171#_c_1646_n 0.00619614f $X=7.22 $Y=6.36 $X2=0
+ $Y2=0
cc_690 N_VGND_c_612_n N_A_528_1171#_c_1622_n 0.00740132f $X=17.945 $Y=0.9
+ $X2=10.215 $Y2=0
cc_691 N_VGND_c_680_n N_A_528_1171#_c_1623_n 0.229481f $X=19.825 $Y=0.51
+ $X2=10.215 $Y2=0
cc_692 N_VGND_c_612_n N_A_528_1171#_M1007_g 0.00452505f $X=17.945 $Y=0.9
+ $X2=10.215 $Y2=8.14
cc_693 N_VGND_c_616_n N_A_528_1171#_M1007_g 0.00616943f $X=18.71 $Y=0.51
+ $X2=10.215 $Y2=8.14
cc_694 N_VGND_c_621_n N_A_528_1171#_M1007_g 5.66437e-19 $X=18.875 $Y=0.98
+ $X2=10.215 $Y2=8.14
cc_695 N_VGND_c_680_n N_A_528_1171#_M1007_g 0.00523016f $X=19.825 $Y=0.51
+ $X2=10.215 $Y2=8.14
cc_696 N_VGND_c_616_n N_A_528_1171#_M1009_g 0.00512208f $X=18.71 $Y=0.51 $X2=0
+ $Y2=0
cc_697 N_VGND_c_621_n N_A_528_1171#_M1009_g 0.010436f $X=18.875 $Y=0.98 $X2=0
+ $Y2=0
cc_698 N_VGND_c_668_n N_A_528_1171#_M1009_g 4.54744e-19 $X=18.875 $Y=0.51 $X2=0
+ $Y2=0
cc_699 N_VGND_c_680_n N_A_528_1171#_M1009_g 0.00435847f $X=19.825 $Y=0.51 $X2=0
+ $Y2=0
cc_700 N_VGND_c_621_n N_A_528_1171#_M1014_g 0.00233719f $X=18.875 $Y=0.98 $X2=0
+ $Y2=0
cc_701 N_VGND_c_624_n N_A_528_1171#_M1014_g 0.00616943f $X=19.62 $Y=0.51 $X2=0
+ $Y2=0
cc_702 N_VGND_c_628_n N_A_528_1171#_M1014_g 5.73449e-19 $X=19.785 $Y=0.98 $X2=0
+ $Y2=0
cc_703 N_VGND_c_680_n N_A_528_1171#_M1014_g 0.00523016f $X=19.825 $Y=0.51 $X2=0
+ $Y2=0
cc_704 N_VGND_c_624_n N_A_528_1171#_M1016_g 0.00512208f $X=19.62 $Y=0.51 $X2=0
+ $Y2=0
cc_705 N_VGND_c_626_n N_A_528_1171#_M1016_g 4.54744e-19 $X=19.785 $Y=0.625 $X2=0
+ $Y2=0
cc_706 N_VGND_c_628_n N_A_528_1171#_M1016_g 0.0121142f $X=19.785 $Y=0.98 $X2=0
+ $Y2=0
cc_707 N_VGND_c_680_n N_A_528_1171#_M1016_g 0.00435847f $X=19.825 $Y=0.51 $X2=0
+ $Y2=0
cc_708 N_VGND_c_615_n N_A_528_1171#_c_1640_n 0.0024426f $X=17.945 $Y=7.16 $X2=0
+ $Y2=0
cc_709 N_VGND_M1018_d N_A_528_1171#_c_1641_n 0.00301575f $X=17.8 $Y=6.645 $X2=0
+ $Y2=0
cc_710 N_VGND_c_615_n N_A_528_1171#_c_1641_n 0.0207726f $X=17.945 $Y=7.16 $X2=0
+ $Y2=0
cc_711 N_VGND_c_618_n N_A_528_1171#_c_1736_n 0.012069f $X=18.69 $Y=7.63 $X2=0
+ $Y2=0
cc_712 N_VGND_c_682_n N_A_528_1171#_c_1736_n 0.00516602f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_713 N_VGND_M1019_d N_A_528_1171#_c_1642_n 0.00229612f $X=18.665 $Y=6.645
+ $X2=0 $Y2=0
cc_714 N_VGND_c_620_n N_A_528_1171#_c_1642_n 0.0194017f $X=18.855 $Y=7.16 $X2=0
+ $Y2=0
cc_715 N_VGND_c_629_n N_A_528_1171#_c_1642_n 0.00167954f $X=19.785 $Y=6.79 $X2=0
+ $Y2=0
cc_716 N_VGND_c_622_n N_A_528_1171#_c_1741_n 0.0163928f $X=19.62 $Y=7.63 $X2=0
+ $Y2=0
cc_717 N_VGND_c_682_n N_A_528_1171#_c_1741_n 0.0076335f $X=21.265 $Y=7.63 $X2=0
+ $Y2=0
cc_718 N_VGND_c_632_n N_A_M1024_g 0.00683317f $X=20.35 $Y=6.79 $X2=0 $Y2=0
cc_719 N_VGND_c_633_n N_A_M1024_g 0.00577902f $X=21.125 $Y=7.63 $X2=0 $Y2=0
cc_720 N_VGND_c_682_n N_A_M1024_g 0.00523016f $X=21.265 $Y=7.63 $X2=0 $Y2=0
cc_721 N_VGND_c_637_n N_A_c_1870_n 0.00196285f $X=21.21 $Y=6.79 $X2=0 $Y2=8.025
cc_722 N_VGND_c_633_n N_A_M1046_g 0.00577902f $X=21.125 $Y=7.63 $X2=0 $Y2=0
cc_723 N_VGND_c_637_n N_A_M1046_g 0.00683317f $X=21.21 $Y=6.79 $X2=0 $Y2=0
cc_724 N_VGND_c_682_n N_A_M1046_g 0.00523016f $X=21.265 $Y=7.63 $X2=0 $Y2=0
cc_725 N_VGND_c_637_n A 0.0215684f $X=21.21 $Y=6.79 $X2=0 $Y2=0
cc_726 N_VGND_c_597_n N_X_c_1920_n 6.48091e-19 $X=1.95 $Y=0.81 $X2=0 $Y2=0
cc_727 N_VGND_c_680_n N_X_c_1920_n 0.00998275f $X=19.825 $Y=0.51 $X2=0 $Y2=0
cc_728 N_VGND_c_597_n N_X_c_1921_n 0.011937f $X=1.95 $Y=0.81 $X2=0 $Y2=0
cc_729 N_VGND_c_597_n N_X_c_1922_n 6.48091e-19 $X=1.95 $Y=0.81 $X2=24.72 $Y2=0
cc_730 N_VGND_c_602_n N_X_c_1922_n 6.48091e-19 $X=3.51 $Y=0.81 $X2=24.72 $Y2=0
cc_731 N_VGND_c_680_n N_X_c_1922_n 0.00998275f $X=19.825 $Y=0.51 $X2=24.72 $Y2=0
cc_732 N_A_262_107#_c_851_n N_A_840_107#_M1012_g 0.00591016f $X=3.515 $Y=2.03
+ $X2=0 $Y2=0
cc_733 N_A_262_107#_c_852_n N_A_840_107#_M1012_g 0.010109f $X=4.06 $Y=0.81 $X2=0
+ $Y2=0
cc_734 N_A_262_107#_c_855_n N_A_840_107#_M1012_g 0.00208822f $X=4.06 $Y=2.03
+ $X2=0 $Y2=0
cc_735 N_A_262_107#_c_868_n N_A_840_107#_M39_noxref_g 0.0127377f $X=4.06 $Y=2.57
+ $X2=0 $Y2=0
cc_736 N_A_262_107#_c_853_n N_A_840_107#_M39_noxref_g 0.0249504f $X=5.51 $Y=2.03
+ $X2=0 $Y2=0
cc_737 N_A_262_107#_c_855_n N_A_840_107#_M39_noxref_g 0.00208952f $X=4.06
+ $Y=2.03 $X2=0 $Y2=0
cc_738 N_A_262_107#_c_853_n N_A_840_107#_c_968_n 0.0116766f $X=5.51 $Y=2.03
+ $X2=0 $Y2=0
cc_739 N_A_262_107#_c_854_n N_A_840_107#_M1034_g 0.0122356f $X=5.62 $Y=0.81
+ $X2=0 $Y2=0
cc_740 N_A_262_107#_c_853_n N_A_840_107#_M40_noxref_g 0.0247919f $X=5.51 $Y=2.03
+ $X2=0.24 $Y2=8.14
cc_741 N_A_262_107#_c_871_n N_A_840_107#_M40_noxref_g 0.00989074f $X=5.62
+ $Y=2.57 $X2=0.24 $Y2=8.14
cc_742 N_A_262_107#_c_853_n N_A_840_107#_c_971_n 0.00155418f $X=5.51 $Y=2.03
+ $X2=0 $Y2=0
cc_743 N_A_262_107#_c_854_n N_A_840_107#_c_971_n 0.00631677f $X=5.62 $Y=0.81
+ $X2=0 $Y2=0
cc_744 N_A_262_107#_c_874_n N_A_840_107#_c_971_n 0.0169051f $X=5.62 $Y=2.03
+ $X2=0 $Y2=0
cc_745 N_A_262_107#_c_871_n N_A_840_107#_c_988_n 0.0175346f $X=5.62 $Y=2.57
+ $X2=24.72 $Y2=8.14
cc_746 N_A_262_107#_c_874_n N_A_840_107#_c_988_n 8.61763e-19 $X=5.62 $Y=2.03
+ $X2=24.72 $Y2=8.14
cc_747 N_A_262_107#_c_853_n N_A_840_107#_c_972_n 0.0351651f $X=5.51 $Y=2.03
+ $X2=10.215 $Y2=0
cc_748 N_A_262_107#_c_853_n N_A_840_107#_c_973_n 0.0316835f $X=5.51 $Y=2.03
+ $X2=10.215 $Y2=0
cc_749 N_A_262_107#_M1011_g N_A_362_1243#_c_1124_n 0.0206068f $X=2.34 $Y=3.925
+ $X2=24.72 $Y2=0
cc_750 N_A_262_107#_M1036_g N_A_362_1243#_c_1124_n 0.0113045f $X=3.12 $Y=3.925
+ $X2=24.72 $Y2=0
cc_751 N_A_262_107#_c_871_n N_A_362_1243#_c_1129_n 0.0296347f $X=5.62 $Y=2.57
+ $X2=10.215 $Y2=0
cc_752 N_A_262_107#_c_871_n N_A_362_1243#_c_1138_n 0.0119787f $X=5.62 $Y=2.57
+ $X2=24.72 $Y2=0
cc_753 N_A_262_107#_M1036_g N_A_528_1171#_c_1614_n 0.0209968f $X=3.12 $Y=3.925
+ $X2=0 $Y2=0
cc_754 N_A_262_107#_M1008_g N_X_c_1920_n 0.0127137f $X=1.56 $Y=1.165 $X2=0 $Y2=0
cc_755 N_A_262_107#_M1008_g N_X_c_1921_n 0.0234116f $X=1.56 $Y=1.165 $X2=0 $Y2=0
cc_756 N_A_262_107#_M1005_g N_X_c_1921_n 0.0234116f $X=1.56 $Y=3.925 $X2=0 $Y2=0
cc_757 N_A_262_107#_c_842_n N_X_c_1921_n 0.00802808f $X=2.09 $Y=2.03 $X2=0 $Y2=0
cc_758 N_A_262_107#_M1030_g N_X_c_1921_n 0.0233336f $X=2.34 $Y=1.165 $X2=0 $Y2=0
cc_759 N_A_262_107#_M1011_g N_X_c_1921_n 0.0233336f $X=2.34 $Y=3.925 $X2=0 $Y2=0
cc_760 N_A_262_107#_c_845_n N_X_c_1921_n 5.27321e-19 $X=2.87 $Y=2.03 $X2=0 $Y2=0
cc_761 N_A_262_107#_c_848_n N_X_c_1921_n 0.0132772f $X=1.56 $Y=2.03 $X2=0 $Y2=0
cc_762 N_A_262_107#_c_849_n N_X_c_1921_n 0.00941644f $X=2.34 $Y=2.03 $X2=0 $Y2=0
cc_763 N_A_262_107#_M1030_g N_X_c_1922_n 0.007192f $X=2.34 $Y=1.165 $X2=24.72
+ $Y2=0
cc_764 N_A_262_107#_M1047_g N_X_c_1922_n 0.00624147f $X=3.12 $Y=1.165 $X2=24.72
+ $Y2=0
cc_765 N_A_262_107#_c_850_n N_X_c_1922_n 0.00435706f $X=3.95 $Y=2.03 $X2=24.72
+ $Y2=0
cc_766 N_A_262_107#_M1011_g N_X_c_1927_n 0.0117782f $X=2.34 $Y=3.925 $X2=0.24
+ $Y2=8.14
cc_767 N_A_262_107#_c_850_n N_X_c_1927_n 0.00435706f $X=3.95 $Y=2.03 $X2=0.24
+ $Y2=8.14
cc_768 N_A_262_107#_c_851_n N_X_c_1927_n 0.0108276f $X=3.515 $Y=2.03 $X2=0.24
+ $Y2=8.14
cc_769 N_A_262_107#_c_845_n N_X_c_1958_n 0.0118894f $X=2.87 $Y=2.03 $X2=0 $Y2=0
cc_770 N_A_262_107#_c_850_n N_X_c_1958_n 0.018713f $X=3.95 $Y=2.03 $X2=0 $Y2=0
cc_771 N_A_262_107#_c_851_n N_X_c_1958_n 2.08086e-19 $X=3.515 $Y=2.03 $X2=0
+ $Y2=0
cc_772 N_A_262_107#_M1005_g X 0.0175006f $X=1.56 $Y=3.925 $X2=24.72 $Y2=8.14
cc_773 N_A_262_107#_M1005_g N_VPWR_c_1988_n 0.00377453f $X=1.56 $Y=3.925 $X2=0
+ $Y2=0
cc_774 N_A_262_107#_c_842_n N_VPWR_c_1988_n 7.39577e-19 $X=2.09 $Y=2.03 $X2=0
+ $Y2=0
cc_775 N_A_262_107#_M1011_g N_VPWR_c_1988_n 0.00377453f $X=2.34 $Y=3.925 $X2=0
+ $Y2=0
cc_776 N_A_262_107#_M1036_g N_VPWR_c_1990_n 0.00417775f $X=3.12 $Y=3.925 $X2=0
+ $Y2=0
cc_777 N_A_262_107#_c_850_n N_VPWR_c_1990_n 0.0164123f $X=3.95 $Y=2.03 $X2=0
+ $Y2=0
cc_778 N_A_262_107#_c_851_n N_VPWR_c_1990_n 0.00520252f $X=3.515 $Y=2.03 $X2=0
+ $Y2=0
cc_779 N_A_262_107#_c_868_n N_VPWR_c_1990_n 0.0563495f $X=4.06 $Y=2.57 $X2=0
+ $Y2=0
cc_780 N_A_262_107#_c_868_n N_VPWR_c_1992_n 0.00237952f $X=4.06 $Y=2.57 $X2=0
+ $Y2=0
cc_781 N_A_262_107#_c_868_n N_VPWR_c_1993_n 0.00410199f $X=4.06 $Y=2.57 $X2=0
+ $Y2=0
cc_782 N_A_262_107#_c_853_n N_VPWR_c_1993_n 0.0143702f $X=5.51 $Y=2.03 $X2=0
+ $Y2=0
cc_783 N_A_262_107#_c_871_n N_VPWR_c_1993_n 0.00410199f $X=5.62 $Y=2.57 $X2=0
+ $Y2=0
cc_784 N_A_262_107#_c_871_n N_VPWR_c_2008_n 0.0101728f $X=5.62 $Y=2.57 $X2=0
+ $Y2=0
cc_785 N_A_262_107#_M1005_g N_VPWR_c_2010_n 0.0138184f $X=1.56 $Y=3.925 $X2=0
+ $Y2=0
cc_786 N_A_262_107#_M1011_g N_VPWR_c_2010_n 0.0138184f $X=2.34 $Y=3.925 $X2=0
+ $Y2=0
cc_787 N_A_262_107#_M1036_g N_VPWR_c_2011_n 0.0138184f $X=3.12 $Y=3.925 $X2=0
+ $Y2=0
cc_788 N_A_262_107#_M39_noxref_s N_VPWR_c_1981_n 0.00250198f $X=3.935 $Y=2.425
+ $X2=0 $Y2=0
cc_789 N_A_262_107#_M40_noxref_d N_VPWR_c_1981_n 0.00250198f $X=5.48 $Y=2.425
+ $X2=0 $Y2=0
cc_790 N_A_262_107#_M1005_g N_VPWR_c_1981_n 0.0144881f $X=1.56 $Y=3.925 $X2=0
+ $Y2=0
cc_791 N_A_262_107#_M1011_g N_VPWR_c_1981_n 0.0144881f $X=2.34 $Y=3.925 $X2=0
+ $Y2=0
cc_792 N_A_262_107#_M1036_g N_VPWR_c_1981_n 0.0144881f $X=3.12 $Y=3.925 $X2=0
+ $Y2=0
cc_793 N_A_262_107#_c_868_n N_VPWR_c_1981_n 0.0271439f $X=4.06 $Y=2.57 $X2=0
+ $Y2=0
cc_794 N_A_262_107#_c_871_n N_VPWR_c_1981_n 0.0263521f $X=5.62 $Y=2.57 $X2=0
+ $Y2=0
cc_795 N_A_262_107#_M1005_g N_VPWR_c_1982_n 0.0297218f $X=1.56 $Y=3.925 $X2=0
+ $Y2=0
cc_796 N_A_262_107#_M1011_g N_VPWR_c_1982_n 0.0297218f $X=2.34 $Y=3.925 $X2=0
+ $Y2=0
cc_797 N_A_262_107#_M1036_g N_VPWR_c_1982_n 0.0297218f $X=3.12 $Y=3.925 $X2=0
+ $Y2=0
cc_798 N_A_840_107#_M1022_g N_A_362_1243#_M1043_g 0.0187199f $X=6.8 $Y=3.605
+ $X2=0 $Y2=0
cc_799 N_A_840_107#_c_997_n N_A_362_1243#_M1043_g 0.0079407f $X=7.97 $Y=3 $X2=0
+ $Y2=0
cc_800 N_A_840_107#_c_1001_n N_A_362_1243#_M1043_g 0.00246719f $X=7.87 $Y=5.07
+ $X2=0 $Y2=0
cc_801 N_A_840_107#_c_1002_n N_A_362_1243#_M1043_g 0.0161883f $X=7.87 $Y=5.07
+ $X2=0 $Y2=0
cc_802 N_A_840_107#_c_988_n N_A_362_1243#_c_1134_n 0.0200332f $X=6.015 $Y=4.905
+ $X2=0.24 $Y2=0
cc_803 N_A_840_107#_M1022_g N_A_362_1243#_c_1134_n 0.0356269f $X=6.8 $Y=3.605
+ $X2=0.24 $Y2=0
cc_804 N_A_840_107#_c_991_n N_A_362_1243#_c_1127_n 0.00339858f $X=6.115 $Y=5.07
+ $X2=0 $Y2=0
cc_805 N_A_840_107#_c_988_n N_A_362_1243#_c_1129_n 0.0383276f $X=6.015 $Y=4.905
+ $X2=10.215 $Y2=0
cc_806 N_A_840_107#_c_990_n N_A_362_1243#_c_1129_n 0.0436687f $X=6.55 $Y=5.07
+ $X2=10.215 $Y2=0
cc_807 N_A_840_107#_M1022_g N_A_362_1243#_c_1129_n 0.0227253f $X=6.8 $Y=3.605
+ $X2=10.215 $Y2=0
cc_808 N_A_840_107#_c_988_n N_A_362_1243#_c_1138_n 0.00367084f $X=6.015 $Y=4.905
+ $X2=24.72 $Y2=0
cc_809 N_A_840_107#_M1022_g N_A_362_1243#_c_1144_n 0.0034221f $X=6.8 $Y=3.605
+ $X2=0.24 $Y2=8.14
cc_810 N_A_840_107#_c_990_n N_A_362_1243#_c_1130_n 0.00354564f $X=6.55 $Y=5.07
+ $X2=24.72 $Y2=8.14
cc_811 N_A_840_107#_c_976_n N_A_2092_381#_c_1221_n 0.00206021f $X=10.65 $Y=5.865
+ $X2=0 $Y2=8.025
cc_812 N_A_840_107#_c_979_n N_A_2092_381#_c_1221_n 0.0338814f $X=12.555 $Y=5.865
+ $X2=0 $Y2=8.025
cc_813 N_A_840_107#_c_1003_n N_A_2092_381#_c_1221_n 0.00285952f $X=10.76
+ $Y=5.865 $X2=0 $Y2=8.025
cc_814 N_A_840_107#_c_979_n N_A_2092_381#_c_1227_n 0.00701338f $X=12.555
+ $Y=5.865 $X2=24.72 $Y2=0
cc_815 N_A_840_107#_c_979_n N_A_2092_381#_M1002_g 0.0118838f $X=12.555 $Y=5.865
+ $X2=0 $Y2=0
cc_816 N_A_840_107#_c_980_n N_A_2092_381#_M1002_g 0.0110787f $X=12.665 $Y=6.36
+ $X2=0 $Y2=0
cc_817 N_A_840_107#_c_975_n N_A_1472_1171#_M1001_g 0.00441776f $X=8.4 $Y=6.36
+ $X2=0 $Y2=0
cc_818 N_A_840_107#_c_975_n N_A_1472_1171#_c_1312_n 0.0120183f $X=8.4 $Y=6.36
+ $X2=0.24 $Y2=0
cc_819 N_A_840_107#_c_976_n N_A_1472_1171#_c_1312_n 0.00204387f $X=10.65
+ $Y=5.865 $X2=0.24 $Y2=0
cc_820 N_A_840_107#_c_977_n N_A_1472_1171#_c_1312_n 0.00645509f $X=8.51 $Y=5.865
+ $X2=0.24 $Y2=0
cc_821 N_A_840_107#_c_974_n N_A_1472_1171#_c_1313_n 2.3241e-19 $X=7.97 $Y=5.755
+ $X2=0 $Y2=0
cc_822 N_A_840_107#_c_977_n N_A_1472_1171#_c_1313_n 0.030241f $X=8.51 $Y=5.865
+ $X2=0 $Y2=0
cc_823 N_A_840_107#_c_975_n N_A_1472_1171#_M1029_g 0.00441776f $X=8.4 $Y=6.36
+ $X2=0 $Y2=0
cc_824 N_A_840_107#_c_974_n N_A_1472_1171#_c_1315_n 0.00300992f $X=7.97 $Y=5.755
+ $X2=0 $Y2=0
cc_825 N_A_840_107#_c_976_n N_A_1472_1171#_c_1315_n 0.0136339f $X=10.65 $Y=5.865
+ $X2=0 $Y2=0
cc_826 N_A_840_107#_c_976_n N_A_1472_1171#_c_1318_n 0.0130802f $X=10.65 $Y=5.865
+ $X2=0 $Y2=0
cc_827 N_A_840_107#_c_978_n N_A_1472_1171#_M1032_g 0.00441776f $X=10.76 $Y=6.36
+ $X2=0 $Y2=0
cc_828 N_A_840_107#_c_976_n N_A_1472_1171#_c_1320_n 0.00171059f $X=10.65
+ $Y=5.865 $X2=0 $Y2=0
cc_829 N_A_840_107#_c_978_n N_A_1472_1171#_c_1320_n 0.0112496f $X=10.76 $Y=6.36
+ $X2=0 $Y2=0
cc_830 N_A_840_107#_c_979_n N_A_1472_1171#_c_1320_n 0.0596852f $X=12.555
+ $Y=5.865 $X2=0 $Y2=0
cc_831 N_A_840_107#_c_1003_n N_A_1472_1171#_c_1320_n 0.0034419f $X=10.76
+ $Y=5.865 $X2=0 $Y2=0
cc_832 N_A_840_107#_c_978_n N_A_1472_1171#_M1041_g 0.00441776f $X=10.76 $Y=6.36
+ $X2=0 $Y2=0
cc_833 N_A_840_107#_c_976_n N_A_1472_1171#_c_1322_n 0.0624517f $X=10.65 $Y=5.865
+ $X2=0.24 $Y2=0
cc_834 N_A_840_107#_c_976_n N_A_1472_1171#_c_1323_n 0.0637912f $X=10.65 $Y=5.865
+ $X2=0 $Y2=0
cc_835 N_A_840_107#_c_991_n N_A_528_1171#_c_1618_n 0.00983382f $X=6.115 $Y=5.07
+ $X2=0.24 $Y2=8.14
cc_836 N_A_840_107#_c_974_n N_A_528_1171#_c_1646_n 0.0207015f $X=7.97 $Y=5.755
+ $X2=0 $Y2=0
cc_837 N_A_840_107#_c_977_n N_A_528_1171#_c_1646_n 0.0092082f $X=8.51 $Y=5.865
+ $X2=0 $Y2=0
cc_838 N_A_840_107#_c_1001_n N_A_528_1171#_c_1646_n 0.00351221f $X=7.87 $Y=5.07
+ $X2=0 $Y2=0
cc_839 N_A_840_107#_c_1002_n N_A_528_1171#_c_1646_n 0.0408941f $X=7.87 $Y=5.07
+ $X2=0 $Y2=0
cc_840 N_A_840_107#_c_996_n N_A_528_1171#_c_1647_n 0.0408941f $X=6.8 $Y=5.07
+ $X2=0 $Y2=0
cc_841 N_A_840_107#_c_997_n N_A_528_1171#_c_1621_n 0.0456725f $X=7.97 $Y=3 $X2=0
+ $Y2=0
cc_842 N_A_840_107#_c_974_n N_A_528_1171#_c_1621_n 0.0074946f $X=7.97 $Y=5.755
+ $X2=0 $Y2=0
cc_843 N_A_840_107#_c_1001_n N_A_528_1171#_c_1621_n 0.00873718f $X=7.87 $Y=5.07
+ $X2=0 $Y2=0
cc_844 N_A_840_107#_c_1002_n N_A_528_1171#_c_1621_n 0.0200332f $X=7.87 $Y=5.07
+ $X2=0 $Y2=0
cc_845 N_A_840_107#_c_990_n N_A_528_1171#_c_1633_n 0.00983382f $X=6.55 $Y=5.07
+ $X2=0 $Y2=0
cc_846 N_A_840_107#_M39_noxref_g N_VPWR_c_1990_n 0.00809852f $X=4.45 $Y=3.175
+ $X2=0 $Y2=0
cc_847 N_A_840_107#_M39_noxref_g N_VPWR_c_1993_n 0.00157749f $X=4.45 $Y=3.175
+ $X2=0 $Y2=0
cc_848 N_A_840_107#_c_968_n N_VPWR_c_1993_n 7.08729e-19 $X=4.98 $Y=2.01 $X2=0
+ $Y2=0
cc_849 N_A_840_107#_M40_noxref_g N_VPWR_c_1993_n 0.00157749f $X=5.23 $Y=3.175
+ $X2=0 $Y2=0
cc_850 N_A_840_107#_c_976_n N_VPWR_c_1997_n 0.00735061f $X=10.65 $Y=5.865 $X2=0
+ $Y2=0
cc_851 N_A_840_107#_c_979_n N_VPWR_c_1997_n 0.0308854f $X=12.555 $Y=5.865 $X2=0
+ $Y2=0
cc_852 N_A_840_107#_c_1003_n N_VPWR_c_1997_n 0.00803194f $X=10.76 $Y=5.865 $X2=0
+ $Y2=0
cc_853 N_A_840_107#_c_976_n N_VPWR_c_1998_n 0.00893992f $X=10.65 $Y=5.865 $X2=0
+ $Y2=0
cc_854 N_A_840_107#_c_979_n N_VPWR_c_2001_n 0.027759f $X=12.555 $Y=5.865 $X2=0
+ $Y2=0
cc_855 N_A_840_107#_c_979_n N_VPWR_c_2007_n 0.00888724f $X=12.555 $Y=5.865 $X2=0
+ $Y2=0
cc_856 N_A_840_107#_M40_noxref_g N_VPWR_c_2008_n 0.023923f $X=5.23 $Y=3.175
+ $X2=0 $Y2=0
cc_857 N_A_840_107#_M1043_d N_VPWR_c_1981_n 7.12537e-19 $X=7.83 $Y=2.855 $X2=0
+ $Y2=0
cc_858 N_A_840_107#_M39_noxref_g N_VPWR_c_1981_n 0.015425f $X=4.45 $Y=3.175
+ $X2=0 $Y2=0
cc_859 N_A_840_107#_M40_noxref_g N_VPWR_c_1981_n 0.00929096f $X=5.23 $Y=3.175
+ $X2=0 $Y2=0
cc_860 N_A_840_107#_c_988_n N_VPWR_c_1981_n 0.0133732f $X=6.015 $Y=4.905 $X2=0
+ $Y2=0
cc_861 N_A_840_107#_M1022_g N_VPWR_c_1981_n 0.0147436f $X=6.8 $Y=3.605 $X2=0
+ $Y2=0
cc_862 N_A_840_107#_c_997_n N_VPWR_c_1981_n 0.0350487f $X=7.97 $Y=3 $X2=0 $Y2=0
cc_863 N_A_840_107#_M1043_d N_VPWR_c_1982_n 3.64366e-19 $X=7.83 $Y=2.855 $X2=0
+ $Y2=0
cc_864 N_A_840_107#_M39_noxref_g N_VPWR_c_1982_n 0.00247029f $X=4.45 $Y=3.175
+ $X2=0 $Y2=0
cc_865 N_A_840_107#_M40_noxref_g N_VPWR_c_1982_n 0.00247029f $X=5.23 $Y=3.175
+ $X2=0 $Y2=0
cc_866 N_A_840_107#_c_988_n N_VPWR_c_1982_n 0.0224473f $X=6.015 $Y=4.905 $X2=0
+ $Y2=0
cc_867 N_A_840_107#_c_990_n N_VPWR_c_1982_n 0.00260696f $X=6.55 $Y=5.07 $X2=0
+ $Y2=0
cc_868 N_A_840_107#_M1022_g N_VPWR_c_1982_n 0.039181f $X=6.8 $Y=3.605 $X2=0
+ $Y2=0
cc_869 N_A_840_107#_c_997_n N_VPWR_c_1982_n 0.0438953f $X=7.97 $Y=3 $X2=0 $Y2=0
cc_870 N_A_840_107#_c_1001_n N_VPWR_c_1982_n 0.0243238f $X=7.87 $Y=5.07 $X2=0
+ $Y2=0
cc_871 N_A_840_107#_c_1002_n N_VPWR_c_1982_n 0.0171453f $X=7.87 $Y=5.07 $X2=0
+ $Y2=0
cc_872 N_A_840_107#_M1022_g N_A_1410_571#_c_2253_n 0.00388367f $X=6.8 $Y=3.605
+ $X2=0 $Y2=8.025
cc_873 N_A_840_107#_c_997_n N_A_1410_571#_c_2253_n 0.00837899f $X=7.97 $Y=3
+ $X2=0 $Y2=8.025
cc_874 N_A_840_107#_c_1002_n N_A_1410_571#_c_2253_n 0.00469412f $X=7.87 $Y=5.07
+ $X2=0 $Y2=8.025
cc_875 N_A_840_107#_M1022_g N_A_1410_571#_c_2254_n 0.00257634f $X=6.8 $Y=3.605
+ $X2=0 $Y2=0
cc_876 N_A_840_107#_M1022_g N_A_1410_571#_c_2262_n 4.56686e-19 $X=6.8 $Y=3.605
+ $X2=0 $Y2=0
cc_877 N_A_840_107#_c_997_n N_A_1410_571#_c_2262_n 0.00448047f $X=7.97 $Y=3
+ $X2=0 $Y2=0
cc_878 N_A_362_1243#_c_1126_n N_A_528_1171#_M1004_g 0.00441776f $X=3.68 $Y=6.36
+ $X2=0 $Y2=0
cc_879 N_A_362_1243#_c_1124_n N_A_528_1171#_c_1613_n 0.00204387f $X=3.57
+ $Y=5.865 $X2=0.24 $Y2=0
cc_880 N_A_362_1243#_c_1126_n N_A_528_1171#_c_1613_n 0.0112496f $X=3.68 $Y=6.36
+ $X2=0.24 $Y2=0
cc_881 N_A_362_1243#_c_1127_n N_A_528_1171#_c_1613_n 0.00204387f $X=5.93
+ $Y=5.865 $X2=0.24 $Y2=0
cc_882 N_A_362_1243#_c_1139_n N_A_528_1171#_c_1613_n 0.00605942f $X=3.68
+ $Y=5.865 $X2=0.24 $Y2=0
cc_883 N_A_362_1243#_c_1123_n N_A_528_1171#_c_1614_n 0.00670407f $X=1.95 $Y=6.36
+ $X2=0 $Y2=0
cc_884 N_A_362_1243#_c_1124_n N_A_528_1171#_c_1614_n 0.063842f $X=3.57 $Y=5.865
+ $X2=0 $Y2=0
cc_885 N_A_362_1243#_c_1126_n N_A_528_1171#_M1010_g 0.00441776f $X=3.68 $Y=6.36
+ $X2=0 $Y2=0
cc_886 N_A_362_1243#_c_1127_n N_A_528_1171#_c_1616_n 0.0130802f $X=5.93 $Y=5.865
+ $X2=24.72 $Y2=0
cc_887 N_A_362_1243#_c_1128_n N_A_528_1171#_M1023_g 0.00441776f $X=6.04 $Y=6.36
+ $X2=0 $Y2=0
cc_888 N_A_362_1243#_c_1127_n N_A_528_1171#_c_1618_n 0.00198257f $X=5.93
+ $Y=5.865 $X2=0.24 $Y2=8.14
cc_889 N_A_362_1243#_c_1128_n N_A_528_1171#_c_1618_n 0.0120486f $X=6.04 $Y=6.36
+ $X2=0.24 $Y2=8.14
cc_890 N_A_362_1243#_c_1130_n N_A_528_1171#_c_1618_n 0.00779303f $X=6.41
+ $Y=5.865 $X2=0.24 $Y2=8.14
cc_891 N_A_362_1243#_c_1128_n N_A_528_1171#_M1040_g 0.00441776f $X=6.04 $Y=6.36
+ $X2=0 $Y2=0
cc_892 N_A_362_1243#_c_1130_n N_A_528_1171#_c_1620_n 0.0034036f $X=6.41 $Y=5.865
+ $X2=0 $Y2=0
cc_893 N_A_362_1243#_c_1129_n N_A_528_1171#_c_1647_n 0.0102184f $X=6.41 $Y=3
+ $X2=0 $Y2=0
cc_894 N_A_362_1243#_c_1134_n N_A_528_1171#_c_1621_n 0.0481957f $X=7.33 $Y=2.35
+ $X2=0 $Y2=0
cc_895 N_A_362_1243#_c_1127_n N_A_528_1171#_c_1631_n 0.0656957f $X=5.93 $Y=5.865
+ $X2=0 $Y2=0
cc_896 N_A_362_1243#_c_1127_n N_A_528_1171#_c_1632_n 0.0656957f $X=5.93 $Y=5.865
+ $X2=0 $Y2=0
cc_897 N_A_362_1243#_c_1129_n N_A_528_1171#_c_1633_n 5.75622e-19 $X=6.41 $Y=3
+ $X2=0 $Y2=0
cc_898 N_A_362_1243#_c_1130_n N_A_528_1171#_c_1633_n 0.0291801f $X=6.41 $Y=5.865
+ $X2=0 $Y2=0
cc_899 N_A_362_1243#_c_1124_n N_X_c_1927_n 0.00613736f $X=3.57 $Y=5.865 $X2=0.24
+ $Y2=8.14
cc_900 N_A_362_1243#_c_1125_n N_VPWR_c_2117_n 0.00668482f $X=2.06 $Y=5.865 $X2=0
+ $Y2=0
cc_901 N_A_362_1243#_c_1124_n N_VPWR_c_2118_n 0.00494461f $X=3.57 $Y=5.865 $X2=0
+ $Y2=0
cc_902 N_A_362_1243#_c_1139_n N_VPWR_c_2118_n 0.00184991f $X=3.68 $Y=5.865 $X2=0
+ $Y2=0
cc_903 N_A_362_1243#_M1022_s N_VPWR_c_1981_n 7.12537e-19 $X=6.285 $Y=2.855 $X2=0
+ $Y2=0
cc_904 N_A_362_1243#_M1043_g N_VPWR_c_1981_n 0.0144787f $X=7.58 $Y=3.605 $X2=0
+ $Y2=0
cc_905 N_A_362_1243#_c_1129_n N_VPWR_c_1981_n 0.0325607f $X=6.41 $Y=3 $X2=0
+ $Y2=0
cc_906 N_A_362_1243#_M1022_s N_VPWR_c_1982_n 3.64366e-19 $X=6.285 $Y=2.855 $X2=0
+ $Y2=0
cc_907 N_A_362_1243#_M1043_g N_VPWR_c_1982_n 0.0116149f $X=7.58 $Y=3.605 $X2=0
+ $Y2=0
cc_908 N_A_362_1243#_c_1129_n N_VPWR_c_1982_n 0.0449203f $X=6.41 $Y=3 $X2=0
+ $Y2=0
cc_909 N_A_362_1243#_M1043_g N_A_1410_571#_c_2253_n 0.00388367f $X=7.58 $Y=3.605
+ $X2=0 $Y2=8.025
cc_910 N_A_362_1243#_c_1129_n N_A_1410_571#_c_2253_n 0.00837899f $X=6.41 $Y=3
+ $X2=0 $Y2=8.025
cc_911 N_A_362_1243#_M1043_g N_A_1410_571#_c_2254_n 0.0122342f $X=7.58 $Y=3.605
+ $X2=0 $Y2=0
cc_912 N_A_362_1243#_c_1134_n N_A_1410_571#_c_2254_n 6.73161e-19 $X=7.33 $Y=2.35
+ $X2=0 $Y2=0
cc_913 N_A_362_1243#_c_1134_n N_A_1410_571#_c_2245_n 0.0214273f $X=7.33 $Y=2.35
+ $X2=0.24 $Y2=0
cc_914 N_A_362_1243#_c_1144_n N_A_1410_571#_c_2245_n 0.00674932f $X=6.83 $Y=2.35
+ $X2=0.24 $Y2=0
cc_915 N_A_362_1243#_c_1134_n N_A_1410_571#_c_2246_n 8.36977e-19 $X=7.33 $Y=2.35
+ $X2=0 $Y2=0
cc_916 N_A_362_1243#_M1043_g N_A_1410_571#_c_2262_n 0.00983498f $X=7.58 $Y=3.605
+ $X2=0 $Y2=0
cc_917 N_A_362_1243#_c_1134_n N_A_1410_571#_c_2262_n 0.00430668f $X=7.33 $Y=2.35
+ $X2=0 $Y2=0
cc_918 N_A_362_1243#_c_1129_n N_A_1410_571#_c_2262_n 0.00106964f $X=6.41 $Y=3
+ $X2=0 $Y2=0
cc_919 N_A_362_1243#_M1043_g N_A_1410_571#_c_2263_n 0.0186168f $X=7.58 $Y=3.605
+ $X2=10.215 $Y2=0
cc_920 N_A_362_1243#_c_1134_n N_A_1410_571#_c_2263_n 0.0259253f $X=7.33 $Y=2.35
+ $X2=10.215 $Y2=0
cc_921 N_A_362_1243#_c_1144_n N_A_1410_571#_c_2263_n 0.00623026f $X=6.83 $Y=2.35
+ $X2=10.215 $Y2=0
cc_922 N_A_2092_381#_M43_noxref_g N_A_1472_1171#_c_1316_n 0.0134488f $X=10.71
+ $Y=3.535 $X2=0 $Y2=0
cc_923 N_A_2092_381#_M44_noxref_g N_A_1472_1171#_c_1316_n 0.0134488f $X=11.49
+ $Y=3.535 $X2=0 $Y2=0
cc_924 N_A_2092_381#_M45_noxref_g N_A_1472_1171#_c_1316_n 0.0134488f $X=12.27
+ $Y=3.535 $X2=0 $Y2=0
cc_925 N_A_2092_381#_M46_noxref_g N_A_1472_1171#_c_1316_n 0.0228224f $X=13.05
+ $Y=3.535 $X2=0 $Y2=0
cc_926 N_A_2092_381#_c_1230_n N_A_1472_1171#_c_1320_n 0.0438407f $X=11.49
+ $Y=5.535 $X2=0 $Y2=0
cc_927 N_A_2092_381#_c_1221_n N_A_1472_1171#_c_1323_n 0.0438407f $X=10.96
+ $Y=5.535 $X2=0 $Y2=0
cc_928 N_A_2092_381#_M46_noxref_g N_A_1472_1171#_c_1335_n 7.21002e-19 $X=13.05
+ $Y=3.535 $X2=24.72 $Y2=0
cc_929 N_A_2092_381#_M46_noxref_g N_A_1472_1171#_c_1324_n 0.00411764f $X=13.05
+ $Y=3.535 $X2=0 $Y2=0
cc_930 N_A_2092_381#_c_1216_n N_SLEEP_B_M1020_g 0.00973513f $X=13.595 $Y=5.59
+ $X2=0 $Y2=0
cc_931 N_A_2092_381#_c_1235_n N_SLEEP_B_M1020_g 0.021518f $X=13.995 $Y=4.43
+ $X2=0 $Y2=0
cc_932 N_A_2092_381#_c_1237_n N_SLEEP_B_M1020_g 0.00704799f $X=13.995 $Y=5.59
+ $X2=0 $Y2=0
cc_933 N_A_2092_381#_c_1217_n N_SLEEP_B_c_1468_n 0.0196534f $X=13.995 $Y=6.36
+ $X2=0 $Y2=0
cc_934 N_A_2092_381#_c_1217_n N_SLEEP_B_c_1470_n 0.00821272f $X=13.995 $Y=6.36
+ $X2=0 $Y2=0
cc_935 N_A_2092_381#_c_1237_n N_SLEEP_B_c_1470_n 0.0158593f $X=13.995 $Y=5.59
+ $X2=0 $Y2=0
cc_936 N_A_2092_381#_M43_noxref_g N_VPWR_c_1994_n 0.00196405f $X=10.71 $Y=3.535
+ $X2=24.72 $Y2=0
cc_937 N_A_2092_381#_M43_noxref_g N_VPWR_c_1995_n 0.00967639f $X=10.71 $Y=3.535
+ $X2=10.215 $Y2=8.14
cc_938 N_A_2092_381#_M43_noxref_g N_VPWR_c_1997_n 0.0367379f $X=10.71 $Y=3.535
+ $X2=0 $Y2=0
cc_939 N_A_2092_381#_c_1220_n N_VPWR_c_1997_n 0.00244421f $X=11.24 $Y=5.535
+ $X2=0 $Y2=0
cc_940 N_A_2092_381#_M44_noxref_g N_VPWR_c_1997_n 0.0351373f $X=11.49 $Y=3.535
+ $X2=0 $Y2=0
cc_941 N_A_2092_381#_M44_noxref_g N_VPWR_c_1999_n 0.00156247f $X=11.49 $Y=3.535
+ $X2=0 $Y2=0
cc_942 N_A_2092_381#_M45_noxref_g N_VPWR_c_1999_n 0.00156247f $X=12.27 $Y=3.535
+ $X2=0 $Y2=0
cc_943 N_A_2092_381#_M44_noxref_g N_VPWR_c_2000_n 0.00405433f $X=11.49 $Y=3.535
+ $X2=0 $Y2=0
cc_944 N_A_2092_381#_M45_noxref_g N_VPWR_c_2000_n 0.00405433f $X=12.27 $Y=3.535
+ $X2=0 $Y2=0
cc_945 N_A_2092_381#_M45_noxref_g N_VPWR_c_2001_n 0.0358388f $X=12.27 $Y=3.535
+ $X2=0 $Y2=0
cc_946 N_A_2092_381#_c_1227_n N_VPWR_c_2001_n 0.00244324f $X=12.8 $Y=5.535 $X2=0
+ $Y2=0
cc_947 N_A_2092_381#_M46_noxref_g N_VPWR_c_2001_n 0.0428339f $X=13.05 $Y=3.535
+ $X2=0 $Y2=0
cc_948 N_A_2092_381#_c_1232_n N_VPWR_c_2001_n 6.73791e-19 $X=12.8 $Y=5.425 $X2=0
+ $Y2=0
cc_949 N_A_2092_381#_c_1233_n N_VPWR_c_2001_n 0.0360609f $X=13.885 $Y=5.59 $X2=0
+ $Y2=0
cc_950 N_A_2092_381#_c_1216_n N_VPWR_c_2001_n 0.00512504f $X=13.595 $Y=5.59
+ $X2=0 $Y2=0
cc_951 N_A_2092_381#_c_1235_n N_VPWR_c_2001_n 0.0118028f $X=13.995 $Y=4.43 $X2=0
+ $Y2=0
cc_952 N_A_2092_381#_M46_noxref_g N_VPWR_c_2002_n 0.00168129f $X=13.05 $Y=3.535
+ $X2=0 $Y2=0
cc_953 N_A_2092_381#_M46_noxref_g N_VPWR_c_2003_n 0.00967639f $X=13.05 $Y=3.535
+ $X2=0 $Y2=0
cc_954 N_A_2092_381#_c_1235_n N_VPWR_c_2003_n 0.0308129f $X=13.995 $Y=4.43 $X2=0
+ $Y2=0
cc_955 N_A_2092_381#_c_1235_n N_VPWR_c_2004_n 0.00134675f $X=13.995 $Y=4.43
+ $X2=0 $Y2=0
cc_956 N_A_2092_381#_c_1235_n N_VPWR_c_2006_n 0.00133858f $X=13.995 $Y=4.43
+ $X2=0 $Y2=0
cc_957 N_A_2092_381#_c_1224_n N_VPWR_c_2007_n 0.00263446f $X=12.02 $Y=5.535
+ $X2=0 $Y2=0
cc_958 N_A_2092_381#_c_1235_n N_VPWR_c_2009_n 0.0102944f $X=13.995 $Y=4.43 $X2=0
+ $Y2=0
cc_959 N_A_2092_381#_M43_noxref_g N_VPWR_c_2013_n 0.0138184f $X=10.71 $Y=3.535
+ $X2=0 $Y2=0
cc_960 N_A_2092_381#_M44_noxref_g N_VPWR_c_2015_n 0.0138184f $X=11.49 $Y=3.535
+ $X2=0 $Y2=0
cc_961 N_A_2092_381#_M45_noxref_g N_VPWR_c_2015_n 0.0138184f $X=12.27 $Y=3.535
+ $X2=0 $Y2=0
cc_962 N_A_2092_381#_M46_noxref_g N_VPWR_c_2016_n 0.0138184f $X=13.05 $Y=3.535
+ $X2=0 $Y2=0
cc_963 N_A_2092_381#_M43_noxref_g N_VPWR_c_1981_n 0.011743f $X=10.71 $Y=3.535
+ $X2=0 $Y2=0
cc_964 N_A_2092_381#_M44_noxref_g N_VPWR_c_1981_n 0.011743f $X=11.49 $Y=3.535
+ $X2=0 $Y2=0
cc_965 N_A_2092_381#_M45_noxref_g N_VPWR_c_1981_n 0.011743f $X=12.27 $Y=3.535
+ $X2=0 $Y2=0
cc_966 N_A_2092_381#_M46_noxref_g N_VPWR_c_1981_n 0.011743f $X=13.05 $Y=3.535
+ $X2=0 $Y2=0
cc_967 N_A_2092_381#_M1020_s N_VPWR_c_1982_n 0.00219125f $X=13.87 $Y=4.285 $X2=0
+ $Y2=0
cc_968 N_A_2092_381#_M43_noxref_g N_VPWR_c_1982_n 0.0161354f $X=10.71 $Y=3.535
+ $X2=0 $Y2=0
cc_969 N_A_2092_381#_M44_noxref_g N_VPWR_c_1982_n 0.0161354f $X=11.49 $Y=3.535
+ $X2=0 $Y2=0
cc_970 N_A_2092_381#_M45_noxref_g N_VPWR_c_1982_n 0.0161354f $X=12.27 $Y=3.535
+ $X2=0 $Y2=0
cc_971 N_A_2092_381#_M46_noxref_g N_VPWR_c_1982_n 0.0161354f $X=13.05 $Y=3.535
+ $X2=0 $Y2=0
cc_972 N_A_2092_381#_c_1235_n N_VPWR_c_1982_n 0.0349366f $X=13.995 $Y=4.43 $X2=0
+ $Y2=0
cc_973 N_A_2092_381#_M43_noxref_g N_A_1410_571#_c_2246_n 0.0134259f $X=10.71
+ $Y=3.535 $X2=0 $Y2=0
cc_974 N_A_2092_381#_M43_noxref_g N_A_1410_571#_c_2257_n 0.00759785f $X=10.71
+ $Y=3.535 $X2=24.72 $Y2=0
cc_975 N_A_2092_381#_M44_noxref_g N_A_1410_571#_c_2257_n 0.00759785f $X=11.49
+ $Y=3.535 $X2=24.72 $Y2=0
cc_976 N_A_2092_381#_M44_noxref_g N_A_1410_571#_c_2248_n 0.0134259f $X=11.49
+ $Y=3.535 $X2=0 $Y2=0
cc_977 N_A_2092_381#_M45_noxref_g N_A_1410_571#_c_2248_n 0.0134259f $X=12.27
+ $Y=3.535 $X2=0 $Y2=0
cc_978 N_A_2092_381#_M45_noxref_g N_A_1410_571#_c_2260_n 0.00759785f $X=12.27
+ $Y=3.535 $X2=0 $Y2=0
cc_979 N_A_2092_381#_M46_noxref_g N_A_1410_571#_c_2260_n 0.00759785f $X=13.05
+ $Y=3.535 $X2=0 $Y2=0
cc_980 N_A_1472_1171#_M1001_g N_A_528_1171#_M1040_g 0.0148916f $X=7.81 $Y=6.715
+ $X2=0 $Y2=0
cc_981 N_A_1472_1171#_c_1313_n N_A_528_1171#_c_1646_n 0.0752391f $X=8.26
+ $Y=5.955 $X2=0 $Y2=0
cc_982 N_A_1472_1171#_c_1315_n N_A_528_1171#_c_1646_n 0.103376f $X=8.865
+ $Y=5.855 $X2=0 $Y2=0
cc_983 N_A_1472_1171#_c_1317_n N_A_528_1171#_c_1621_n 0.103376f $X=8.965
+ $Y=1.435 $X2=0 $Y2=0
cc_984 N_A_1472_1171#_c_1317_n N_A_528_1171#_c_1622_n 0.370299f $X=8.965
+ $Y=1.435 $X2=10.215 $Y2=0
cc_985 N_A_1472_1171#_c_1325_n N_A_528_1171#_c_1622_n 0.10665f $X=18.28 $Y=1.455
+ $X2=10.215 $Y2=0
cc_986 N_A_1472_1171#_c_1326_n N_A_528_1171#_c_1622_n 0.00218009f $X=14.295
+ $Y=1.455 $X2=10.215 $Y2=0
cc_987 N_A_1472_1171#_c_1325_n N_A_528_1171#_c_1624_n 0.0243408f $X=18.28
+ $Y=1.455 $X2=24.72 $Y2=0
cc_988 N_A_1472_1171#_c_1325_n N_A_528_1171#_c_1625_n 0.00608982f $X=18.28
+ $Y=1.455 $X2=0 $Y2=0
cc_989 N_A_1472_1171#_c_1325_n N_A_528_1171#_M1007_g 0.0165335f $X=18.28
+ $Y=1.455 $X2=10.215 $Y2=8.14
cc_990 N_A_1472_1171#_c_1338_n N_A_528_1171#_c_1655_n 0.00203651f $X=18.43
+ $Y=2.505 $X2=24.72 $Y2=8.14
cc_991 N_A_1472_1171#_c_1339_n N_A_528_1171#_c_1655_n 0.00843595f $X=18.43
+ $Y=3.2 $X2=24.72 $Y2=8.14
cc_992 N_A_1472_1171#_c_1338_n N_A_528_1171#_c_1659_n 4.27055e-19 $X=18.43
+ $Y=2.505 $X2=0 $Y2=0
cc_993 N_A_1472_1171#_c_1339_n N_A_528_1171#_c_1659_n 0.0093403f $X=18.43 $Y=3.2
+ $X2=0 $Y2=0
cc_994 N_A_1472_1171#_c_1344_n N_A_528_1171#_c_1659_n 0.00908519f $X=19.165
+ $Y=2.42 $X2=0 $Y2=0
cc_995 N_A_1472_1171#_c_1347_n N_A_528_1171#_c_1659_n 7.59177e-19 $X=19.33
+ $Y=3.2 $X2=0 $Y2=0
cc_996 N_A_1472_1171#_c_1327_n N_A_528_1171#_M1009_g 0.0134748f $X=19.27 $Y=1.48
+ $X2=0 $Y2=0
cc_997 N_A_1472_1171#_c_1339_n N_A_528_1171#_c_1663_n 7.59177e-19 $X=18.43
+ $Y=3.2 $X2=0 $Y2=0
cc_998 N_A_1472_1171#_c_1344_n N_A_528_1171#_c_1663_n 0.00908519f $X=19.165
+ $Y=2.42 $X2=0 $Y2=0
cc_999 N_A_1472_1171#_c_1347_n N_A_528_1171#_c_1663_n 0.0093403f $X=19.33 $Y=3.2
+ $X2=0 $Y2=0
cc_1000 N_A_1472_1171#_c_1428_p N_A_528_1171#_c_1663_n 4.27055e-19 $X=19.33
+ $Y=2.5 $X2=0 $Y2=0
cc_1001 N_A_1472_1171#_c_1327_n N_A_528_1171#_M1014_g 0.0141141f $X=19.27
+ $Y=1.48 $X2=0 $Y2=0
cc_1002 N_A_1472_1171#_c_1347_n N_A_528_1171#_c_1667_n 0.0138014f $X=19.33
+ $Y=3.2 $X2=0 $Y2=0
cc_1003 N_A_1472_1171#_c_1353_n N_A_528_1171#_c_1667_n 0.0144581f $X=19.71
+ $Y=2.42 $X2=0 $Y2=0
cc_1004 N_A_1472_1171#_c_1329_n N_A_528_1171#_c_1667_n 0.00696961f $X=19.825
+ $Y=2.335 $X2=0 $Y2=0
cc_1005 N_A_1472_1171#_c_1428_p N_A_528_1171#_c_1667_n 9.50925e-19 $X=19.33
+ $Y=2.5 $X2=0 $Y2=0
cc_1006 N_A_1472_1171#_c_1328_n N_A_528_1171#_M1016_g 0.0190067f $X=19.71
+ $Y=1.48 $X2=0 $Y2=0
cc_1007 N_A_1472_1171#_c_1329_n N_A_528_1171#_M1016_g 0.0190395f $X=19.825
+ $Y=2.335 $X2=0 $Y2=0
cc_1008 N_A_1472_1171#_c_1313_n N_A_528_1171#_c_1633_n 0.0148916f $X=8.26
+ $Y=5.955 $X2=0 $Y2=0
cc_1009 N_A_1472_1171#_c_1325_n N_A_528_1171#_c_1635_n 0.0189135f $X=18.28
+ $Y=1.455 $X2=0 $Y2=0
cc_1010 N_A_1472_1171#_c_1325_n N_A_528_1171#_c_1636_n 0.0692391f $X=18.28
+ $Y=1.455 $X2=0 $Y2=0
cc_1011 N_A_1472_1171#_c_1338_n N_A_528_1171#_c_1636_n 0.0237598f $X=18.43
+ $Y=2.505 $X2=0 $Y2=0
cc_1012 N_A_1472_1171#_c_1327_n N_A_528_1171#_c_1636_n 0.0555696f $X=19.27
+ $Y=1.48 $X2=0 $Y2=0
cc_1013 N_A_1472_1171#_c_1344_n N_A_528_1171#_c_1636_n 0.0393875f $X=19.165
+ $Y=2.42 $X2=0 $Y2=0
cc_1014 N_A_1472_1171#_c_1328_n N_A_528_1171#_c_1636_n 0.00188044f $X=19.71
+ $Y=1.48 $X2=0 $Y2=0
cc_1015 N_A_1472_1171#_c_1329_n N_A_528_1171#_c_1636_n 0.0266022f $X=19.825
+ $Y=2.335 $X2=0 $Y2=0
cc_1016 N_A_1472_1171#_c_1330_n N_A_528_1171#_c_1636_n 0.021475f $X=18.405
+ $Y=1.455 $X2=0 $Y2=0
cc_1017 N_A_1472_1171#_c_1428_p N_A_528_1171#_c_1636_n 0.0219285f $X=19.33
+ $Y=2.5 $X2=0 $Y2=0
cc_1018 N_A_1472_1171#_c_1331_n N_A_528_1171#_c_1636_n 0.0146029f $X=19.355
+ $Y=1.48 $X2=0 $Y2=0
cc_1019 N_A_1472_1171#_c_1338_n N_A_528_1171#_c_1644_n 0.00144444f $X=18.43
+ $Y=2.505 $X2=0 $Y2=0
cc_1020 N_A_1472_1171#_c_1327_n N_A_528_1171#_c_1644_n 0.00336308f $X=19.27
+ $Y=1.48 $X2=0 $Y2=0
cc_1021 N_A_1472_1171#_c_1344_n N_A_528_1171#_c_1644_n 0.00131212f $X=19.165
+ $Y=2.42 $X2=0 $Y2=0
cc_1022 N_A_1472_1171#_c_1330_n N_A_528_1171#_c_1644_n 0.00326139f $X=18.405
+ $Y=1.455 $X2=0 $Y2=0
cc_1023 N_A_1472_1171#_c_1428_p N_A_528_1171#_c_1644_n 0.00144162f $X=19.33
+ $Y=2.5 $X2=0 $Y2=0
cc_1024 N_A_1472_1171#_c_1331_n N_A_528_1171#_c_1644_n 0.00232957f $X=19.355
+ $Y=1.48 $X2=0 $Y2=0
cc_1025 N_A_1472_1171#_c_1320_n N_VPWR_c_1997_n 0.00100185f $X=10.9 $Y=5.955
+ $X2=0 $Y2=0
cc_1026 N_A_1472_1171#_c_1323_n N_VPWR_c_1997_n 4.82835e-19 $X=10.17 $Y=5.955
+ $X2=0 $Y2=0
cc_1027 N_A_1472_1171#_c_1323_n N_VPWR_c_1998_n 0.00124225f $X=10.17 $Y=5.955
+ $X2=0 $Y2=0
cc_1028 N_A_1472_1171#_c_1316_n N_VPWR_c_2002_n 0.00665071f $X=13.965 $Y=1.435
+ $X2=0 $Y2=0
cc_1029 N_A_1472_1171#_c_1335_n N_VPWR_c_2002_n 0.010242f $X=14.13 $Y=1.78 $X2=0
+ $Y2=0
cc_1030 N_A_1472_1171#_c_1324_n N_VPWR_c_2002_n 0.00234257f $X=14.13 $Y=1.78
+ $X2=0 $Y2=0
cc_1031 N_A_1472_1171#_c_1315_n N_VPWR_c_1981_n 0.0153416f $X=8.865 $Y=5.855
+ $X2=0 $Y2=0
cc_1032 N_A_1472_1171#_c_1339_n N_VPWR_c_1981_n 0.002574f $X=18.43 $Y=3.2 $X2=0
+ $Y2=0
cc_1033 N_A_1472_1171#_c_1347_n N_VPWR_c_1981_n 0.002574f $X=19.33 $Y=3.2 $X2=0
+ $Y2=0
cc_1034 N_A_1472_1171#_c_1315_n N_VPWR_c_1982_n 0.022562f $X=8.865 $Y=5.855
+ $X2=0 $Y2=0
cc_1035 N_A_1472_1171#_c_1315_n N_A_1410_571#_c_2246_n 0.0236262f $X=8.865
+ $Y=5.855 $X2=0 $Y2=0
cc_1036 N_A_1472_1171#_c_1316_n N_A_1410_571#_c_2246_n 0.0729684f $X=13.965
+ $Y=1.435 $X2=0 $Y2=0
cc_1037 N_A_1472_1171#_c_1316_n N_A_1410_571#_c_2248_n 0.0514307f $X=13.965
+ $Y=1.435 $X2=0 $Y2=0
cc_1038 N_A_1472_1171#_c_1316_n N_A_1410_571#_c_2249_n 0.0105968f $X=13.965
+ $Y=1.435 $X2=12.48 $Y2=0
cc_1039 N_SLEEP_B_M1020_g N_VPWR_c_2003_n 0.00379137f $X=14.385 $Y=4.66 $X2=0
+ $Y2=0
cc_1040 N_SLEEP_B_M1020_g N_VPWR_c_2004_n 9.491e-19 $X=14.385 $Y=4.66 $X2=0
+ $Y2=0
cc_1041 N_SLEEP_B_M1020_g N_VPWR_c_2006_n 0.00277795f $X=14.385 $Y=4.66 $X2=0
+ $Y2=0
cc_1042 N_SLEEP_B_c_1469_n N_VPWR_c_2006_n 0.0043047f $X=14.82 $Y=5.71 $X2=0
+ $Y2=0
cc_1043 N_SLEEP_B_c_1470_n N_VPWR_c_2006_n 0.00871549f $X=14.82 $Y=5.71 $X2=0
+ $Y2=0
cc_1044 N_SLEEP_B_M1020_g N_VPWR_c_2009_n 0.0238988f $X=14.385 $Y=4.66 $X2=0
+ $Y2=0
cc_1045 N_SLEEP_B_M1020_g N_VPWR_c_1981_n 0.00227564f $X=14.385 $Y=4.66 $X2=0
+ $Y2=0
cc_1046 N_SLEEP_B_M1020_g N_VPWR_c_1982_n 0.026804f $X=14.385 $Y=4.66 $X2=0
+ $Y2=0
cc_1047 N_A_3617_1198#_c_1508_n N_A_528_1171#_c_1639_n 0.0050126f $X=18.175
+ $Y=5.99 $X2=0 $Y2=0
cc_1048 N_A_3617_1198#_c_1500_n N_A_528_1171#_c_1639_n 0.0266022f $X=19.725
+ $Y=6.19 $X2=0 $Y2=0
cc_1049 N_A_3617_1198#_c_1507_n N_A_528_1171#_c_1639_n 0.0190395f $X=19.525
+ $Y=6.197 $X2=0 $Y2=0
cc_1050 N_A_3617_1198#_c_1508_n N_A_528_1171#_c_1682_n 0.0180205f $X=18.175
+ $Y=5.99 $X2=0 $Y2=0
cc_1051 N_A_3617_1198#_M1018_g N_A_528_1171#_c_1640_n 0.0190067f $X=18.16
+ $Y=7.015 $X2=0 $Y2=0
cc_1052 N_A_3617_1198#_c_1500_n N_A_528_1171#_c_1640_n 0.00188044f $X=19.725
+ $Y=6.19 $X2=0 $Y2=0
cc_1053 N_A_3617_1198#_c_1508_n N_A_528_1171#_c_1684_n 0.014949f $X=18.175
+ $Y=5.99 $X2=0 $Y2=0
cc_1054 N_A_3617_1198#_c_1511_n N_A_528_1171#_c_1684_n 0.0103122f $X=18.625
+ $Y=5.99 $X2=0 $Y2=0
cc_1055 N_A_3617_1198#_c_1514_n N_A_528_1171#_c_1684_n 6.45594e-19 $X=19.075
+ $Y=5.99 $X2=0 $Y2=0
cc_1056 N_A_3617_1198#_M1019_g N_A_528_1171#_c_1642_n 0.0141141f $X=18.59
+ $Y=7.015 $X2=0 $Y2=0
cc_1057 N_A_3617_1198#_M1027_g N_A_528_1171#_c_1642_n 0.0133424f $X=19.07
+ $Y=7.015 $X2=0 $Y2=0
cc_1058 N_A_3617_1198#_M1033_g N_A_528_1171#_c_1642_n 0.00187357f $X=19.54
+ $Y=7.015 $X2=0 $Y2=0
cc_1059 N_A_3617_1198#_c_1500_n N_A_528_1171#_c_1642_n 0.0770446f $X=19.725
+ $Y=6.19 $X2=0 $Y2=0
cc_1060 N_A_3617_1198#_c_1507_n N_A_528_1171#_c_1642_n 0.00662447f $X=19.525
+ $Y=6.197 $X2=0 $Y2=0
cc_1061 N_A_3617_1198#_c_1511_n N_A_528_1171#_c_1688_n 0.0120074f $X=18.625
+ $Y=5.99 $X2=0 $Y2=0
cc_1062 N_A_3617_1198#_c_1514_n N_A_528_1171#_c_1688_n 0.0120074f $X=19.075
+ $Y=5.99 $X2=0 $Y2=0
cc_1063 N_A_3617_1198#_c_1500_n N_A_528_1171#_c_1688_n 0.0393875f $X=19.725
+ $Y=6.19 $X2=0 $Y2=0
cc_1064 N_A_3617_1198#_c_1507_n N_A_528_1171#_c_1688_n 0.00131212f $X=19.525
+ $Y=6.197 $X2=0 $Y2=0
cc_1065 N_A_3617_1198#_c_1514_n N_A_528_1171#_c_1690_n 4.27055e-19 $X=19.075
+ $Y=5.99 $X2=0 $Y2=0
cc_1066 N_A_3617_1198#_c_1517_n N_A_528_1171#_c_1690_n 0.00203208f $X=19.525
+ $Y=5.99 $X2=0 $Y2=0
cc_1067 N_A_3617_1198#_c_1500_n N_A_528_1171#_c_1690_n 0.0237598f $X=19.725
+ $Y=6.19 $X2=0 $Y2=0
cc_1068 N_A_3617_1198#_c_1507_n N_A_528_1171#_c_1690_n 0.00144444f $X=19.525
+ $Y=6.197 $X2=0 $Y2=0
cc_1069 N_A_3617_1198#_c_1511_n N_A_528_1171#_c_1691_n 6.45594e-19 $X=18.625
+ $Y=5.99 $X2=0 $Y2=0
cc_1070 N_A_3617_1198#_c_1514_n N_A_528_1171#_c_1691_n 0.0103122f $X=19.075
+ $Y=5.99 $X2=0 $Y2=0
cc_1071 N_A_3617_1198#_c_1517_n N_A_528_1171#_c_1691_n 0.00957191f $X=19.525
+ $Y=5.99 $X2=0 $Y2=0
cc_1072 N_A_3617_1198#_c_1508_n N_A_528_1171#_c_1696_n 0.00226699f $X=18.175
+ $Y=5.99 $X2=0 $Y2=0
cc_1073 N_A_3617_1198#_c_1508_n N_A_528_1171#_c_1847_n 9.50925e-19 $X=18.175
+ $Y=5.99 $X2=0 $Y2=0
cc_1074 N_A_3617_1198#_c_1511_n N_A_528_1171#_c_1847_n 4.27055e-19 $X=18.625
+ $Y=5.99 $X2=0 $Y2=0
cc_1075 N_A_3617_1198#_c_1500_n N_A_528_1171#_c_1847_n 0.0219285f $X=19.725
+ $Y=6.19 $X2=0 $Y2=0
cc_1076 N_A_3617_1198#_c_1507_n N_A_528_1171#_c_1847_n 0.00144162f $X=19.525
+ $Y=6.197 $X2=0 $Y2=0
cc_1077 N_A_3617_1198#_c_1500_n N_A_528_1171#_c_1643_n 0.0146029f $X=19.725
+ $Y=6.19 $X2=0 $Y2=0
cc_1078 N_A_3617_1198#_c_1507_n N_A_528_1171#_c_1643_n 0.00232957f $X=19.525
+ $Y=6.197 $X2=0 $Y2=0
cc_1079 N_A_3617_1198#_c_1502_n N_A_c_1874_n 0.0033656f $X=20.785 $Y=4.94 $X2=0
+ $Y2=0
cc_1080 N_A_3617_1198#_c_1504_n N_A_c_1874_n 0.00340125f $X=19.94 $Y=6.19 $X2=0
+ $Y2=0
cc_1081 N_A_3617_1198#_c_1501_n N_A_c_1867_n 0.010937f $X=20.615 $Y=6.295 $X2=0
+ $Y2=0
cc_1082 N_A_3617_1198#_c_1502_n N_A_c_1867_n 0.00342021f $X=20.785 $Y=4.94 $X2=0
+ $Y2=0
cc_1083 N_A_3617_1198#_c_1505_n N_A_c_1867_n 0.00149998f $X=20.757 $Y=6.295
+ $X2=0 $Y2=0
cc_1084 N_A_3617_1198#_c_1502_n N_A_c_1876_n 0.016332f $X=20.785 $Y=4.94 $X2=0
+ $Y2=0
cc_1085 N_A_3617_1198#_c_1504_n N_A_c_1876_n 2.22502e-19 $X=19.94 $Y=6.19 $X2=0
+ $Y2=0
cc_1086 N_A_3617_1198#_c_1503_n N_A_M1024_g 0.00828462f $X=20.78 $Y=6.79 $X2=0
+ $Y2=0
cc_1087 N_A_3617_1198#_c_1506_n N_A_M1024_g 0.00881083f $X=20.78 $Y=6.625 $X2=0
+ $Y2=0
cc_1088 N_A_3617_1198#_c_1505_n N_A_c_1869_n 0.0059624f $X=20.757 $Y=6.295 $X2=0
+ $Y2=0
cc_1089 N_A_3617_1198#_c_1506_n N_A_c_1869_n 0.00424976f $X=20.78 $Y=6.625 $X2=0
+ $Y2=0
cc_1090 N_A_3617_1198#_c_1502_n N_A_c_1870_n 0.0016147f $X=20.785 $Y=4.94 $X2=0
+ $Y2=8.025
cc_1091 N_A_3617_1198#_c_1505_n N_A_c_1870_n 0.00118692f $X=20.757 $Y=6.295
+ $X2=0 $Y2=8.025
cc_1092 N_A_3617_1198#_c_1503_n N_A_M1046_g 0.00950623f $X=20.78 $Y=6.79 $X2=0
+ $Y2=0
cc_1093 N_A_3617_1198#_c_1506_n N_A_M1046_g 0.00465421f $X=20.78 $Y=6.625 $X2=0
+ $Y2=0
cc_1094 N_A_3617_1198#_c_1502_n N_A_c_1883_n 0.0021175f $X=20.785 $Y=4.94
+ $X2=0.24 $Y2=0
cc_1095 N_A_3617_1198#_c_1501_n N_A_c_1872_n 0.0102472f $X=20.615 $Y=6.295 $X2=0
+ $Y2=0
cc_1096 N_A_3617_1198#_c_1505_n N_A_c_1872_n 3.29575e-19 $X=20.757 $Y=6.295
+ $X2=0 $Y2=0
cc_1097 N_A_3617_1198#_c_1506_n N_A_c_1872_n 0.00215258f $X=20.78 $Y=6.625 $X2=0
+ $Y2=0
cc_1098 N_A_3617_1198#_c_1502_n A 0.0163467f $X=20.785 $Y=4.94 $X2=0 $Y2=0
cc_1099 N_A_3617_1198#_c_1505_n A 0.0181008f $X=20.757 $Y=6.295 $X2=0 $Y2=0
cc_1100 N_A_3617_1198#_c_1506_n A 0.00367389f $X=20.78 $Y=6.625 $X2=0 $Y2=0
cc_1101 N_A_3617_1198#_c_1508_n N_VPWR_c_1982_n 0.00884289f $X=18.175 $Y=5.99
+ $X2=0 $Y2=0
cc_1102 N_A_3617_1198#_c_1511_n N_VPWR_c_1982_n 0.00855479f $X=18.625 $Y=5.99
+ $X2=0 $Y2=0
cc_1103 N_A_3617_1198#_c_1514_n N_VPWR_c_1982_n 0.00855479f $X=19.075 $Y=5.99
+ $X2=0 $Y2=0
cc_1104 N_A_3617_1198#_c_1517_n N_VPWR_c_1982_n 0.00884289f $X=19.525 $Y=5.99
+ $X2=0 $Y2=0
cc_1105 N_A_3617_1198#_c_1502_n N_VPWR_c_1982_n 0.00957445f $X=20.785 $Y=4.94
+ $X2=0 $Y2=0
cc_1106 N_A_528_1171#_c_1621_n N_VPWR_c_1981_n 0.012621f $X=8.365 $Y=5.445 $X2=0
+ $Y2=0
cc_1107 N_A_528_1171#_c_1655_n N_VPWR_c_1981_n 0.00387811f $X=18.205 $Y=2.15
+ $X2=0 $Y2=0
cc_1108 N_A_528_1171#_c_1659_n N_VPWR_c_1981_n 0.00359001f $X=18.655 $Y=2.15
+ $X2=0 $Y2=0
cc_1109 N_A_528_1171#_c_1663_n N_VPWR_c_1981_n 0.00359001f $X=19.105 $Y=2.15
+ $X2=0 $Y2=0
cc_1110 N_A_528_1171#_c_1667_n N_VPWR_c_1981_n 0.00387811f $X=19.555 $Y=2.15
+ $X2=0 $Y2=0
cc_1111 N_A_528_1171#_c_1634_n N_VPWR_c_1981_n 0.036594f $X=17.27 $Y=5.635 $X2=0
+ $Y2=0
cc_1112 N_A_528_1171#_c_1621_n N_VPWR_c_1982_n 0.0213855f $X=8.365 $Y=5.445
+ $X2=0 $Y2=0
cc_1113 N_A_528_1171#_c_1634_n N_VPWR_c_1982_n 0.046032f $X=17.27 $Y=5.635 $X2=0
+ $Y2=0
cc_1114 N_A_528_1171#_c_1684_n N_VPWR_c_1982_n 0.0110699f $X=18.4 $Y=4.94 $X2=0
+ $Y2=0
cc_1115 N_A_528_1171#_c_1691_n N_VPWR_c_1982_n 0.0110699f $X=19.3 $Y=4.94 $X2=0
+ $Y2=0
cc_1116 N_A_528_1171#_c_1621_n N_A_1410_571#_c_2245_n 0.0115846f $X=8.365
+ $Y=5.445 $X2=0.24 $Y2=0
cc_1117 N_A_528_1171#_c_1621_n N_A_1410_571#_c_2246_n 0.0299202f $X=8.365
+ $Y=5.445 $X2=0 $Y2=0
cc_1118 N_A_528_1171#_c_1622_n N_A_1410_571#_c_2246_n 0.0109634f $X=17.465
+ $Y=1.022 $X2=0 $Y2=0
cc_1119 N_A_528_1171#_c_1621_n N_A_1410_571#_c_2263_n 0.00125896f $X=8.365
+ $Y=5.445 $X2=10.215 $Y2=0
cc_1120 N_A_c_1876_n N_VPWR_c_1982_n 0.00866342f $X=20.56 $Y=5.99 $X2=0 $Y2=0
cc_1121 N_A_c_1883_n N_VPWR_c_1982_n 0.00804022f $X=21.01 $Y=5.99 $X2=0 $Y2=0
cc_1122 N_X_c_1921_n N_VPWR_c_1988_n 0.0143699f $X=2.62 $Y=2.03 $X2=0 $Y2=0
cc_1123 N_X_c_1927_n N_VPWR_c_1988_n 0.00995267f $X=2.73 $Y=2.57 $X2=0 $Y2=0
cc_1124 X N_VPWR_c_1988_n 0.00995267f $X=1.085 $Y=1.98 $X2=0 $Y2=0
cc_1125 N_X_c_1927_n N_VPWR_c_1990_n 0.00995267f $X=2.73 $Y=2.57 $X2=0 $Y2=0
cc_1126 N_X_c_1927_n N_VPWR_c_2117_n 6.82011e-19 $X=2.73 $Y=2.57 $X2=0 $Y2=0
cc_1127 X N_VPWR_c_2117_n 6.82011e-19 $X=1.085 $Y=1.98 $X2=0 $Y2=0
cc_1128 N_X_c_1927_n N_VPWR_c_2010_n 0.00470914f $X=2.73 $Y=2.57 $X2=0 $Y2=0
cc_1129 X N_VPWR_c_2010_n 0.00470914f $X=1.085 $Y=1.98 $X2=0 $Y2=0
cc_1130 N_X_c_1927_n N_VPWR_c_2118_n 6.82011e-19 $X=2.73 $Y=2.57 $X2=0 $Y2=0
cc_1131 N_X_c_1927_n N_VPWR_c_2011_n 0.00470914f $X=2.73 $Y=2.57 $X2=0 $Y2=0
cc_1132 N_X_M1005_s N_VPWR_c_1981_n 7.12537e-19 $X=1.045 $Y=2.425 $X2=0 $Y2=0
cc_1133 N_X_M1011_s N_VPWR_c_1981_n 9.06866e-19 $X=2.59 $Y=2.425 $X2=0 $Y2=0
cc_1134 N_X_c_1927_n N_VPWR_c_1981_n 0.0322386f $X=2.73 $Y=2.57 $X2=0 $Y2=0
cc_1135 X N_VPWR_c_1981_n 0.0350487f $X=1.085 $Y=1.98 $X2=0 $Y2=0
cc_1136 N_X_M1005_s N_VPWR_c_1982_n 0.00219125f $X=1.045 $Y=2.425 $X2=0 $Y2=0
cc_1137 N_X_M1011_s N_VPWR_c_1982_n 0.00278887f $X=2.59 $Y=2.425 $X2=0 $Y2=0
cc_1138 N_X_c_1927_n N_VPWR_c_1982_n 0.0383084f $X=2.73 $Y=2.57 $X2=0 $Y2=0
cc_1139 X N_VPWR_c_1982_n 0.0390242f $X=1.085 $Y=1.98 $X2=0 $Y2=0
cc_1140 N_VPWR_c_1981_n N_A_1410_571#_M1022_d 6.7971e-19 $X=13.62 $Y=3.63 $X2=0
+ $Y2=0
cc_1141 N_VPWR_c_1982_n N_A_1410_571#_M1022_d 3.88657e-19 $X=14.77 $Y=4.51 $X2=0
+ $Y2=0
cc_1142 N_VPWR_c_1981_n N_A_1410_571#_M43_noxref_d 9.06866e-19 $X=13.62 $Y=3.63
+ $X2=0 $Y2=0
cc_1143 N_VPWR_c_1982_n N_A_1410_571#_M43_noxref_d 0.00104903f $X=14.77 $Y=4.51
+ $X2=0 $Y2=0
cc_1144 N_VPWR_c_1981_n N_A_1410_571#_M45_noxref_d 9.06866e-19 $X=13.62 $Y=3.63
+ $X2=0 $Y2=0
cc_1145 N_VPWR_c_1982_n N_A_1410_571#_M45_noxref_d 0.00104903f $X=14.77 $Y=4.51
+ $X2=0 $Y2=0
cc_1146 N_VPWR_c_1981_n N_A_1410_571#_c_2253_n 0.0327821f $X=13.62 $Y=3.63 $X2=0
+ $Y2=8.025
cc_1147 N_VPWR_c_1982_n N_A_1410_571#_c_2253_n 0.0112297f $X=14.77 $Y=4.51 $X2=0
+ $Y2=8.025
cc_1148 N_VPWR_c_1994_n N_A_1410_571#_c_2246_n 0.0161483f $X=10.32 $Y=2.18 $X2=0
+ $Y2=0
cc_1149 N_VPWR_c_1994_n N_A_1410_571#_c_2257_n 0.00405296f $X=10.32 $Y=2.18
+ $X2=24.72 $Y2=0
cc_1150 N_VPWR_c_1995_n N_A_1410_571#_c_2257_n 0.0064384f $X=10.32 $Y=3.88
+ $X2=24.72 $Y2=0
cc_1151 N_VPWR_c_1997_n N_A_1410_571#_c_2257_n 0.00866266f $X=11.77 $Y=5.145
+ $X2=24.72 $Y2=0
cc_1152 N_VPWR_c_1999_n N_A_1410_571#_c_2257_n 0.00405296f $X=11.88 $Y=2.18
+ $X2=24.72 $Y2=0
cc_1153 N_VPWR_c_2000_n N_A_1410_571#_c_2257_n 0.0064384f $X=11.88 $Y=3.88
+ $X2=24.72 $Y2=0
cc_1154 N_VPWR_c_2013_n N_A_1410_571#_c_2257_n 0.00470914f $X=10.5 $Y=3.63
+ $X2=24.72 $Y2=0
cc_1155 N_VPWR_c_2015_n N_A_1410_571#_c_2257_n 0.00470914f $X=12.06 $Y=3.63
+ $X2=24.72 $Y2=0
cc_1156 N_VPWR_c_1981_n N_A_1410_571#_c_2257_n 0.0298862f $X=13.62 $Y=3.63
+ $X2=24.72 $Y2=0
cc_1157 N_VPWR_c_1982_n N_A_1410_571#_c_2257_n 0.0324723f $X=14.77 $Y=4.51
+ $X2=24.72 $Y2=0
cc_1158 N_VPWR_c_1999_n N_A_1410_571#_c_2248_n 0.0161483f $X=11.88 $Y=2.18 $X2=0
+ $Y2=0
cc_1159 N_VPWR_c_1999_n N_A_1410_571#_c_2260_n 0.00405296f $X=11.88 $Y=2.18
+ $X2=0 $Y2=0
cc_1160 N_VPWR_c_2000_n N_A_1410_571#_c_2260_n 0.0064384f $X=11.88 $Y=3.88 $X2=0
+ $Y2=0
cc_1161 N_VPWR_c_2001_n N_A_1410_571#_c_2260_n 0.00866266f $X=13.33 $Y=5.145
+ $X2=0 $Y2=0
cc_1162 N_VPWR_c_2002_n N_A_1410_571#_c_2260_n 0.00405296f $X=13.44 $Y=2.18
+ $X2=0 $Y2=0
cc_1163 N_VPWR_c_2003_n N_A_1410_571#_c_2260_n 0.0064384f $X=13.44 $Y=3.88 $X2=0
+ $Y2=0
cc_1164 N_VPWR_c_2015_n N_A_1410_571#_c_2260_n 0.00470914f $X=12.06 $Y=3.63
+ $X2=0 $Y2=0
cc_1165 N_VPWR_c_2016_n N_A_1410_571#_c_2260_n 0.00470914f $X=13.62 $Y=3.63
+ $X2=0 $Y2=0
cc_1166 N_VPWR_c_1981_n N_A_1410_571#_c_2260_n 0.0298862f $X=13.62 $Y=3.63 $X2=0
+ $Y2=0
cc_1167 N_VPWR_c_1982_n N_A_1410_571#_c_2260_n 0.0324723f $X=14.77 $Y=4.51 $X2=0
+ $Y2=0
cc_1168 N_VPWR_c_1981_n N_A_1410_571#_c_2262_n 0.00132323f $X=13.62 $Y=3.63
+ $X2=0 $Y2=0
