* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VNB VPB VPWR X
X0 a_30_207# a_30_1337# a_187_207# VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X1 a_30_443# a_30_1337# a_30_207# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X2 X a_389_141# a_187_207# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X5 X a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X6 a_389_141# a_389_1337# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X7 a_187_207# a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X8 a_389_141# a_30_207# a_187_207# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X9 a_389_141# a_30_207# a_187_207# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X10 VPWR A a_30_1337# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=500000u
X11 a_30_1337# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=420000u l=500000u
X12 LVPWR a_389_141# a_389_1337# LVPWR sky130_fd_pr__pfet_01v8_hvt w=1.12e+06u l=150000u
X13 a_389_141# a_30_207# a_187_207# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X14 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X15 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
.ends
