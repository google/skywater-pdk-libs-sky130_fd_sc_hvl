* File: sky130_fd_sc_hvl__sdfxbp_1.pex.spice
* Created: Fri Aug 28 09:40:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%VNB 5 7 11
c119 11 0 1.67566e-19 $X=0.24 $Y=0
r120 7 11 0.000362043 $w=1.968e-05 $l=5.7e-08 $layer=MET1_cond $X=9.84 $Y=0.057
+ $X2=9.84 $Y2=0
r121 5 11 0.453659 $w=1.7e-07 $l=3.485e-06 $layer=mcon $count=20 $X=19.44 $Y=0
+ $X2=19.44 $Y2=0
r122 5 11 0.453659 $w=1.7e-07 $l=3.485e-06 $layer=mcon $count=20 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%VPB 4 6 14
c177 6 0 1.50317e-20 $X=9.84 $Y=4.013
r178 10 14 0.453659 $w=1.7e-07 $l=3.485e-06 $layer=mcon $count=20 $X=19.44
+ $Y=4.07 $X2=19.44 $Y2=4.07
r179 9 14 1252.62 $w=1.68e-07 $l=1.92e-05 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=19.44 $Y2=4.07
r180 9 10 0.453659 $w=1.7e-07 $l=3.485e-06 $layer=mcon $count=20 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r181 6 10 0.000362043 $w=1.968e-05 $l=5.7e-08 $layer=MET1_cond $X=9.84 $Y=4.013
+ $X2=9.84 $Y2=4.07
r182 4 14 8.87805 $w=1.7e-07 $l=1.94825e-05 $layer=licon1_NTAP_notbjt $count=20
+ $X=0 $Y=3.985 $X2=19.44 $Y2=4.07
r183 4 9 8.87805 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=20
+ $X=0 $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%SCE 3 7 11 15 17 18 19 20 21 30 35 36 39
+ 49 50
c72 11 0 3.21733e-20 $X=2.585 $Y=0.745
c73 3 0 6.15916e-20 $X=0.665 $Y=2.785
r74 49 50 2.80859 $w=3.3e-07 $l=2.35e-07 $layer=LI1_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=1.75
r75 47 49 0.254485 $w=4.68e-07 $l=1e-08 $layer=LI1_cond $X=0.72 $Y=1.985
+ $X2=0.73 $Y2=1.985
r76 35 38 50.2236 $w=5.7e-07 $l=5.25e-07 $layer=POLY_cond $X=2.62 $Y=2.26
+ $X2=2.62 $Y2=2.785
r77 35 37 18.3095 $w=5.7e-07 $l=1.85e-07 $layer=POLY_cond $X=2.62 $Y=2.26
+ $X2=2.62 $Y2=2.075
r78 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.59
+ $Y=2.26 $X2=2.59 $Y2=2.26
r79 30 33 39.9482 $w=9.3e-07 $l=5.25e-07 $layer=POLY_cond $X=0.88 $Y=1.715
+ $X2=0.88 $Y2=2.24
r80 30 32 45.7534 $w=9.3e-07 $l=6.3e-07 $layer=POLY_cond $X=0.88 $Y=1.715
+ $X2=0.88 $Y2=1.085
r81 21 39 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=1.65 $X2=2.425
+ $Y2=1.65
r82 21 36 13.5837 $w=4.98e-07 $l=5.1e-07 $layer=LI1_cond $X=2.59 $Y=1.75
+ $X2=2.59 $Y2=2.26
r83 20 39 14.6955 $w=1.98e-07 $l=2.65e-07 $layer=LI1_cond $X=2.16 $Y=1.65
+ $X2=2.425 $Y2=1.65
r84 19 20 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.65
+ $X2=2.16 $Y2=1.65
r85 18 19 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.65 $X2=1.68
+ $Y2=1.65
r86 18 40 16.9136 $w=1.98e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=1.65
+ $X2=0.895 $Y2=1.65
r87 17 50 2.77883 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=0.73 $Y=1.65 $X2=0.73
+ $Y2=1.75
r88 17 40 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=1.65 $X2=0.895
+ $Y2=1.65
r89 17 47 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.72 $Y=1.75
+ $X2=0.72 $Y2=1.985
r90 17 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.73
+ $Y=1.715 $X2=0.73 $Y2=1.715
r91 15 38 77.0442 $w=5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.655 $Y=3.505
+ $X2=2.655 $Y2=2.785
r92 11 37 142.318 $w=5e-07 $l=1.33e-06 $layer=POLY_cond $X=2.585 $Y=0.745
+ $X2=2.585 $Y2=2.075
r93 7 32 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.095 $Y=0.745 $X2=1.095
+ $Y2=1.085
r94 3 33 58.3182 $w=5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.665 $Y=2.785
+ $X2=0.665 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%SCD 1 4 8 10
r28 7 10 159.439 $w=5e-07 $l=1.49e-06 $layer=POLY_cond $X=1.875 $Y=2.015
+ $X2=1.875 $Y2=3.505
r29 7 8 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.81 $Y=2.015
+ $X2=1.81 $Y2=2.015
r30 4 7 135.897 $w=5e-07 $l=1.27e-06 $layer=POLY_cond $X=1.875 $Y=0.745
+ $X2=1.875 $Y2=2.015
r31 1 8 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=1.77 $Y=2.035 $X2=1.77
+ $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_30_515# 1 2 9 12 15 19 23 24 27 29 34 35
+ 37 39 40
r86 40 43 50.2236 $w=5.7e-07 $l=5.25e-07 $layer=POLY_cond $X=3.33 $Y=1.34
+ $X2=3.33 $Y2=1.865
r87 40 42 24.8801 $w=5.7e-07 $l=2.55e-07 $layer=POLY_cond $X=3.33 $Y=1.34
+ $X2=3.33 $Y2=1.085
r88 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.23
+ $Y=1.34 $X2=3.23 $Y2=1.34
r89 34 35 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.275 $Y=2.785
+ $X2=0.275 $Y2=2.555
r90 30 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.87 $Y=1.26
+ $X2=0.705 $Y2=1.26
r91 29 39 4.40896 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.065 $Y=1.26
+ $X2=3.197 $Y2=1.26
r92 29 30 143.203 $w=1.68e-07 $l=2.195e-06 $layer=LI1_cond $X=3.065 $Y=1.26
+ $X2=0.87 $Y2=1.26
r93 25 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.175
+ $X2=0.705 $Y2=1.26
r94 25 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.705 $Y=1.175
+ $X2=0.705 $Y2=0.745
r95 23 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.54 $Y=1.26
+ $X2=0.705 $Y2=1.26
r96 23 24 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.54 $Y=1.26
+ $X2=0.28 $Y2=1.26
r97 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.195 $Y=1.345
+ $X2=0.28 $Y2=1.26
r98 21 35 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=0.195 $Y=1.345
+ $X2=0.195 $Y2=2.555
r99 17 19 66.3437 $w=5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.365 $Y=2.61
+ $X2=3.985 $Y2=2.61
r100 13 19 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.985 $Y=2.86
+ $X2=3.985 $Y2=2.61
r101 13 15 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.985 $Y=2.86
+ $X2=3.985 $Y2=3.2
r102 12 17 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.365 $Y=2.36
+ $X2=3.365 $Y2=2.61
r103 12 43 52.9679 $w=5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.365 $Y=2.36
+ $X2=3.365 $Y2=1.865
r104 9 42 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.365 $Y=0.745
+ $X2=3.365 $Y2=1.085
r105 2 34 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.575 $X2=0.275 $Y2=2.785
r106 1 27 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.535 $X2=0.705 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%D 3 7 9 10 11 20
c43 3 0 2.41303e-19 $X=4.075 $Y=0.745
r44 18 20 28.675 $w=7.8e-07 $l=4.35e-07 $layer=POLY_cond $X=4.33 $Y=1.475
+ $X2=4.765 $Y2=1.475
r45 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.33
+ $Y=1.34 $X2=4.33 $Y2=1.34
r46 15 18 16.8095 $w=7.8e-07 $l=2.55e-07 $layer=POLY_cond $X=4.075 $Y=1.475
+ $X2=4.33 $Y2=1.475
r47 10 11 8.67743 $w=5.08e-07 $l=3.7e-07 $layer=LI1_cond $X=4.42 $Y=1.665
+ $X2=4.42 $Y2=2.035
r48 10 19 7.62207 $w=5.08e-07 $l=3.25e-07 $layer=LI1_cond $X=4.42 $Y=1.665
+ $X2=4.42 $Y2=1.34
r49 9 19 1.05536 $w=5.08e-07 $l=4.5e-08 $layer=LI1_cond $X=4.42 $Y=1.295
+ $X2=4.42 $Y2=1.34
r50 5 20 13.1928 $w=5e-07 $l=3.9e-07 $layer=POLY_cond $X=4.765 $Y=1.865
+ $X2=4.765 $Y2=1.475
r51 5 7 142.853 $w=5e-07 $l=1.335e-06 $layer=POLY_cond $X=4.765 $Y=1.865
+ $X2=4.765 $Y2=3.2
r52 1 15 13.1928 $w=5e-07 $l=3.9e-07 $layer=POLY_cond $X=4.075 $Y=1.085
+ $X2=4.075 $Y2=1.475
r53 1 3 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.075 $Y=1.085 $X2=4.075
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1124_81# 1 2 7 9 10 12 13 19 20 22 24 27
+ 28 32
c92 22 0 1.87436e-19 $X=7.91 $Y=2.98
r93 32 34 11.4306 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=8.78 $Y=1.11
+ $X2=8.78 $Y2=1.36
r94 27 34 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=8.7 $Y=2.135
+ $X2=8.7 $Y2=1.36
r95 22 24 26.7367 $w=2.48e-07 $l=5.8e-07 $layer=LI1_cond $X=7.91 $Y=2.98
+ $X2=8.49 $Y2=2.98
r96 21 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=2.22
+ $X2=7.825 $Y2=2.22
r97 20 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.615 $Y=2.22
+ $X2=8.7 $Y2=2.135
r98 20 21 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=8.615 $Y=2.22
+ $X2=7.91 $Y2=2.22
r99 19 22 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.825 $Y=2.855
+ $X2=7.91 $Y2=2.98
r100 18 19 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.825 $Y=2.555
+ $X2=7.825 $Y2=2.855
r101 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.485
+ $Y=2.39 $X2=6.485 $Y2=2.39
r102 13 18 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.825 $Y=2.43
+ $X2=7.825 $Y2=2.555
r103 13 28 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.825 $Y=2.43
+ $X2=7.825 $Y2=2.22
r104 13 15 57.8526 $w=2.48e-07 $l=1.255e-06 $layer=LI1_cond $X=7.74 $Y=2.43
+ $X2=6.485 $Y2=2.43
r105 10 16 20.4123 $w=8.59e-07 $l=2.38694e-07 $layer=POLY_cond $X=6.095 $Y=2.605
+ $X2=6.145 $Y2=2.39
r106 10 12 58.804 $w=5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.095 $Y=2.605
+ $X2=6.095 $Y2=3.215
r107 7 16 64.1795 $w=8.59e-07 $l=1.12412e-06 $layer=POLY_cond $X=5.87 $Y=1.395
+ $X2=6.145 $Y2=2.39
r108 7 9 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=5.87 $Y=1.395 $X2=5.87
+ $Y2=0.91
r109 2 24 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=8.35
+ $Y=2.895 $X2=8.49 $Y2=3.02
r110 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.64
+ $Y=0.9 $X2=8.78 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1067_107# 1 2 3 4 13 15 18 22 26 30 31
+ 32 34 36 40 41 47 53 56 60
c163 53 0 4.11115e-20 $X=7.39 $Y=1.645
c164 13 0 8.01934e-20 $X=7.02 $Y=1.395
r165 60 63 24.3474 $w=3.53e-07 $l=7.5e-07 $layer=LI1_cond $X=13.617 $Y=2.35
+ $X2=13.617 $Y2=3.1
r166 52 53 39.5922 $w=5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.02 $Y=1.645
+ $X2=7.39 $Y2=1.645
r167 47 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.145
+ $X2=13.68 $Y2=3.145
r168 44 56 8.87693 $w=3.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.605 $Y=3.145
+ $X2=5.605 $Y2=2.86
r169 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.145
+ $X2=5.52 $Y2=3.145
r170 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=3.145
+ $X2=5.52 $Y2=3.145
r171 40 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.535 $Y=3.145
+ $X2=13.68 $Y2=3.145
r172 40 41 9.74008 $w=1.4e-07 $l=7.87e-06 $layer=MET1_cond $X=13.535 $Y=3.145
+ $X2=5.665 $Y2=3.145
r173 39 63 6.00569 $w=3.53e-07 $l=1.85e-07 $layer=LI1_cond $X=13.617 $Y=3.285
+ $X2=13.617 $Y2=3.1
r174 36 38 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=12.315 $Y=1.075
+ $X2=12.315 $Y2=1.245
r175 33 56 33.7946 $w=3.68e-07 $l=1.085e-06 $layer=LI1_cond $X=5.605 $Y=1.775
+ $X2=5.605 $Y2=2.86
r176 33 34 2.73602 $w=3.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=5.605 $Y=1.775
+ $X2=5.552 $Y2=1.69
r177 31 39 7.97992 $w=1.7e-07 $l=2.15346e-07 $layer=LI1_cond $X=13.44 $Y=3.37
+ $X2=13.617 $Y2=3.285
r178 31 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=13.44 $Y=3.37
+ $X2=12.48 $Y2=3.37
r179 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.395 $Y=3.285
+ $X2=12.48 $Y2=3.37
r180 30 38 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=12.395 $Y=3.285
+ $X2=12.395 $Y2=1.245
r181 27 52 6.95538 $w=5e-07 $l=6.5e-08 $layer=POLY_cond $X=6.955 $Y=1.645
+ $X2=7.02 $Y2=1.645
r182 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.955
+ $Y=1.69 $X2=6.955 $Y2=1.69
r183 24 34 4.03347 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=5.79 $Y=1.69
+ $X2=5.552 $Y2=1.69
r184 24 26 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=5.79 $Y=1.69
+ $X2=6.955 $Y2=1.69
r185 20 34 2.73602 $w=3.5e-07 $l=1.15521e-07 $layer=LI1_cond $X=5.48 $Y=1.605
+ $X2=5.552 $Y2=1.69
r186 20 22 31.6049 $w=3.28e-07 $l=9.05e-07 $layer=LI1_cond $X=5.48 $Y=1.605
+ $X2=5.48 $Y2=0.7
r187 16 53 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.39 $Y=1.895
+ $X2=7.39 $Y2=1.645
r188 16 18 129.477 $w=5e-07 $l=1.21e-06 $layer=POLY_cond $X=7.39 $Y=1.895
+ $X2=7.39 $Y2=3.105
r189 13 52 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.02 $Y=1.395
+ $X2=7.02 $Y2=1.645
r190 13 15 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.02 $Y=1.395 $X2=7.02
+ $Y2=1.075
r191 4 63 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=13.465
+ $Y=2.225 $X2=13.605 $Y2=3.1
r192 4 60 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=13.465
+ $Y=2.225 $X2=13.605 $Y2=2.35
r193 3 56 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=5.58
+ $Y=2.715 $X2=5.705 $Y2=2.86
r194 2 36 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=12.17
+ $Y=0.865 $X2=12.315 $Y2=1.075
r195 1 22 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=5.335
+ $Y=0.535 $X2=5.48 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1570_457# 1 2 9 14 15 17 18 20 21 23 24
+ 25 26 29 31 34 36 37 39 43 48 49 50 52 53 59 61 63 66 68 71 73 78 81 82
c187 81 0 1.08168e-19 $X=8.135 $Y=2.285
c188 73 0 1.52106e-19 $X=13.525 $Y=1.62
c189 66 0 1.6142e-19 $X=10.66 $Y=1.25
c190 25 0 3.19798e-19 $X=8.28 $Y=1.93
c191 24 0 1.93647e-20 $X=8.28 $Y=1.43
r192 83 85 34.554 $w=4.8e-07 $l=3.1e-07 $layer=POLY_cond $X=10.23 $Y=1.305
+ $X2=10.54 $Y2=1.305
r193 75 83 1.84115 $w=5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.23 $Y=1.545
+ $X2=10.23 $Y2=1.305
r194 71 90 3.3884 $w=5.69e-07 $l=4e-08 $layer=POLY_cond $X=13.445 $Y=1.755
+ $X2=13.485 $Y2=1.755
r195 71 88 19.4833 $w=5.69e-07 $l=2.3e-07 $layer=POLY_cond $X=13.445 $Y=1.755
+ $X2=13.215 $Y2=1.755
r196 70 73 4.0085 $w=2.28e-07 $l=8e-08 $layer=LI1_cond $X=13.445 $Y=1.62
+ $X2=13.525 $Y2=1.62
r197 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.445
+ $Y=1.62 $X2=13.445 $Y2=1.62
r198 66 85 13.3757 $w=4.8e-07 $l=1.2e-07 $layer=POLY_cond $X=10.66 $Y=1.305
+ $X2=10.54 $Y2=1.305
r199 65 68 8.61591 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.66 $Y=1.23
+ $X2=10.825 $Y2=1.23
r200 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.66
+ $Y=1.25 $X2=10.66 $Y2=1.25
r201 59 78 74.9041 $w=5e-07 $l=7e-07 $layer=POLY_cond $X=10.23 $Y=2.015
+ $X2=10.23 $Y2=2.715
r202 59 75 50.2928 $w=5e-07 $l=4.7e-07 $layer=POLY_cond $X=10.23 $Y=2.015
+ $X2=10.23 $Y2=1.545
r203 58 61 3.76308 $w=2.43e-07 $l=8e-08 $layer=LI1_cond $X=10.19 $Y=2.017
+ $X2=10.27 $Y2=2.017
r204 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.19
+ $Y=2.015 $X2=10.19 $Y2=2.015
r205 53 55 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.92 $Y=2.58
+ $X2=8.92 $Y2=2.835
r206 52 73 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=13.525 $Y=1.505
+ $X2=13.525 $Y2=1.62
r207 51 52 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=13.525 $Y=0.645
+ $X2=13.525 $Y2=1.505
r208 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.44 $Y=0.56
+ $X2=13.525 $Y2=0.645
r209 49 50 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=13.44 $Y=0.56
+ $X2=11.875 $Y2=0.56
r210 46 48 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=11.75 $Y=1.095
+ $X2=11.75 $Y2=0.745
r211 45 50 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=11.75 $Y=0.645
+ $X2=11.875 $Y2=0.56
r212 45 48 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=11.75 $Y=0.645
+ $X2=11.75 $Y2=0.745
r213 41 43 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=11.44 $Y=2.47
+ $X2=11.44 $Y2=2.485
r214 39 46 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=11.625 $Y=1.18
+ $X2=11.75 $Y2=1.095
r215 39 68 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=11.625 $Y=1.18
+ $X2=10.825 $Y2=1.18
r216 38 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.355 $Y=2.385
+ $X2=10.27 $Y2=2.385
r217 37 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=11.315 $Y=2.385
+ $X2=11.44 $Y2=2.47
r218 37 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.315 $Y=2.385
+ $X2=10.355 $Y2=2.385
r219 35 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.27 $Y=2.47
+ $X2=10.27 $Y2=2.385
r220 35 36 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.27 $Y=2.47
+ $X2=10.27 $Y2=2.75
r221 34 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.27 $Y=2.3
+ $X2=10.27 $Y2=2.385
r222 33 61 2.87745 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=10.27 $Y=2.14
+ $X2=10.27 $Y2=2.017
r223 33 34 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=10.27 $Y=2.14
+ $X2=10.27 $Y2=2.3
r224 32 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.005 $Y=2.835
+ $X2=8.92 $Y2=2.835
r225 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.185 $Y=2.835
+ $X2=10.27 $Y2=2.75
r226 31 32 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=10.185 $Y=2.835
+ $X2=9.005 $Y2=2.835
r227 29 82 21.1255 $w=5.7e-07 $l=2.15e-07 $layer=POLY_cond $X=8.135 $Y=2.57
+ $X2=8.135 $Y2=2.785
r228 29 81 27.696 $w=5.7e-07 $l=2.85e-07 $layer=POLY_cond $X=8.135 $Y=2.57
+ $X2=8.135 $Y2=2.285
r229 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.255
+ $Y=2.57 $X2=8.255 $Y2=2.57
r230 26 53 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.835 $Y=2.58
+ $X2=8.92 $Y2=2.58
r231 26 28 33.8565 $w=1.88e-07 $l=5.8e-07 $layer=LI1_cond $X=8.835 $Y=2.58
+ $X2=8.255 $Y2=2.58
r232 25 81 37.9871 $w=5e-07 $l=3.55e-07 $layer=POLY_cond $X=8.17 $Y=1.93
+ $X2=8.17 $Y2=2.285
r233 24 25 35.7064 $w=7.2e-07 $l=5e-07 $layer=POLY_cond $X=8.28 $Y=1.43 $X2=8.28
+ $Y2=1.93
r234 21 90 5.89942 $w=5e-07 $l=3.6e-07 $layer=POLY_cond $X=13.485 $Y=1.395
+ $X2=13.485 $Y2=1.755
r235 21 23 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=13.485 $Y=1.395
+ $X2=13.485 $Y2=1.075
r236 18 88 5.89942 $w=5e-07 $l=3.6e-07 $layer=POLY_cond $X=13.215 $Y=2.115
+ $X2=13.215 $Y2=1.755
r237 18 20 58.804 $w=5e-07 $l=6.1e-07 $layer=POLY_cond $X=13.215 $Y=2.115
+ $X2=13.215 $Y2=2.725
r238 15 85 1.84115 $w=5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.54 $Y=1.065
+ $X2=10.54 $Y2=1.305
r239 15 17 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.54 $Y=1.065
+ $X2=10.54 $Y2=0.745
r240 14 24 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.39 $Y=1.11 $X2=8.39
+ $Y2=1.43
r241 9 82 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.1 $Y=3.105 $X2=8.1
+ $Y2=2.785
r242 2 43 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=11.26
+ $Y=2.34 $X2=11.4 $Y2=2.485
r243 1 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.57
+ $Y=0.535 $X2=11.71 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1726_453# 1 2 9 13 15 17 20 25 31 33 34
+ 36 41 42 45 51 55
c105 55 0 1.52106e-19 $X=12.34 $Y=1.745
c106 36 0 4.27966e-19 $X=9.235 $Y=1.71
c107 13 0 1.09959e-19 $X=12.34 $Y=2.435
c108 9 0 1.50317e-20 $X=8.88 $Y=3.105
r109 46 55 32.2192 $w=5.61e-07 $l=3.75e-07 $layer=POLY_cond $X=11.965 $Y=1.745
+ $X2=12.34 $Y2=1.745
r110 45 48 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=11.965 $Y=1.56
+ $X2=11.965 $Y2=1.63
r111 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.965
+ $Y=1.56 $X2=11.965 $Y2=1.56
r112 41 42 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.84 $Y=2.485
+ $X2=9.84 $Y2=2.32
r113 37 51 64.2035 $w=5e-07 $l=6e-07 $layer=POLY_cond $X=9.17 $Y=1.71 $X2=9.17
+ $Y2=1.11
r114 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.235
+ $Y=1.71 $X2=9.235 $Y2=1.71
r115 33 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.8 $Y=1.63
+ $X2=11.965 $Y2=1.63
r116 33 34 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=11.8 $Y=1.63
+ $X2=10.315 $Y2=1.63
r117 29 34 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.15 $Y=1.63
+ $X2=10.315 $Y2=1.63
r118 29 38 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.15 $Y=1.63
+ $X2=9.76 $Y2=1.63
r119 29 31 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=10.15 $Y=1.545
+ $X2=10.15 $Y2=0.745
r120 27 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.76 $Y=1.715
+ $X2=9.76 $Y2=1.63
r121 27 42 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=9.76 $Y=1.715
+ $X2=9.76 $Y2=2.32
r122 26 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.4 $Y=1.63
+ $X2=9.235 $Y2=1.63
r123 25 38 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.675 $Y=1.63
+ $X2=9.76 $Y2=1.63
r124 25 26 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.675 $Y=1.63
+ $X2=9.4 $Y2=1.63
r125 21 37 59.3883 $w=5e-07 $l=5.55e-07 $layer=POLY_cond $X=9.17 $Y=2.265
+ $X2=9.17 $Y2=1.71
r126 20 21 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=9.17 $Y=2.515
+ $X2=9.17 $Y2=2.265
r127 18 20 31.0317 $w=5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.88 $Y=2.515
+ $X2=9.17 $Y2=2.515
r128 15 55 31.3601 $w=5.61e-07 $l=5.10857e-07 $layer=POLY_cond $X=12.705
+ $Y=1.395 $X2=12.34 $Y2=1.745
r129 15 17 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=12.705 $Y=1.395
+ $X2=12.705 $Y2=1.075
r130 11 55 5.56718 $w=5e-07 $l=3.5e-07 $layer=POLY_cond $X=12.34 $Y=2.095
+ $X2=12.34 $Y2=1.745
r131 11 13 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=12.34 $Y=2.095
+ $X2=12.34 $Y2=2.435
r132 7 18 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.88 $Y=2.765 $X2=8.88
+ $Y2=2.515
r133 7 9 36.382 $w=5e-07 $l=3.4e-07 $layer=POLY_cond $X=8.88 $Y=2.765 $X2=8.88
+ $Y2=3.105
r134 2 41 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=9.715
+ $Y=2.34 $X2=9.84 $Y2=2.485
r135 1 31 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=10.005
+ $Y=0.535 $X2=10.15 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%CLK 1 3 4 6 8 9
c40 9 0 1.09959e-19 $X=11.28 $Y=2.035
r41 13 16 7.61053 $w=4.75e-07 $l=6.5e-08 $layer=POLY_cond $X=10.945 $Y=1.992
+ $X2=11.01 $Y2=1.992
r42 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.945
+ $Y=2.01 $X2=10.945 $Y2=2.01
r43 9 14 17.1586 $w=2.23e-07 $l=3.35e-07 $layer=LI1_cond $X=11.28 $Y=2.007
+ $X2=10.945 $Y2=2.007
r44 8 14 7.42686 $w=2.23e-07 $l=1.45e-07 $layer=LI1_cond $X=10.8 $Y=2.007
+ $X2=10.945 $Y2=2.007
r45 4 16 36.2964 $w=4.75e-07 $l=3.1e-07 $layer=POLY_cond $X=11.32 $Y=1.992
+ $X2=11.01 $Y2=1.992
r46 4 6 108.076 $w=5e-07 $l=1.01e-06 $layer=POLY_cond $X=11.32 $Y=1.755
+ $X2=11.32 $Y2=0.745
r47 1 16 1.58534 $w=5e-07 $l=2.38e-07 $layer=POLY_cond $X=11.01 $Y=2.23
+ $X2=11.01 $Y2=1.992
r48 1 3 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.01 $Y=2.23 $X2=11.01
+ $Y2=2.715
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_2789_147# 1 2 9 11 13 16 20 24 28 30 33
+ 37 44 45 46 48 49 51 52 54 68
r110 67 68 25.6814 $w=5e-07 $l=2.4e-07 $layer=POLY_cond $X=17.405 $Y=1.665
+ $X2=17.645 $Y2=1.665
r111 63 65 27.8215 $w=5e-07 $l=2.6e-07 $layer=POLY_cond $X=16.51 $Y=1.665
+ $X2=16.77 $Y2=1.665
r112 58 60 39.5922 $w=5e-07 $l=3.7e-07 $layer=POLY_cond $X=14.195 $Y=2.355
+ $X2=14.565 $Y2=2.355
r113 55 67 55.108 $w=5e-07 $l=5.15e-07 $layer=POLY_cond $X=16.89 $Y=1.665
+ $X2=17.405 $Y2=1.665
r114 55 65 12.8407 $w=5e-07 $l=1.2e-07 $layer=POLY_cond $X=16.89 $Y=1.665
+ $X2=16.77 $Y2=1.665
r115 54 57 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=16.89 $Y=1.67
+ $X2=16.89 $Y2=1.835
r116 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.89
+ $Y=1.67 $X2=16.89 $Y2=1.67
r117 51 52 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=15.8 $Y=2.86
+ $X2=15.8 $Y2=2.695
r118 48 57 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=16.81 $Y=3.635
+ $X2=16.81 $Y2=1.835
r119 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=16.725 $Y=3.72
+ $X2=16.81 $Y2=3.635
r120 45 46 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=16.725 $Y=3.72
+ $X2=15.995 $Y2=3.72
r121 42 46 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=15.8 $Y=3.635
+ $X2=15.995 $Y2=3.72
r122 42 44 1.92074 $w=3.88e-07 $l=6.5e-08 $layer=LI1_cond $X=15.8 $Y=3.635
+ $X2=15.8 $Y2=3.57
r123 41 51 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=15.8 $Y=2.89
+ $X2=15.8 $Y2=2.86
r124 41 44 20.0939 $w=3.88e-07 $l=6.8e-07 $layer=LI1_cond $X=15.8 $Y=2.89
+ $X2=15.8 $Y2=3.57
r125 39 49 4.24487 $w=3.15e-07 $l=1.97864e-07 $layer=LI1_cond $X=15.69 $Y=2.515
+ $X2=15.545 $Y2=2.39
r126 39 52 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=15.69 $Y=2.515
+ $X2=15.69 $Y2=2.695
r127 35 49 4.24487 $w=3.15e-07 $l=1.25e-07 $layer=LI1_cond $X=15.545 $Y=2.265
+ $X2=15.545 $Y2=2.39
r128 35 37 41.7327 $w=4.58e-07 $l=1.605e-06 $layer=LI1_cond $X=15.545 $Y=2.265
+ $X2=15.545 $Y2=0.66
r129 33 60 6.95538 $w=5e-07 $l=6.5e-08 $layer=POLY_cond $X=14.63 $Y=2.355
+ $X2=14.565 $Y2=2.355
r130 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.63
+ $Y=2.39 $X2=14.63 $Y2=2.39
r131 30 49 2.18656 $w=2.5e-07 $l=2.3e-07 $layer=LI1_cond $X=15.315 $Y=2.39
+ $X2=15.545 $Y2=2.39
r132 30 32 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=15.315 $Y=2.39
+ $X2=14.63 $Y2=2.39
r133 26 68 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=17.645 $Y=1.915
+ $X2=17.645 $Y2=1.665
r134 26 28 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=17.645 $Y=1.915
+ $X2=17.645 $Y2=2.42
r135 22 67 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=17.405 $Y=1.415
+ $X2=17.405 $Y2=1.665
r136 22 24 71.6939 $w=5e-07 $l=6.7e-07 $layer=POLY_cond $X=17.405 $Y=1.415
+ $X2=17.405 $Y2=0.745
r137 18 65 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=16.77 $Y=1.915
+ $X2=16.77 $Y2=1.665
r138 18 20 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=16.77 $Y=1.915
+ $X2=16.77 $Y2=2.795
r139 14 63 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=16.51 $Y=1.415
+ $X2=16.51 $Y2=1.665
r140 14 16 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=16.51 $Y=1.415
+ $X2=16.51 $Y2=0.91
r141 11 60 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=14.565 $Y=2.605
+ $X2=14.565 $Y2=2.355
r142 11 13 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=14.565 $Y=2.605
+ $X2=14.565 $Y2=2.925
r143 7 58 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=14.195 $Y=2.105
+ $X2=14.195 $Y2=2.355
r144 7 9 110.216 $w=5e-07 $l=1.03e-06 $layer=POLY_cond $X=14.195 $Y=2.105
+ $X2=14.195 $Y2=1.075
r145 2 51 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.69
+ $Y=2.715 $X2=15.83 $Y2=2.86
r146 2 44 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=15.69
+ $Y=2.715 $X2=15.83 $Y2=3.57
r147 1 37 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=15.34
+ $Y=0.535 $X2=15.48 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_2518_445# 1 2 7 9 12 16 18 21 22 26 33
+ 38
r80 37 38 37.4521 $w=5e-07 $l=3.5e-07 $layer=POLY_cond $X=15.09 $Y=1.645
+ $X2=15.44 $Y2=1.645
r81 30 33 4.5451 $w=4.98e-07 $l=1.9e-07 $layer=LI1_cond $X=12.905 $Y=1.075
+ $X2=13.095 $Y2=1.075
r82 27 37 12.8407 $w=5e-07 $l=1.2e-07 $layer=POLY_cond $X=14.97 $Y=1.645
+ $X2=15.09 $Y2=1.645
r83 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.97
+ $Y=1.71 $X2=14.97 $Y2=1.71
r84 24 26 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=14.97 $Y=1.915
+ $X2=14.97 $Y2=1.71
r85 23 29 2.45823 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.99 $Y=2
+ $X2=12.825 $Y2=2
r86 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=14.805 $Y=2
+ $X2=14.97 $Y2=1.915
r87 22 23 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=14.805 $Y=2
+ $X2=12.99 $Y2=2
r88 21 29 5.36411 $w=2.28e-07 $l=1.18427e-07 $layer=LI1_cond $X=12.905 $Y=1.915
+ $X2=12.825 $Y2=2
r89 20 30 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=12.905 $Y=1.325
+ $X2=12.905 $Y2=1.075
r90 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.905 $Y=1.325
+ $X2=12.905 $Y2=1.915
r91 16 29 14.8553 $w=3.3e-07 $l=3.7e-07 $layer=LI1_cond $X=12.825 $Y=2.37
+ $X2=12.825 $Y2=2
r92 16 18 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=12.825 $Y=2.37
+ $X2=12.825 $Y2=3.02
r93 10 38 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=15.44 $Y=1.895
+ $X2=15.44 $Y2=1.645
r94 10 12 141.248 $w=5e-07 $l=1.32e-06 $layer=POLY_cond $X=15.44 $Y=1.895
+ $X2=15.44 $Y2=3.215
r95 7 37 2.83073 $w=5e-07 $l=2.5e-07 $layer=POLY_cond $X=15.09 $Y=1.395
+ $X2=15.09 $Y2=1.645
r96 7 9 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=15.09 $Y=1.395 $X2=15.09
+ $Y2=0.91
r97 2 18 600 $w=1.7e-07 $l=9.04903e-07 $layer=licon1_PDIFF $count=1 $X=12.59
+ $Y=2.225 $X2=12.825 $Y2=3.02
r98 2 16 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=12.59
+ $Y=2.225 $X2=12.825 $Y2=2.37
r99 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.955
+ $Y=0.865 $X2=13.095 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_3531_107# 1 2 9 13 17 21 25 27 28 32
r40 28 35 40.6478 $w=5.55e-07 $l=4.15e-07 $layer=POLY_cond $X=18.967 $Y=1.67
+ $X2=18.967 $Y2=2.085
r41 28 34 25.2235 $w=5.55e-07 $l=2.55e-07 $layer=POLY_cond $X=18.967 $Y=1.67
+ $X2=18.967 $Y2=1.415
r42 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=18.875
+ $Y=1.67 $X2=18.875 $Y2=1.67
r43 25 31 4.57321 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.2 $Y=1.67
+ $X2=18.115 $Y2=1.67
r44 25 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=18.2 $Y=1.67
+ $X2=18.875 $Y2=1.67
r45 23 31 2.16928 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.115 $Y=1.835
+ $X2=18.115 $Y2=1.67
r46 23 32 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=18.115 $Y=1.835
+ $X2=18.115 $Y2=2.025
r47 21 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=18.035 $Y=2.19
+ $X2=18.035 $Y2=2.025
r48 15 31 17.9908 $w=2.17e-07 $l=3.2e-07 $layer=LI1_cond $X=17.795 $Y=1.67
+ $X2=18.115 $Y2=1.67
r49 15 17 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=17.795 $Y=1.505
+ $X2=17.795 $Y2=0.745
r50 13 35 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=18.995 $Y=2.965
+ $X2=18.995 $Y2=2.085
r51 9 34 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=18.995 $Y=0.91
+ $X2=18.995 $Y2=1.415
r52 2 21 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=17.895
+ $Y=2.045 $X2=18.035 $Y2=2.19
r53 1 17 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=17.655
+ $Y=0.535 $X2=17.795 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%VPWR 1 2 3 4 5 6 7 22 25 32 46 50 57 68 77
+ 82
c129 82 0 1.87436e-19 $X=18.855 $Y=3.59
r130 80 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.855 $Y=3.59
+ $X2=18.855 $Y2=3.59
r131 77 80 25.3406 $w=5.88e-07 $l=1.25e-06 $layer=LI1_cond $X=18.675 $Y=2.34
+ $X2=18.675 $Y2=3.59
r132 74 82 0.500997 $w=3.7e-07 $l=1.305e-06 $layer=MET1_cond $X=17.55 $Y=3.63
+ $X2=18.855 $Y2=3.63
r133 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.55 $Y=3.59
+ $X2=17.55 $Y2=3.59
r134 71 73 11.9608 $w=5.88e-07 $l=5.9e-07 $layer=LI1_cond $X=17.37 $Y=3
+ $X2=17.37 $Y2=3.59
r135 68 71 16.4207 $w=5.88e-07 $l=8.1e-07 $layer=LI1_cond $X=17.37 $Y=2.19
+ $X2=17.37 $Y2=3
r136 65 74 0.85227 $w=3.7e-07 $l=2.22e-06 $layer=MET1_cond $X=15.33 $Y=3.63
+ $X2=17.55 $Y2=3.63
r137 63 65 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=14.61 $Y=3.63
+ $X2=15.33 $Y2=3.63
r138 62 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.33 $Y=3.59
+ $X2=15.33 $Y2=3.59
r139 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.61 $Y=3.59
+ $X2=14.61 $Y2=3.59
r140 60 62 5.05525 $w=9.03e-07 $l=3.75e-07 $layer=LI1_cond $X=14.972 $Y=3.215
+ $X2=14.972 $Y2=3.59
r141 57 60 4.78564 $w=9.03e-07 $l=3.55e-07 $layer=LI1_cond $X=14.972 $Y=2.86
+ $X2=14.972 $Y2=3.215
r142 54 63 1.38206 $w=3.7e-07 $l=3.6e-06 $layer=MET1_cond $X=11.01 $Y=3.63
+ $X2=14.61 $Y2=3.63
r143 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.01 $Y=3.59
+ $X2=11.01 $Y2=3.59
r144 50 53 14.1908 $w=5.88e-07 $l=7e-07 $layer=LI1_cond $X=10.83 $Y=2.89
+ $X2=10.83 $Y2=3.59
r145 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.125 $Y=3.59
+ $X2=7.125 $Y2=3.59
r146 42 47 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=6.405 $Y=3.63
+ $X2=7.125 $Y2=3.63
r147 41 46 28.6124 $w=2.88e-07 $l=7.2e-07 $layer=LI1_cond $X=6.405 $Y=3.61
+ $X2=7.125 $Y2=3.61
r148 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.405 $Y=3.59
+ $X2=6.405 $Y2=3.59
r149 38 42 1.46652 $w=3.7e-07 $l=3.82e-06 $layer=MET1_cond $X=2.585 $Y=3.63
+ $X2=6.405 $Y2=3.63
r150 36 38 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.865 $Y=3.63
+ $X2=2.585 $Y2=3.63
r151 35 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.585 $Y=3.59
+ $X2=2.585 $Y2=3.59
r152 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.865 $Y=3.59
+ $X2=1.865 $Y2=3.59
r153 32 35 1.09158 $w=9.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=3.505
+ $X2=2.225 $Y2=3.59
r154 29 36 0.291768 $w=3.7e-07 $l=7.6e-07 $layer=MET1_cond $X=1.105 $Y=3.63
+ $X2=1.865 $Y2=3.63
r155 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.105 $Y=3.59
+ $X2=1.105 $Y2=3.59
r156 25 28 16.3194 $w=5.88e-07 $l=8.05e-07 $layer=LI1_cond $X=0.925 $Y=2.785
+ $X2=0.925 $Y2=3.59
r157 22 54 0.449169 $w=3.7e-07 $l=1.17e-06 $layer=MET1_cond $X=9.84 $Y=3.63
+ $X2=11.01 $Y2=3.63
r158 22 47 1.0423 $w=3.7e-07 $l=2.715e-06 $layer=MET1_cond $X=9.84 $Y=3.63
+ $X2=7.125 $Y2=3.63
r159 7 80 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=18.46
+ $Y=2.215 $X2=18.605 $Y2=3.59
r160 7 77 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=18.46
+ $Y=2.215 $X2=18.605 $Y2=2.34
r161 6 71 300 $w=1.7e-07 $l=1.02261e-06 $layer=licon1_PDIFF $count=2 $X=17.02
+ $Y=2.045 $X2=17.16 $Y2=3
r162 6 68 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=17.02
+ $Y=2.045 $X2=17.16 $Y2=2.19
r163 5 60 300 $w=1.7e-07 $l=6.06218e-07 $layer=licon1_PDIFF $count=2 $X=14.815
+ $Y=2.715 $X2=15.05 $Y2=3.215
r164 5 57 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=14.815
+ $Y=2.715 $X2=15.05 $Y2=2.86
r165 4 50 600 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=1 $X=10.48
+ $Y=2.34 $X2=10.62 $Y2=2.89
r166 3 41 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=6.345
+ $Y=2.715 $X2=6.485 $Y2=3.57
r167 2 32 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.125
+ $Y=3.295 $X2=2.265 $Y2=3.505
r168 1 25 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.915
+ $Y=2.575 $X2=1.055 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_268_659# 1 2 9 11 12 15
c32 9 0 6.15916e-20 $X=1.485 $Y=3.505
r33 13 15 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=3.555 $Y=3.095
+ $X2=3.555 $Y2=3.2
r34 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.43 $Y=3.01
+ $X2=3.555 $Y2=3.095
r35 11 12 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=3.43 $Y=3.01
+ $X2=1.57 $Y2=3.01
r36 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.485 $Y=3.095
+ $X2=1.57 $Y2=3.01
r37 7 9 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.485 $Y=3.095
+ $X2=1.485 $Y2=3.505
r38 2 15 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=2.99 $X2=3.595 $Y2=3.2
r39 1 9 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=3.295 $X2=1.485 $Y2=3.505
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_581_659# 1 2 9 11 12 14 15 16 19
r46 17 19 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=5.115 $Y=2.85
+ $X2=5.115 $Y2=3.2
r47 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.99 $Y=2.765
+ $X2=5.115 $Y2=2.85
r48 15 16 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.99 $Y=2.765
+ $X2=4.03 $Y2=2.765
r49 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.945 $Y=2.85
+ $X2=4.03 $Y2=2.765
r50 13 14 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.945 $Y=2.85
+ $X2=3.945 $Y2=3.61
r51 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.86 $Y=3.695
+ $X2=3.945 $Y2=3.61
r52 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.86 $Y=3.695
+ $X2=3.21 $Y2=3.695
r53 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.045 $Y=3.61
+ $X2=3.21 $Y2=3.695
r54 7 9 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.045 $Y=3.61
+ $X2=3.045 $Y2=3.505
r55 2 19 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.015
+ $Y=2.99 $X2=5.155 $Y2=3.2
r56 1 9 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.905
+ $Y=3.295 $X2=3.045 $Y2=3.505
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_567_107# 1 2 3 4 13 16 17 18 21 23 24 26
+ 27 28 30 32 34 35 36 37 38 39 42 43 45 48 52 53 54 59 64
c189 59 0 4.11115e-20 $X=8 $Y=1.11
c190 42 0 1.93647e-20 $X=7.385 $Y=1.955
c191 28 0 7.37372e-20 $X=5.135 $Y=0.35
c192 13 0 3.21733e-20 $X=3.51 $Y=0.91
r193 64 66 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=9.27 $Y=3.185
+ $X2=9.27 $Y2=3.37
r194 59 61 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=8 $Y=1.11 $X2=8
+ $Y2=1.34
r195 54 56 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.475 $Y=3.2
+ $X2=7.475 $Y2=3.37
r196 48 50 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=0.745
+ $X2=2.975 $Y2=0.91
r197 46 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.56 $Y=3.37
+ $X2=7.475 $Y2=3.37
r198 45 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.105 $Y=3.37
+ $X2=9.27 $Y2=3.37
r199 45 46 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=9.105 $Y=3.37
+ $X2=7.56 $Y2=3.37
r200 44 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=1.34
+ $X2=7.385 $Y2=1.34
r201 43 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.835 $Y=1.34 $X2=8
+ $Y2=1.34
r202 43 44 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.835 $Y=1.34
+ $X2=7.47 $Y2=1.34
r203 41 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.385 $Y=1.425
+ $X2=7.385 $Y2=1.34
r204 41 42 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.385 $Y=1.425
+ $X2=7.385 $Y2=1.955
r205 40 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.14 $Y=3.2
+ $X2=6.055 $Y2=3.2
r206 39 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.39 $Y=3.2
+ $X2=7.475 $Y2=3.2
r207 39 40 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=7.39 $Y=3.2
+ $X2=6.14 $Y2=3.2
r208 37 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.3 $Y=2.04
+ $X2=7.385 $Y2=1.955
r209 37 38 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=7.3 $Y=2.04
+ $X2=6.14 $Y2=2.04
r210 35 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.3 $Y=1.34
+ $X2=7.385 $Y2=1.34
r211 35 36 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=7.3 $Y=1.34
+ $X2=5.995 $Y2=1.34
r212 33 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=3.285
+ $X2=6.055 $Y2=3.2
r213 33 34 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.055 $Y=3.285
+ $X2=6.055 $Y2=3.635
r214 32 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=3.115
+ $X2=6.055 $Y2=3.2
r215 31 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.055 $Y=2.125
+ $X2=6.14 $Y2=2.04
r216 31 32 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=6.055 $Y=2.125
+ $X2=6.055 $Y2=3.115
r217 30 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.91 $Y=1.255
+ $X2=5.995 $Y2=1.34
r218 29 30 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=5.91 $Y=0.435
+ $X2=5.91 $Y2=1.255
r219 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.825 $Y=0.35
+ $X2=5.91 $Y2=0.435
r220 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.825 $Y=0.35
+ $X2=5.135 $Y2=0.35
r221 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.05 $Y=0.435
+ $X2=5.135 $Y2=0.35
r222 25 26 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=5.05 $Y=0.435
+ $X2=5.05 $Y2=2.33
r223 23 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.97 $Y=3.72
+ $X2=6.055 $Y2=3.635
r224 23 24 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=5.97 $Y=3.72
+ $X2=4.54 $Y2=3.72
r225 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.375 $Y=3.635
+ $X2=4.54 $Y2=3.72
r226 19 21 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=4.375 $Y=3.635
+ $X2=4.375 $Y2=3.2
r227 17 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.965 $Y=2.415
+ $X2=5.05 $Y2=2.33
r228 17 18 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=4.965 $Y=2.415
+ $X2=3.68 $Y2=2.415
r229 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.595 $Y=2.33
+ $X2=3.68 $Y2=2.415
r230 15 16 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=3.595 $Y=0.995
+ $X2=3.595 $Y2=2.33
r231 14 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=0.91
+ $X2=2.975 $Y2=0.91
r232 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.51 $Y=0.91
+ $X2=3.595 $Y2=0.995
r233 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.51 $Y=0.91
+ $X2=3.14 $Y2=0.91
r234 4 64 600 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_PDIFF $count=1 $X=9.13
+ $Y=2.895 $X2=9.27 $Y2=3.185
r235 3 21 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.235
+ $Y=2.99 $X2=4.375 $Y2=3.2
r236 2 59 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.855
+ $Y=0.9 $X2=8 $Y2=1.11
r237 1 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.835
+ $Y=0.535 $X2=2.975 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_2365_445# 1 2 9 11 12 15
r39 13 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=14.175 $Y=3.635
+ $X2=14.175 $Y2=2.925
r40 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=14.01 $Y=3.72
+ $X2=14.175 $Y2=3.635
r41 11 12 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=14.01 $Y=3.72
+ $X2=12.115 $Y2=3.72
r42 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.95 $Y=3.635
+ $X2=12.115 $Y2=3.72
r43 7 9 41.907 $w=3.28e-07 $l=1.2e-06 $layer=LI1_cond $X=11.95 $Y=3.635
+ $X2=11.95 $Y2=2.435
r44 2 15 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=14.05
+ $Y=2.715 $X2=14.175 $Y2=2.925
r45 1 9 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=11.825
+ $Y=2.225 $X2=11.95 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%Q 1 2 9 11 12 13 14 24 39
r28 37 39 6.34654 $w=4.88e-07 $l=2.6e-07 $layer=LI1_cond $X=16.12 $Y=2.27
+ $X2=16.38 $Y2=2.27
r29 22 37 3.05139 $w=3.3e-07 $l=2.45e-07 $layer=LI1_cond $X=16.12 $Y=2.025
+ $X2=16.12 $Y2=2.27
r30 14 37 0.976391 $w=4.88e-07 $l=4e-08 $layer=LI1_cond $X=16.08 $Y=2.27
+ $X2=16.12 $Y2=2.27
r31 14 22 1.32706 $w=3.28e-07 $l=3.8e-08 $layer=LI1_cond $X=16.12 $Y=1.987
+ $X2=16.12 $Y2=2.025
r32 13 14 11.245 $w=3.28e-07 $l=3.22e-07 $layer=LI1_cond $X=16.12 $Y=1.665
+ $X2=16.12 $Y2=1.987
r33 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=16.12 $Y=1.295
+ $X2=16.12 $Y2=1.665
r34 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=16.12 $Y=0.925
+ $X2=16.12 $Y2=1.295
r35 11 24 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=16.12 $Y=0.925
+ $X2=16.12 $Y2=0.66
r36 7 39 3.05139 $w=3.3e-07 $l=2.45e-07 $layer=LI1_cond $X=16.38 $Y=2.515
+ $X2=16.38 $Y2=2.27
r37 7 9 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=16.38 $Y=2.515
+ $X2=16.38 $Y2=3.37
r38 2 39 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=16.255
+ $Y=2.045 $X2=16.38 $Y2=2.19
r39 2 9 300 $w=1.7e-07 $l=1.38609e-06 $layer=licon1_PDIFF $count=2 $X=16.255
+ $Y=2.045 $X2=16.38 $Y2=3.37
r40 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=15.975
+ $Y=0.535 $X2=16.12 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%Q_N 1 2 7 8 9 10 11 12 13 22
r13 13 40 15.3086 $w=3.33e-07 $l=4.45e-07 $layer=LI1_cond $X=19.387 $Y=3.145
+ $X2=19.387 $Y2=3.59
r14 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=19.387 $Y=2.775
+ $X2=19.387 $Y2=3.145
r15 11 12 14.9646 $w=3.33e-07 $l=4.35e-07 $layer=LI1_cond $X=19.387 $Y=2.34
+ $X2=19.387 $Y2=2.775
r16 10 11 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=19.387 $Y=2.035
+ $X2=19.387 $Y2=2.34
r17 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=19.387 $Y=1.665
+ $X2=19.387 $Y2=2.035
r18 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=19.387 $Y=1.295
+ $X2=19.387 $Y2=1.665
r19 7 8 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=19.387 $Y=0.925
+ $X2=19.387 $Y2=1.295
r20 7 22 9.11634 $w=3.33e-07 $l=2.65e-07 $layer=LI1_cond $X=19.387 $Y=0.925
+ $X2=19.387 $Y2=0.66
r21 2 40 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=19.245
+ $Y=2.215 $X2=19.385 $Y2=3.59
r22 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=19.245
+ $Y=2.215 $X2=19.385 $Y2=2.34
r23 1 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=19.245
+ $Y=0.535 $X2=19.385 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%VGND 1 2 3 4 5 6 7 22 25 34 43 52 61 72 83
+ 87
c110 87 0 1.6142e-19 $X=18.95 $Y=0.48
r111 84 87 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=18.23 $Y=0.44
+ $X2=18.95 $Y2=0.44
r112 83 89 2.44 $w=8.98e-07 $l=1.8e-07 $layer=LI1_cond $X=18.59 $Y=0.48
+ $X2=18.59 $Y2=0.66
r113 83 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=18.95 $Y=0.48
+ $X2=18.95 $Y2=0.48
r114 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=18.23 $Y=0.48
+ $X2=18.23 $Y2=0.48
r115 78 80 6.42105 $w=9.48e-07 $l=5e-07 $layer=LI1_cond $X=16.94 $Y=0.66
+ $X2=16.94 $Y2=1.16
r116 76 84 0.357032 $w=3.7e-07 $l=9.3e-07 $layer=MET1_cond $X=17.3 $Y=0.44
+ $X2=18.23 $Y2=0.44
r117 73 76 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=16.58 $Y=0.44
+ $X2=17.3 $Y2=0.44
r118 72 78 2.31158 $w=9.48e-07 $l=1.8e-07 $layer=LI1_cond $X=16.94 $Y=0.48
+ $X2=16.94 $Y2=0.66
r119 72 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=17.3 $Y=0.48
+ $X2=17.3 $Y2=0.48
r120 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=16.58 $Y=0.48
+ $X2=16.58 $Y2=0.48
r121 67 69 6.42105 $w=9.48e-07 $l=5e-07 $layer=LI1_cond $X=14.39 $Y=0.66
+ $X2=14.39 $Y2=1.16
r122 65 73 0.702547 $w=3.7e-07 $l=1.83e-06 $layer=MET1_cond $X=14.75 $Y=0.44
+ $X2=16.58 $Y2=0.44
r123 62 65 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=14.03 $Y=0.44
+ $X2=14.75 $Y2=0.44
r124 61 67 2.31158 $w=9.48e-07 $l=1.8e-07 $layer=LI1_cond $X=14.39 $Y=0.48
+ $X2=14.39 $Y2=0.66
r125 61 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.75 $Y=0.48
+ $X2=14.75 $Y2=0.48
r126 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.03 $Y=0.48
+ $X2=14.03 $Y2=0.48
r127 56 62 1.03654 $w=3.7e-07 $l=2.7e-06 $layer=MET1_cond $X=11.33 $Y=0.44
+ $X2=14.03 $Y2=0.44
r128 53 56 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=10.61 $Y=0.44
+ $X2=11.33 $Y2=0.44
r129 52 58 3.40316 $w=9.48e-07 $l=2.65e-07 $layer=LI1_cond $X=10.97 $Y=0.48
+ $X2=10.97 $Y2=0.745
r130 52 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.33 $Y=0.48
+ $X2=11.33 $Y2=0.48
r131 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.61 $Y=0.48
+ $X2=10.61 $Y2=0.48
r132 44 47 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=6.26 $Y=0.44
+ $X2=6.98 $Y2=0.44
r133 43 49 4.72921 $w=8.88e-07 $l=3.45e-07 $layer=LI1_cond $X=6.62 $Y=0.48
+ $X2=6.62 $Y2=0.825
r134 43 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.98 $Y=0.48
+ $X2=6.98 $Y2=0.48
r135 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.26 $Y=0.48
+ $X2=6.26 $Y2=0.48
r136 38 44 0.606571 $w=3.7e-07 $l=1.58e-06 $layer=MET1_cond $X=4.68 $Y=0.44
+ $X2=6.26 $Y2=0.44
r137 35 38 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=3.96 $Y=0.44
+ $X2=4.68 $Y2=0.44
r138 34 40 3.49514 $w=9.23e-07 $l=2.65e-07 $layer=LI1_cond $X=4.322 $Y=0.48
+ $X2=4.322 $Y2=0.745
r139 34 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.68 $Y=0.48
+ $X2=4.68 $Y2=0.48
r140 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.96 $Y=0.48
+ $X2=3.96 $Y2=0.48
r141 29 35 0.796604 $w=3.7e-07 $l=2.075e-06 $layer=MET1_cond $X=1.885 $Y=0.44
+ $X2=3.96 $Y2=0.44
r142 26 29 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=1.165 $Y=0.44
+ $X2=1.885 $Y2=0.44
r143 25 31 3.40316 $w=9.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.525 $Y=0.48
+ $X2=1.525 $Y2=0.745
r144 25 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.885 $Y=0.48
+ $X2=1.885 $Y2=0.48
r145 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.165 $Y=0.48
+ $X2=1.165 $Y2=0.48
r146 22 53 0.295607 $w=3.7e-07 $l=7.7e-07 $layer=MET1_cond $X=9.84 $Y=0.44
+ $X2=10.61 $Y2=0.44
r147 22 47 1.09797 $w=3.7e-07 $l=2.86e-06 $layer=MET1_cond $X=9.84 $Y=0.44
+ $X2=6.98 $Y2=0.44
r148 7 89 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=18.46
+ $Y=0.535 $X2=18.605 $Y2=0.66
r149 6 80 182 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_NDIFF $count=1 $X=16.76
+ $Y=0.535 $X2=16.9 $Y2=1.16
r150 6 78 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=16.76
+ $Y=0.535 $X2=16.9 $Y2=0.66
r151 5 69 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=14.445
+ $Y=0.865 $X2=14.7 $Y2=1.16
r152 5 67 182 $w=1.7e-07 $l=3.42491e-07 $layer=licon1_NDIFF $count=1 $X=14.445
+ $Y=0.865 $X2=14.7 $Y2=0.66
r153 4 58 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.79
+ $Y=0.535 $X2=10.93 $Y2=0.745
r154 3 49 182 $w=1.7e-07 $l=3.84578e-07 $layer=licon1_NDIFF $count=1 $X=6.12
+ $Y=0.535 $X2=6.34 $Y2=0.825
r155 2 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.325
+ $Y=0.535 $X2=4.465 $Y2=0.745
r156 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.345
+ $Y=0.535 $X2=1.485 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__SDFXBP_1%A_1454_173# 1 2 7 11 13
c30 7 0 8.01934e-20 $X=9.395 $Y=0.675
r31 13 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=7.41 $Y=0.675
+ $X2=7.41 $Y2=0.99
r32 9 11 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=9.56 $Y=0.76 $X2=9.56
+ $Y2=1.11
r33 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.575 $Y=0.675
+ $X2=7.41 $Y2=0.675
r34 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.395 $Y=0.675
+ $X2=9.56 $Y2=0.76
r35 7 8 118.738 $w=1.68e-07 $l=1.82e-06 $layer=LI1_cond $X=9.395 $Y=0.675
+ $X2=7.575 $Y2=0.675
r36 2 11 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.42
+ $Y=0.9 $X2=9.56 $Y2=1.11
r37 1 16 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=7.27
+ $Y=0.865 $X2=7.41 $Y2=0.99
.ends

