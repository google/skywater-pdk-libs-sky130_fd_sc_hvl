* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbuflv2hv_1 A LVPWR VGND VNB VPB VPWR X
X0 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X1 a_686_151# a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X2 a_1711_885# a_504_1221# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X3 a_1711_885# a_504_1221# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X4 a_404_1133# A a_686_151# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VPWR a_1711_885# X VPB sky130_fd_pr__pfet_g5v0d10v5 w=1.5e+06u l=500000u
X6 a_404_1133# A LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X7 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X8 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X9 a_1197_107# a_504_1221# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X10 a_686_151# a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X11 a_686_151# a_404_1133# a_772_151# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 LVPWR a_404_1133# a_772_151# LVPWR sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 a_686_151# a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X14 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X15 a_504_1221# a_1197_107# a_1606_563# VPB sky130_fd_pr__pfet_g5v0d10v5 w=420000u l=1e+06u
X16 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X17 VGND a_1711_885# X VNB sky130_fd_pr__nfet_g5v0d10v5 w=750000u l=500000u
X18 a_1197_107# a_772_151# a_686_151# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
X19 a_1197_107# a_772_151# a_686_151# VNB sky130_fd_pr__nfet_g5v0d10v5 w=1.5e+06u l=500000u
.ends
