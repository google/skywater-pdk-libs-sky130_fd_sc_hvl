# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__mux2_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__mux2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A0
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 1.785000 2.905000 1.955000 ;
        RECT 2.295000 1.955000 2.625000 2.235000 ;
        RECT 2.735000 1.095000 3.685000 1.390000 ;
        RECT 2.735000 1.390000 2.905000 1.785000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.085000 1.570000 3.685000 1.955000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 1.705000 1.765000 3.095000 ;
        RECT 1.435000 3.095000 3.230000 3.265000 ;
        RECT 3.060000 2.135000 4.675000 2.305000 ;
        RECT 3.060000 2.305000 3.230000 3.095000 ;
        RECT 4.365000 1.550000 4.675000 2.135000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.495000 0.415000 1.925000 ;
        RECT 0.125000 1.925000 0.495000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 5.280000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 5.280000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 5.280000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 5.280000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.985000 5.280000 4.155000 ;
      RECT 0.595000  0.365000 2.205000 1.175000 ;
      RECT 0.620000  1.355000 2.555000 1.525000 ;
      RECT 0.620000  1.525000 0.950000 1.745000 ;
      RECT 0.675000  2.175000 1.255000 3.755000 ;
      RECT 1.945000  1.525000 2.115000 2.415000 ;
      RECT 1.945000  2.415000 2.880000 2.585000 ;
      RECT 2.385000  0.495000 2.880000 0.915000 ;
      RECT 2.385000  0.915000 2.555000 1.355000 ;
      RECT 2.550000  2.585000 2.880000 2.915000 ;
      RECT 3.060000  0.365000 4.720000 0.915000 ;
      RECT 3.410000  2.495000 4.720000 3.705000 ;
      RECT 3.865000  1.105000 5.150000 1.275000 ;
      RECT 3.865000  1.275000 4.115000 1.775000 ;
      RECT 4.900000  0.495000 5.150000 1.105000 ;
      RECT 4.900000  1.275000 5.150000 2.915000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.595000  0.395000 0.765000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.700000  3.505000 0.870000 3.675000 ;
      RECT 0.955000  0.395000 1.125000 0.565000 ;
      RECT 1.060000  3.505000 1.230000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.315000  0.395000 1.485000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.675000  0.395000 1.845000 0.565000 ;
      RECT 2.035000  0.395000 2.205000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.085000  0.395000 3.255000 0.565000 ;
      RECT 3.440000  3.505000 3.610000 3.675000 ;
      RECT 3.445000  0.395000 3.615000 0.565000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.800000  3.505000 3.970000 3.675000 ;
      RECT 3.805000  0.395000 3.975000 0.565000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.160000  3.505000 4.330000 3.675000 ;
      RECT 4.165000  0.395000 4.335000 0.565000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.520000  3.505000 4.690000 3.675000 ;
      RECT 4.525000  0.395000 4.695000 0.565000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
  END
END sky130_fd_sc_hvl__mux2_1
END LIBRARY
