* File: sky130_fd_sc_hvl__lsbufhv2lv_simple_1.pxi.spice
* Created: Wed Sep  2 09:07:35 2020
* 
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%VNB N_VNB_M0_noxref_b VNB VNB
+ N_VNB_c_9_p VNB PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%VNB
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%VPB N_VPB_X4_noxref_D1
+ N_VPB_X6_noxref_D1 VPB N_VPB_c_26_n N_VPB_c_27_n N_VPB_c_28_n
+ PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%VPB
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%LVPWR N_LVPWR_M1001_d N_LVPWR_M1001_b
+ N_LVPWR_c_47_n N_LVPWR_c_48_n LVPWR N_LVPWR_c_54_p
+ PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%LVPWR
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%A_662_81# N_A_662_81#_M1_noxref_d
+ N_A_662_81#_M1003_d N_A_662_81#_M0_noxref_g N_A_662_81#_M1001_g
+ N_A_662_81#_c_80_n N_A_662_81#_c_81_n N_A_662_81#_c_82_n N_A_662_81#_c_115_p
+ N_A_662_81#_c_83_n N_A_662_81#_c_85_n N_A_662_81#_c_86_n N_A_662_81#_c_87_n
+ PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%A_662_81#
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%A A A A A A N_A_M1_noxref_g
+ N_A_c_132_n N_A_M1003_g PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%A
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%X N_X_M0_noxref_s N_X_M1001_s X X X X
+ X X X N_X_c_150_n X N_X_c_157_n PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%X
x_PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%VGND N_VGND_M0_noxref_d VGND VGND
+ N_VGND_c_171_n N_VGND_c_173_n PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%VGND
cc_1 N_VNB_M0_noxref_b N_VPB_c_26_n 0.0021751f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_2 N_VNB_M0_noxref_b N_VPB_c_27_n 0.0021751f $X=-0.33 $Y=-0.265 $X2=8.4
+ $Y2=4.07
cc_3 N_VNB_M0_noxref_b N_VPB_c_28_n 0.0830934f $X=-0.33 $Y=-0.265 $X2=8.4
+ $Y2=4.07
cc_4 N_VNB_M0_noxref_b LVPWR 0.211657f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_5 N_VNB_M0_noxref_b N_A_662_81#_c_80_n 0.00140289f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_6 N_VNB_M0_noxref_b N_A_662_81#_c_81_n 0.0581956f $X=-0.33 $Y=-0.265 $X2=0.24
+ $Y2=4.07
cc_7 N_VNB_M0_noxref_b N_A_662_81#_c_82_n 0.0121633f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_8 N_VNB_M0_noxref_b N_A_662_81#_c_83_n 0.0310211f $X=-0.33 $Y=-0.265 $X2=8.4
+ $Y2=4.07
cc_9 N_VNB_c_9_p N_A_662_81#_c_83_n 5.81195e-19 $X=0.24 $Y=0 $X2=8.4 $Y2=4.07
cc_10 N_VNB_M0_noxref_b N_A_662_81#_c_85_n 0.030449f $X=-0.33 $Y=-0.265 $X2=4.32
+ $Y2=4.07
cc_11 N_VNB_M0_noxref_b N_A_662_81#_c_86_n 0.00770964f $X=-0.33 $Y=-0.265
+ $X2=8.4 $Y2=4.07
cc_12 N_VNB_M0_noxref_b N_A_662_81#_c_87_n 0.0441687f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_c_9_p N_A_662_81#_c_87_n 5.86481e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_14 N_VNB_M0_noxref_b N_A_M1_noxref_g 0.128583f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_15 N_VNB_c_9_p N_A_M1_noxref_g 5.86481e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_16 N_VNB_M0_noxref_b N_X_c_150_n 0.0685484f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_17 N_VNB_c_9_p N_X_c_150_n 6.04631e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_18 N_VNB_M0_noxref_b VGND 0.545305f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_19 VNB VGND 0.925009f $X=0 $Y=8.025 $X2=0 $Y2=0
cc_20 N_VNB_M0_noxref_b N_VGND_c_171_n 0.0622807f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_21 N_VNB_c_9_p N_VGND_c_171_n 0.0035518f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_22 N_VNB_M0_noxref_b N_VGND_c_173_n 0.437531f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_23 N_VNB_c_9_p N_VGND_c_173_n 0.924731f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_24 N_VNB_M0_noxref_b VPWR 0.098711f $X=-0.33 $Y=-0.265 $X2=0 $Y2=3.985
cc_25 N_VNB_M0_noxref_b VPWR 0.224313f $X=-0.33 $Y=-0.265 $X2=7.755 $Y2=3.985
cc_26 N_VPB_c_28_n N_LVPWR_M1001_b 0.0212813f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_27 N_VPB_c_28_n N_LVPWR_c_47_n 0.0587624f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_28 N_VPB_c_28_n N_LVPWR_c_48_n 0.0557866f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_29 N_VPB_X4_noxref_D1 LVPWR 0.050189f $X=-0.33 $Y=1.885 $X2=0.24 $Y2=0
cc_30 N_VPB_X6_noxref_D1 LVPWR 0.0721485f $X=7.425 $Y=1.885 $X2=0.24 $Y2=0
cc_31 N_VPB_c_28_n X 0.00120061f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_32 N_VPB_X4_noxref_D1 VPWR 0.0336658f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_33 N_VPB_X6_noxref_D1 VPWR 0.0422033f $X=7.425 $Y=1.885 $X2=0 $Y2=0
cc_34 N_VPB_c_26_n VPWR 0.00613319f $X=0.24 $Y=4.07 $X2=0 $Y2=0
cc_35 N_VPB_c_27_n VPWR 0.00931478f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_36 N_VPB_c_28_n VPWR 0.916941f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_37 N_VPB_X4_noxref_D1 VPWR 0.0565882f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_38 N_VPB_X6_noxref_D1 VPWR 0.078157f $X=7.425 $Y=1.885 $X2=0 $Y2=0
cc_39 N_VPB_c_26_n VPWR 0.00613319f $X=0.24 $Y=4.07 $X2=0 $Y2=0
cc_40 N_VPB_c_27_n VPWR 0.00931478f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_41 N_VPB_c_28_n VPWR 0.903541f $X=8.4 $Y=4.07 $X2=0 $Y2=0
cc_42 N_LVPWR_M1001_b N_A_662_81#_M1001_g 0.0612552f $X=2.8 $Y=1.885 $X2=0
+ $Y2=8.025
cc_43 N_LVPWR_c_48_n N_A_662_81#_M1001_g 0.00855416f $X=3.897 $Y=3.955 $X2=0
+ $Y2=8.025
cc_44 LVPWR N_A_662_81#_M1001_g 0.00959355f $X=0.07 $Y=3.02 $X2=0 $Y2=8.025
cc_45 N_LVPWR_c_54_p N_A_662_81#_M1001_g 0.0868446f $X=4.055 $Y=2.34 $X2=0
+ $Y2=8.025
cc_46 N_LVPWR_c_54_p N_A_662_81#_c_80_n 0.0107918f $X=4.055 $Y=2.34 $X2=0.24
+ $Y2=0
cc_47 N_LVPWR_M1001_b N_A_662_81#_c_81_n 0.00408238f $X=2.8 $Y=1.885 $X2=0.24
+ $Y2=0
cc_48 N_LVPWR_M1001_b N_A_662_81#_c_85_n 0.0493968f $X=2.8 $Y=1.885 $X2=0 $Y2=0
cc_49 LVPWR N_A_662_81#_c_85_n 0.0162923f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_50 N_LVPWR_M1001_b N_A_M1_noxref_g 0.0623628f $X=2.8 $Y=1.885 $X2=0 $Y2=8.025
cc_51 LVPWR N_A_M1_noxref_g 0.0114705f $X=0.07 $Y=3.02 $X2=0 $Y2=8.025
cc_52 N_LVPWR_c_54_p N_A_M1_noxref_g 0.00863521f $X=4.055 $Y=2.34 $X2=0
+ $Y2=8.025
cc_53 N_LVPWR_M1001_b N_A_c_132_n 0.00696568f $X=2.8 $Y=1.885 $X2=0.24 $Y2=0
cc_54 LVPWR N_A_c_132_n 0.0443244f $X=0.07 $Y=3.02 $X2=0.24 $Y2=0
cc_55 N_LVPWR_c_54_p N_A_c_132_n 0.0813128f $X=4.055 $Y=2.34 $X2=0.24 $Y2=0
cc_56 N_LVPWR_M1001_b N_X_c_150_n 0.0159909f $X=2.8 $Y=1.885 $X2=0 $Y2=0
cc_57 N_LVPWR_M1001_b X 0.0468726f $X=2.8 $Y=1.885 $X2=0 $Y2=0
cc_58 N_LVPWR_c_48_n X 0.0194349f $X=3.897 $Y=3.955 $X2=0 $Y2=0
cc_59 LVPWR X 0.057874f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_60 N_LVPWR_M1001_b N_X_c_157_n 0.0133803f $X=2.8 $Y=1.885 $X2=0 $Y2=0
cc_61 N_LVPWR_c_54_p N_X_c_157_n 0.1117f $X=4.055 $Y=2.34 $X2=0 $Y2=0
cc_62 N_LVPWR_M1001_d VPWR 2.10522e-19 $X=3.915 $Y=2.215 $X2=0 $Y2=0
cc_63 N_LVPWR_M1001_b VPWR 0.0293317f $X=2.8 $Y=1.885 $X2=0 $Y2=0
cc_64 N_LVPWR_c_47_n VPWR 0.00738401f $X=4.89 $Y=4.07 $X2=0 $Y2=0
cc_65 N_LVPWR_c_48_n VPWR 0.00252876f $X=3.897 $Y=3.955 $X2=0 $Y2=0
cc_66 LVPWR VPWR 0.912095f $X=0.07 $Y=3.02 $X2=0 $Y2=0
cc_67 N_LVPWR_c_54_p VPWR 0.0545982f $X=4.055 $Y=2.34 $X2=0 $Y2=0
cc_68 N_LVPWR_M1001_b VPWR 0.115262f $X=2.8 $Y=1.885 $X2=0 $Y2=0
cc_69 N_LVPWR_c_47_n VPWR 0.0642888f $X=4.89 $Y=4.07 $X2=0 $Y2=0
cc_70 N_LVPWR_c_48_n VPWR 0.0722445f $X=3.897 $Y=3.955 $X2=0 $Y2=0
cc_71 N_A_662_81#_c_80_n N_A_M1_noxref_g 0.00392032f $X=3.73 $Y=1.58 $X2=0
+ $Y2=8.025
cc_72 N_A_662_81#_c_81_n N_A_M1_noxref_g 0.041181f $X=3.73 $Y=1.58 $X2=0
+ $Y2=8.025
cc_73 N_A_662_81#_c_82_n N_A_M1_noxref_g 0.034515f $X=4.865 $Y=1.2 $X2=0
+ $Y2=8.025
cc_74 N_A_662_81#_c_83_n N_A_M1_noxref_g 0.0090774f $X=4.95 $Y=0.745 $X2=0
+ $Y2=8.025
cc_75 N_A_662_81#_c_85_n N_A_M1_noxref_g 0.0335927f $X=4.95 $Y=2.34 $X2=0
+ $Y2=8.025
cc_76 N_A_662_81#_c_87_n N_A_M1_noxref_g 0.0184277f $X=3.612 $Y=1.395 $X2=0
+ $Y2=8.025
cc_77 N_A_662_81#_M1001_g N_A_c_132_n 3.29035e-19 $X=3.665 $Y=2.965 $X2=0.24
+ $Y2=0
cc_78 N_A_662_81#_c_80_n N_A_c_132_n 0.00936991f $X=3.73 $Y=1.58 $X2=0.24 $Y2=0
cc_79 N_A_662_81#_c_81_n N_A_c_132_n 0.00392409f $X=3.73 $Y=1.58 $X2=0.24 $Y2=0
cc_80 N_A_662_81#_c_82_n N_A_c_132_n 0.0238596f $X=4.865 $Y=1.2 $X2=0.24 $Y2=0
cc_81 N_A_662_81#_c_85_n N_A_c_132_n 0.0853873f $X=4.95 $Y=2.34 $X2=0.24 $Y2=0
cc_82 N_A_662_81#_M1001_g N_X_c_150_n 0.0116649f $X=3.665 $Y=2.965 $X2=0 $Y2=0
cc_83 N_A_662_81#_c_80_n N_X_c_150_n 0.0227476f $X=3.73 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A_662_81#_c_87_n N_X_c_150_n 0.0243181f $X=3.612 $Y=1.395 $X2=0 $Y2=0
cc_85 N_A_662_81#_M1001_g X 0.0215851f $X=3.665 $Y=2.965 $X2=0 $Y2=0
cc_86 N_A_662_81#_M1001_g N_X_c_157_n 0.00584083f $X=3.665 $Y=2.965 $X2=0 $Y2=0
cc_87 N_A_662_81#_c_81_n N_X_c_157_n 0.0045161f $X=3.73 $Y=1.58 $X2=0 $Y2=0
cc_88 N_A_662_81#_c_82_n N_VGND_M0_noxref_d 0.00985042f $X=4.865 $Y=1.2 $X2=0
+ $Y2=0
cc_89 N_A_662_81#_c_115_p N_VGND_M0_noxref_d 2.97932e-19 $X=3.895 $Y=1.2 $X2=0
+ $Y2=0
cc_90 N_A_662_81#_c_81_n N_VGND_c_171_n 3.04803e-19 $X=3.73 $Y=1.58 $X2=-0.33
+ $Y2=-0.265
cc_91 N_A_662_81#_c_82_n N_VGND_c_171_n 0.0543159f $X=4.865 $Y=1.2 $X2=-0.33
+ $Y2=-0.265
cc_92 N_A_662_81#_c_115_p N_VGND_c_171_n 0.0208495f $X=3.895 $Y=1.2 $X2=-0.33
+ $Y2=-0.265
cc_93 N_A_662_81#_c_83_n N_VGND_c_171_n 0.0192683f $X=4.95 $Y=0.745 $X2=-0.33
+ $Y2=-0.265
cc_94 N_A_662_81#_c_87_n N_VGND_c_171_n 0.0421821f $X=3.612 $Y=1.395 $X2=-0.33
+ $Y2=-0.265
cc_95 N_A_662_81#_M1_noxref_d N_VGND_c_173_n 6.76135e-19 $X=4.81 $Y=0.535 $X2=0
+ $Y2=0
cc_96 N_A_662_81#_c_82_n N_VGND_c_173_n 0.008626f $X=4.865 $Y=1.2 $X2=0 $Y2=0
cc_97 N_A_662_81#_c_115_p N_VGND_c_173_n 0.00135661f $X=3.895 $Y=1.2 $X2=0 $Y2=0
cc_98 N_A_662_81#_c_83_n N_VGND_c_173_n 0.0275143f $X=4.95 $Y=0.745 $X2=0 $Y2=0
cc_99 N_A_662_81#_c_87_n N_VGND_c_173_n 0.00910554f $X=3.612 $Y=1.395 $X2=0
+ $Y2=0
cc_100 N_A_662_81#_M1001_g VPWR 0.00308323f $X=3.665 $Y=2.965 $X2=0 $Y2=0
cc_101 N_A_M1_noxref_g N_VGND_c_171_n 0.0443101f $X=4.56 $Y=0.745 $X2=-0.33
+ $Y2=-0.265
cc_102 N_A_M1_noxref_g N_VGND_c_173_n 0.00552997f $X=4.56 $Y=0.745 $X2=0 $Y2=0
cc_103 N_A_M1_noxref_g VPWR 7.73971e-19 $X=4.56 $Y=0.745 $X2=0 $Y2=0
cc_104 N_A_c_132_n VPWR 0.00226714f $X=4.52 $Y=1.55 $X2=0 $Y2=0
cc_105 N_X_c_150_n N_VGND_c_171_n 0.0192718f $X=3.17 $Y=0.68 $X2=-0.33
+ $Y2=-0.265
cc_106 N_X_M0_noxref_s N_VGND_c_173_n 0.00221032f $X=3.045 $Y=0.535 $X2=0 $Y2=0
cc_107 N_X_c_150_n N_VGND_c_173_n 0.0283937f $X=3.17 $Y=0.68 $X2=0 $Y2=0
cc_108 X VPWR 0.0394062f $X=3.12 $Y=2.405 $X2=0 $Y2=0
