# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hvl__buf_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hvl__buf_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.775000 4.215000 2.120000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.260000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.550000 1.390000 1.780000 ;
        RECT 1.220000 0.495000 1.470000 1.205000 ;
        RECT 1.220000 1.205000 3.030000 1.375000 ;
        RECT 1.220000 1.375000 1.390000 1.550000 ;
        RECT 1.220000 1.780000 1.390000 1.905000 ;
        RECT 1.220000 1.905000 3.110000 2.075000 ;
        RECT 1.220000 2.075000 1.470000 3.755000 ;
        RECT 2.780000 0.495000 3.030000 1.205000 ;
        RECT 2.780000 2.075000 3.110000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 4.800000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 4.800000 0.115000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 4.800000 4.185000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 4.800000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.985000 4.800000 4.155000 ;
      RECT 0.090000  0.365000 1.040000 1.325000 ;
      RECT 0.090000  2.175000 1.040000 3.755000 ;
      RECT 1.570000  1.555000 4.670000 1.595000 ;
      RECT 1.570000  1.595000 3.600000 1.725000 ;
      RECT 1.650000  0.365000 2.600000 1.025000 ;
      RECT 1.650000  2.255000 2.600000 3.755000 ;
      RECT 3.210000  0.365000 4.160000 1.245000 ;
      RECT 3.290000  2.300000 4.240000 3.755000 ;
      RECT 3.430000  1.425000 4.670000 1.555000 ;
      RECT 4.340000  0.495000 4.670000 1.425000 ;
      RECT 4.420000  1.595000 4.670000 3.755000 ;
    LAYER mcon ;
      RECT 0.120000  0.395000 0.290000 0.565000 ;
      RECT 0.120000  3.505000 0.290000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.480000  0.395000 0.650000 0.565000 ;
      RECT 0.480000  3.505000 0.650000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.840000  0.395000 1.010000 0.565000 ;
      RECT 0.840000  3.505000 1.010000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.680000  0.395000 1.850000 0.565000 ;
      RECT 1.680000  3.505000 1.850000 3.675000 ;
      RECT 2.040000  0.395000 2.210000 0.565000 ;
      RECT 2.040000  3.505000 2.210000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.400000  0.395000 2.570000 0.565000 ;
      RECT 2.400000  3.505000 2.570000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.240000  0.395000 3.410000 0.565000 ;
      RECT 3.320000  3.505000 3.490000 3.675000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.600000  0.395000 3.770000 0.565000 ;
      RECT 3.680000  3.505000 3.850000 3.675000 ;
      RECT 3.960000  0.395000 4.130000 0.565000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.040000  3.505000 4.210000 3.675000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
  END
END sky130_fd_sc_hvl__buf_4
