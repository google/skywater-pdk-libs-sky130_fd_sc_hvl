* File: sky130_fd_sc_hvl__buf_2.pxi.spice
* Created: Wed Sep  2 09:04:05 2020
* 
x_PM_SKY130_FD_SC_HVL__BUF_2%VNB N_VNB_M1002_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__BUF_2%VNB
x_PM_SKY130_FD_SC_HVL__BUF_2%VPB N_VPB_M1001_b VPB N_VPB_c_24_p VPB
+ PM_SKY130_FD_SC_HVL__BUF_2%VPB
x_PM_SKY130_FD_SC_HVL__BUF_2%A_129_279# N_A_129_279#_M1004_d
+ N_A_129_279#_M1000_d N_A_129_279#_c_54_n N_A_129_279#_M1001_g
+ N_A_129_279#_c_45_n N_A_129_279#_M1002_g N_A_129_279#_M1003_g
+ N_A_129_279#_c_47_n N_A_129_279#_M1005_g N_A_129_279#_c_49_n
+ N_A_129_279#_c_50_n N_A_129_279#_c_51_n N_A_129_279#_c_69_p
+ N_A_129_279#_c_52_n N_A_129_279#_c_53_n PM_SKY130_FD_SC_HVL__BUF_2%A_129_279#
x_PM_SKY130_FD_SC_HVL__BUF_2%A N_A_M1000_g N_A_M1004_g A A N_A_c_102_n
+ N_A_c_103_n N_A_c_106_n PM_SKY130_FD_SC_HVL__BUF_2%A
x_PM_SKY130_FD_SC_HVL__BUF_2%VPWR N_VPWR_M1001_s N_VPWR_M1003_s VPWR
+ N_VPWR_c_125_n N_VPWR_c_128_n N_VPWR_c_131_n PM_SKY130_FD_SC_HVL__BUF_2%VPWR
x_PM_SKY130_FD_SC_HVL__BUF_2%X N_X_M1002_d N_X_M1001_d N_X_c_152_n N_X_c_149_n X
+ X X PM_SKY130_FD_SC_HVL__BUF_2%X
x_PM_SKY130_FD_SC_HVL__BUF_2%VGND N_VGND_M1002_s N_VGND_M1005_s VGND
+ N_VGND_c_175_n N_VGND_c_177_n N_VGND_c_179_n PM_SKY130_FD_SC_HVL__BUF_2%VGND
cc_1 N_VNB_M1002_b N_A_129_279#_c_45_n 0.0444239f $X=-0.33 $Y=-0.265 $X2=0.915
+ $Y2=1.395
cc_2 N_VNB_c_2_p N_A_129_279#_c_45_n 5.86481e-19 $X=0.24 $Y=0 $X2=0.915
+ $Y2=1.395
cc_3 N_VNB_M1002_b N_A_129_279#_c_47_n 0.0426704f $X=-0.33 $Y=-0.265 $X2=1.695
+ $Y2=1.395
cc_4 N_VNB_c_2_p N_A_129_279#_c_47_n 5.86481e-19 $X=0.24 $Y=0 $X2=1.695
+ $Y2=1.395
cc_5 N_VNB_M1002_b N_A_129_279#_c_49_n 0.0145627f $X=-0.33 $Y=-0.265 $X2=2.98
+ $Y2=1.51
cc_6 N_VNB_M1002_b N_A_129_279#_c_50_n 0.0148195f $X=-0.33 $Y=-0.265 $X2=3.065
+ $Y2=2.34
cc_7 N_VNB_M1002_b N_A_129_279#_c_51_n 0.0280653f $X=-0.33 $Y=-0.265 $X2=3.085
+ $Y2=1.075
cc_8 N_VNB_M1002_b N_A_129_279#_c_52_n 0.00852418f $X=-0.33 $Y=-0.265 $X2=3.115
+ $Y2=1.51
cc_9 N_VNB_M1002_b N_A_129_279#_c_53_n 0.103893f $X=-0.33 $Y=-0.265 $X2=1.695
+ $Y2=1.75
cc_10 N_VNB_M1002_b A 0.00545491f $X=-0.33 $Y=-0.265 $X2=0.895 $Y2=2.965
cc_11 N_VNB_M1002_b N_A_c_102_n 0.0512249f $X=-0.33 $Y=-0.265 $X2=0.915 $Y2=0.91
cc_12 N_VNB_M1002_b N_A_c_103_n 0.0454459f $X=-0.33 $Y=-0.265 $X2=1.675
+ $Y2=2.965
cc_13 N_VNB_M1002_b N_X_c_149_n 0.00827821f $X=-0.33 $Y=-0.265 $X2=1.675
+ $Y2=2.965
cc_14 N_VNB_c_2_p N_X_c_149_n 3.93713e-19 $X=0.24 $Y=0 $X2=1.675 $Y2=2.965
cc_15 N_VNB_M1002_b X 0.0242117f $X=-0.33 $Y=-0.265 $X2=1.695 $Y2=0.91
cc_16 N_VNB_M1002_b N_VGND_c_175_n 0.0961733f $X=-0.33 $Y=-0.265 $X2=0.915
+ $Y2=1.395
cc_17 N_VNB_c_2_p N_VGND_c_175_n 0.00269049f $X=0.24 $Y=0 $X2=0.915 $Y2=1.395
cc_18 N_VNB_M1002_b N_VGND_c_177_n 0.0738976f $X=-0.33 $Y=-0.265 $X2=1.695
+ $Y2=0.91
cc_19 N_VNB_c_2_p N_VGND_c_177_n 0.00354191f $X=0.24 $Y=0 $X2=1.695 $Y2=0.91
cc_20 N_VNB_M1002_b N_VGND_c_179_n 0.0782508f $X=-0.33 $Y=-0.265 $X2=3.115
+ $Y2=2.34
cc_21 N_VNB_c_2_p N_VGND_c_179_n 0.359281f $X=0.24 $Y=0 $X2=3.115 $Y2=2.34
cc_22 N_VPB_M1001_b N_A_129_279#_c_54_n 0.0387543f $X=-0.33 $Y=1.885 $X2=0.895
+ $Y2=2.105
cc_23 VPB N_A_129_279#_c_54_n 0.00970178f $X=0 $Y=3.955 $X2=0.895 $Y2=2.105
cc_24 N_VPB_c_24_p N_A_129_279#_c_54_n 0.0152133f $X=3.12 $Y=4.07 $X2=0.895
+ $Y2=2.105
cc_25 N_VPB_M1001_b N_A_129_279#_M1003_g 0.0571164f $X=-0.33 $Y=1.885 $X2=1.675
+ $Y2=2.965
cc_26 VPB N_A_129_279#_M1003_g 0.00970178f $X=0 $Y=3.955 $X2=1.675 $Y2=2.965
cc_27 N_VPB_c_24_p N_A_129_279#_M1003_g 0.0152133f $X=3.12 $Y=4.07 $X2=1.675
+ $Y2=2.965
cc_28 N_VPB_M1001_b N_A_129_279#_c_50_n 0.0527693f $X=-0.33 $Y=1.885 $X2=3.065
+ $Y2=2.34
cc_29 N_VPB_M1001_b N_A_129_279#_c_53_n 0.0324531f $X=-0.33 $Y=1.885 $X2=1.695
+ $Y2=1.75
cc_30 N_VPB_M1001_b A 0.00767318f $X=-0.33 $Y=1.885 $X2=0.895 $Y2=2.965
cc_31 N_VPB_M1001_b N_A_c_102_n 0.0229742f $X=-0.33 $Y=1.885 $X2=0.915 $Y2=0.91
cc_32 N_VPB_M1001_b N_A_c_106_n 0.0422619f $X=-0.33 $Y=1.885 $X2=1.675 $Y2=2.965
cc_33 N_VPB_M1001_b N_VPWR_c_125_n 0.0825346f $X=-0.33 $Y=1.885 $X2=0.915
+ $Y2=1.395
cc_34 VPB N_VPWR_c_125_n 0.00349285f $X=0 $Y=3.955 $X2=0.915 $Y2=1.395
cc_35 N_VPB_c_24_p N_VPWR_c_125_n 0.0475576f $X=3.12 $Y=4.07 $X2=0.915 $Y2=1.395
cc_36 N_VPB_M1001_b N_VPWR_c_128_n 0.0331845f $X=-0.33 $Y=1.885 $X2=2.98
+ $Y2=1.51
cc_37 VPB N_VPWR_c_128_n 0.00447364f $X=0 $Y=3.955 $X2=2.98 $Y2=1.51
cc_38 N_VPB_c_24_p N_VPWR_c_128_n 0.0644672f $X=3.12 $Y=4.07 $X2=2.98 $Y2=1.51
cc_39 N_VPB_M1001_b N_VPWR_c_131_n 0.0574803f $X=-0.33 $Y=1.885 $X2=3.085
+ $Y2=1.075
cc_40 VPB N_VPWR_c_131_n 0.357521f $X=0 $Y=3.955 $X2=3.085 $Y2=1.075
cc_41 N_VPB_c_24_p N_VPWR_c_131_n 0.0158542f $X=3.12 $Y=4.07 $X2=3.085 $Y2=1.075
cc_42 N_VPB_M1001_b N_X_c_152_n 0.00790968f $X=-0.33 $Y=1.885 $X2=0.895
+ $Y2=2.965
cc_43 VPB N_X_c_152_n 5.14916e-19 $X=0 $Y=3.955 $X2=0.895 $Y2=2.965
cc_44 N_VPB_c_24_p N_X_c_152_n 0.00887752f $X=3.12 $Y=4.07 $X2=0.895 $Y2=2.965
cc_45 N_A_129_279#_M1003_g A 0.00422806f $X=1.675 $Y=2.965 $X2=0 $Y2=0
cc_46 N_A_129_279#_c_49_n A 0.0530016f $X=2.98 $Y=1.51 $X2=0 $Y2=0
cc_47 N_A_129_279#_c_50_n A 0.024569f $X=3.065 $Y=2.34 $X2=0 $Y2=0
cc_48 N_A_129_279#_c_53_n A 0.00244686f $X=1.695 $Y=1.75 $X2=0 $Y2=0
cc_49 N_A_129_279#_M1003_g N_A_c_102_n 0.0170835f $X=1.675 $Y=2.965 $X2=0 $Y2=0
cc_50 N_A_129_279#_c_49_n N_A_c_102_n 0.0379174f $X=2.98 $Y=1.51 $X2=0 $Y2=0
cc_51 N_A_129_279#_c_50_n N_A_c_102_n 0.0185373f $X=3.065 $Y=2.34 $X2=0 $Y2=0
cc_52 N_A_129_279#_c_69_p N_A_c_102_n 9.89615e-19 $X=1.717 $Y=1.51 $X2=0 $Y2=0
cc_53 N_A_129_279#_c_53_n N_A_c_102_n 0.0131328f $X=1.695 $Y=1.75 $X2=0 $Y2=0
cc_54 N_A_129_279#_c_47_n N_A_c_103_n 0.0106668f $X=1.695 $Y=1.395 $X2=0 $Y2=0
cc_55 N_A_129_279#_c_51_n N_A_c_103_n 0.00836499f $X=3.085 $Y=1.075 $X2=0 $Y2=0
cc_56 N_A_129_279#_c_50_n N_A_c_106_n 0.00878462f $X=3.065 $Y=2.34 $X2=0 $Y2=0
cc_57 N_A_129_279#_c_54_n N_VPWR_c_125_n 0.0813488f $X=0.895 $Y=2.105 $X2=0.24
+ $Y2=0
cc_58 N_A_129_279#_M1003_g N_VPWR_c_128_n 0.0775691f $X=1.675 $Y=2.965 $X2=0
+ $Y2=0
cc_59 N_A_129_279#_c_50_n N_VPWR_c_128_n 0.0297448f $X=3.065 $Y=2.34 $X2=0 $Y2=0
cc_60 N_A_129_279#_c_69_p N_VPWR_c_128_n 0.00898391f $X=1.717 $Y=1.51 $X2=0
+ $Y2=0
cc_61 N_A_129_279#_c_54_n N_VPWR_c_131_n 0.00829406f $X=0.895 $Y=2.105 $X2=0
+ $Y2=0
cc_62 N_A_129_279#_M1003_g N_VPWR_c_131_n 0.00841417f $X=1.675 $Y=2.965 $X2=0
+ $Y2=0
cc_63 N_A_129_279#_c_50_n N_VPWR_c_131_n 0.011836f $X=3.065 $Y=2.34 $X2=0 $Y2=0
cc_64 N_A_129_279#_c_54_n N_X_c_152_n 0.00313915f $X=0.895 $Y=2.105 $X2=0 $Y2=0
cc_65 N_A_129_279#_M1003_g N_X_c_152_n 0.0065902f $X=1.675 $Y=2.965 $X2=0 $Y2=0
cc_66 N_A_129_279#_c_53_n N_X_c_152_n 0.0169982f $X=1.695 $Y=1.75 $X2=0 $Y2=0
cc_67 N_A_129_279#_c_45_n N_X_c_149_n 0.00308135f $X=0.915 $Y=1.395 $X2=0 $Y2=0
cc_68 N_A_129_279#_c_47_n N_X_c_149_n 0.00373379f $X=1.695 $Y=1.395 $X2=0 $Y2=0
cc_69 N_A_129_279#_c_69_p N_X_c_149_n 0.008418f $X=1.717 $Y=1.51 $X2=0 $Y2=0
cc_70 N_A_129_279#_c_53_n N_X_c_149_n 0.0144434f $X=1.695 $Y=1.75 $X2=0 $Y2=0
cc_71 N_A_129_279#_c_69_p X 0.015286f $X=1.717 $Y=1.51 $X2=0 $Y2=0
cc_72 N_A_129_279#_c_53_n X 0.0573539f $X=1.695 $Y=1.75 $X2=0 $Y2=0
cc_73 N_A_129_279#_c_45_n N_VGND_c_175_n 0.0579063f $X=0.915 $Y=1.395 $X2=0.24
+ $Y2=0
cc_74 N_A_129_279#_c_47_n N_VGND_c_175_n 6.27588e-19 $X=1.695 $Y=1.395 $X2=0.24
+ $Y2=0
cc_75 N_A_129_279#_c_53_n N_VGND_c_175_n 6.36121e-19 $X=1.695 $Y=1.75 $X2=0.24
+ $Y2=0
cc_76 N_A_129_279#_c_45_n N_VGND_c_177_n 6.0418e-19 $X=0.915 $Y=1.395 $X2=0
+ $Y2=0
cc_77 N_A_129_279#_c_47_n N_VGND_c_177_n 0.0524473f $X=1.695 $Y=1.395 $X2=0
+ $Y2=0
cc_78 N_A_129_279#_c_49_n N_VGND_c_177_n 0.0676614f $X=2.98 $Y=1.51 $X2=0 $Y2=0
cc_79 N_A_129_279#_c_51_n N_VGND_c_177_n 0.0183139f $X=3.085 $Y=1.075 $X2=0
+ $Y2=0
cc_80 N_A_129_279#_c_69_p N_VGND_c_177_n 0.022445f $X=1.717 $Y=1.51 $X2=0 $Y2=0
cc_81 N_A_129_279#_c_45_n N_VGND_c_179_n 0.00774885f $X=0.915 $Y=1.395 $X2=1.68
+ $Y2=0.057
cc_82 N_A_129_279#_c_47_n N_VGND_c_179_n 0.00774885f $X=1.695 $Y=1.395 $X2=1.68
+ $Y2=0.057
cc_83 N_A_129_279#_c_51_n N_VGND_c_179_n 0.0137969f $X=3.085 $Y=1.075 $X2=1.68
+ $Y2=0.057
cc_84 A N_VPWR_c_128_n 0.056015f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_85 N_A_c_106_n N_VPWR_c_128_n 0.0677433f $X=2.685 $Y=2.105 $X2=0 $Y2=0
cc_86 N_A_c_106_n N_VPWR_c_131_n 0.00357298f $X=2.685 $Y=2.105 $X2=0 $Y2=0
cc_87 A N_X_c_152_n 0.010268f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_88 N_A_c_103_n N_VGND_c_177_n 0.0482894f $X=2.685 $Y=1.395 $X2=0 $Y2=0
cc_89 N_A_c_103_n N_VGND_c_179_n 0.00411567f $X=2.685 $Y=1.395 $X2=1.68
+ $Y2=0.057
cc_90 N_VPWR_c_131_n N_X_M1001_d 0.00442064f $X=2.715 $Y=3.59 $X2=0 $Y2=0
cc_91 N_VPWR_c_125_n N_X_c_152_n 0.0676307f $X=0.505 $Y=2.34 $X2=0.24 $Y2=4.07
cc_92 N_VPWR_c_128_n N_X_c_152_n 0.0612155f $X=2.065 $Y=2.385 $X2=0.24 $Y2=4.07
cc_93 N_VPWR_c_131_n N_X_c_152_n 0.0229352f $X=2.715 $Y=3.59 $X2=0.24 $Y2=4.07
cc_94 N_VPWR_c_125_n X 0.0397037f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_95 N_X_c_149_n N_VGND_c_175_n 0.0362614f $X=1.305 $Y=0.66 $X2=0.24 $Y2=0
cc_96 X N_VGND_c_175_n 0.0613864f $X=1.115 $Y=1.58 $X2=0.24 $Y2=0
cc_97 N_X_c_149_n N_VGND_c_177_n 0.0316484f $X=1.305 $Y=0.66 $X2=0 $Y2=0
cc_98 N_X_M1002_d N_VGND_c_179_n 0.00442064f $X=1.165 $Y=0.535 $X2=1.68
+ $Y2=0.057
cc_99 N_X_c_149_n N_VGND_c_179_n 0.0174197f $X=1.305 $Y=0.66 $X2=1.68 $Y2=0.057
