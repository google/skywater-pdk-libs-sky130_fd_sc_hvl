* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1 A LVPWR VGND VNB VPB VPWR X
M1000 a_1197_107# a_772_151# a_686_151# VNB nhv w=1.5e+06u l=500000u
+  ad=1.215e+12p pd=1.062e+07u as=7.95e+11p ps=7.06e+06u
M1001 VGND a_573_897# a_816_1221# VNB nhv w=1.5e+06u l=500000u
+  ad=1.03875e+12p pd=9.21e+06u as=4.2e+11p ps=3.56e+06u
M1002 a_1400_777# a_816_1221# a_1606_563# VPB phv w=420000u l=1e+06u
+  ad=2.457e+11p pd=2.14e+06u as=4.599e+11p ps=4.13e+06u
M1003 a_1606_563# a_1406_429# a_1400_777# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_816_1221# a_573_897# VGND VNB nhv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1005 LVPWR A a_573_897# LVPWR phighvt w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=2.478e+11p ps=2.27e+06u
M1006 a_1606_563# a_1406_429# a_816_1221# VPB phv w=420000u l=1e+06u
+  ad=0p pd=0u as=1.0092e+12p ps=9.05e+06u
M1007 X a_1406_429# VGND VNB nhv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u
M1008 VPWR a_1400_777# a_816_1221# VPB phv w=1.5e+06u l=500000u
+  ad=9.75e+11p pd=7.3e+06u as=0p ps=0u
M1009 a_816_1221# a_1400_777# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1197_107# a_1406_429# a_1400_777# VNB nhv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=4.2e+11p ps=3.56e+06u
M1011 VGND a_816_1221# a_1406_429# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u
M1012 a_686_151# a_772_151# a_1197_107# VNB nhv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_816_1221# a_1406_429# VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=3.975e+11p ps=3.53e+06u
M1014 X a_1406_429# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=3.975e+11p pd=3.53e+06u as=0p ps=0u
M1015 a_686_151# A a_573_897# VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=2.478e+11p ps=2.27e+06u
M1016 a_772_151# a_573_897# a_686_151# VNB nshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1017 a_772_151# a_573_897# LVPWR LVPWR phighvt w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1018 a_1400_777# a_1406_429# a_1197_107# VNB nhv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
