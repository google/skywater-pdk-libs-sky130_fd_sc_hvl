* File: sky130_fd_sc_hvl__buf_16.pxi.spice
* Created: Fri Aug 28 09:32:50 2020
* 
x_PM_SKY130_FD_SC_HVL__BUF_16%VNB N_VNB_M1006_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__BUF_16%VNB
x_PM_SKY130_FD_SC_HVL__BUF_16%VPB N_VPB_M1000_b VPB N_VPB_c_91_p N_VPB_c_92_p
+ VPB PM_SKY130_FD_SC_HVL__BUF_16%VPB
x_PM_SKY130_FD_SC_HVL__BUF_16%A N_A_c_227_n N_A_M1006_g N_A_M1000_g N_A_c_229_n
+ N_A_M1016_g N_A_M1005_g N_A_c_231_n N_A_M1019_g N_A_M1011_g N_A_c_233_n
+ N_A_M1026_g N_A_M1023_g N_A_c_235_n N_A_M1040_g N_A_M1029_g N_A_c_237_n
+ N_A_M1043_g N_A_M1036_g A A A A A A A N_A_c_239_n N_A_c_240_n
+ PM_SKY130_FD_SC_HVL__BUF_16%A
x_PM_SKY130_FD_SC_HVL__BUF_16%A_183_141# N_A_183_141#_M1006_s
+ N_A_183_141#_M1019_s N_A_183_141#_M1040_s N_A_183_141#_M1000_s
+ N_A_183_141#_M1011_s N_A_183_141#_M1029_s N_A_183_141#_c_359_n
+ N_A_183_141#_M1002_g N_A_183_141#_M1001_g N_A_183_141#_c_361_n
+ N_A_183_141#_M1004_g N_A_183_141#_M1003_g N_A_183_141#_c_363_n
+ N_A_183_141#_M1007_g N_A_183_141#_M1008_g N_A_183_141#_c_365_n
+ N_A_183_141#_M1009_g N_A_183_141#_M1010_g N_A_183_141#_c_367_n
+ N_A_183_141#_M1014_g N_A_183_141#_M1012_g N_A_183_141#_c_369_n
+ N_A_183_141#_M1017_g N_A_183_141#_M1013_g N_A_183_141#_c_371_n
+ N_A_183_141#_M1020_g N_A_183_141#_M1015_g N_A_183_141#_c_373_n
+ N_A_183_141#_M1024_g N_A_183_141#_M1018_g N_A_183_141#_c_375_n
+ N_A_183_141#_M1027_g N_A_183_141#_M1021_g N_A_183_141#_c_377_n
+ N_A_183_141#_M1028_g N_A_183_141#_M1022_g N_A_183_141#_c_379_n
+ N_A_183_141#_M1030_g N_A_183_141#_M1025_g N_A_183_141#_c_381_n
+ N_A_183_141#_M1032_g N_A_183_141#_M1031_g N_A_183_141#_c_383_n
+ N_A_183_141#_M1034_g N_A_183_141#_M1033_g N_A_183_141#_c_385_n
+ N_A_183_141#_M1035_g N_A_183_141#_M1038_g N_A_183_141#_c_387_n
+ N_A_183_141#_M1037_g N_A_183_141#_M1039_g N_A_183_141#_c_389_n
+ N_A_183_141#_M1041_g N_A_183_141#_M1042_g N_A_183_141#_c_391_n
+ N_A_183_141#_c_457_n N_A_183_141#_c_472_n N_A_183_141#_c_476_n
+ N_A_183_141#_c_479_n N_A_183_141#_c_483_n N_A_183_141#_c_392_n
+ N_A_183_141#_c_460_n N_A_183_141#_c_490_n N_A_183_141#_c_494_n
+ N_A_183_141#_c_463_n N_A_183_141#_c_393_n N_A_183_141#_c_502_n
+ N_A_183_141#_c_504_n N_A_183_141#_c_507_n N_A_183_141#_c_511_n
+ N_A_183_141#_c_514_n N_A_183_141#_c_517_n N_A_183_141#_c_546_p
+ N_A_183_141#_c_636_p N_A_183_141#_c_394_n N_A_183_141#_c_547_p
+ N_A_183_141#_c_395_n N_A_183_141#_c_549_p N_A_183_141#_c_647_p
+ N_A_183_141#_c_396_n N_A_183_141#_c_556_p N_A_183_141#_c_397_n
+ N_A_183_141#_c_558_p N_A_183_141#_c_657_p N_A_183_141#_c_398_n
+ N_A_183_141#_c_565_p N_A_183_141#_c_399_n N_A_183_141#_c_567_p
+ N_A_183_141#_c_667_p N_A_183_141#_c_400_n N_A_183_141#_c_574_p
+ N_A_183_141#_c_401_n N_A_183_141#_c_576_p N_A_183_141#_c_677_p
+ N_A_183_141#_c_402_n N_A_183_141#_c_583_p N_A_183_141#_c_403_n
+ N_A_183_141#_c_585_p N_A_183_141#_c_687_p N_A_183_141#_c_404_n
+ N_A_183_141#_c_592_p N_A_183_141#_c_405_n N_A_183_141#_c_594_p
+ N_A_183_141#_c_697_p N_A_183_141#_c_601_p N_A_183_141#_c_406_n
+ N_A_183_141#_c_407_n N_A_183_141#_c_520_n N_A_183_141#_c_523_n
+ PM_SKY130_FD_SC_HVL__BUF_16%A_183_141#
x_PM_SKY130_FD_SC_HVL__BUF_16%VPWR N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_M1023_d
+ N_VPWR_M1036_d N_VPWR_M1003_s N_VPWR_M1010_s N_VPWR_M1013_s N_VPWR_M1018_s
+ N_VPWR_M1022_s N_VPWR_M1031_s N_VPWR_M1038_s N_VPWR_M1042_s VPWR
+ N_VPWR_c_841_n N_VPWR_c_844_n N_VPWR_c_846_n N_VPWR_c_848_n N_VPWR_c_850_n
+ N_VPWR_c_853_n N_VPWR_c_856_n N_VPWR_c_859_n N_VPWR_c_862_n N_VPWR_c_865_n
+ N_VPWR_c_868_n N_VPWR_c_871_n N_VPWR_c_874_n PM_SKY130_FD_SC_HVL__BUF_16%VPWR
x_PM_SKY130_FD_SC_HVL__BUF_16%X N_X_M1002_s N_X_M1007_s N_X_M1014_s N_X_M1020_s
+ N_X_M1027_s N_X_M1030_s N_X_M1034_s N_X_M1037_s N_X_M1001_d N_X_M1008_d
+ N_X_M1012_d N_X_M1015_d N_X_M1021_d N_X_M1025_d N_X_M1033_d N_X_M1039_d X
+ N_X_c_1046_n N_X_c_1049_n N_X_c_1052_n N_X_c_1055_n N_X_c_1058_n N_X_c_1061_n
+ N_X_c_1064_n N_X_c_1067_n N_X_c_1148_n N_X_c_1152_n N_X_c_1153_n N_X_c_1157_n
+ N_X_c_1158_n N_X_c_1162_n N_X_c_1163_n N_X_c_1167_n X N_X_c_1168_n
+ N_X_c_1172_n N_X_c_1173_n N_X_c_1177_n N_X_c_1178_n N_X_c_1182_n
+ PM_SKY130_FD_SC_HVL__BUF_16%X
x_PM_SKY130_FD_SC_HVL__BUF_16%VGND N_VGND_M1006_d N_VGND_M1016_d N_VGND_M1026_d
+ N_VGND_M1043_d N_VGND_M1004_d N_VGND_M1009_d N_VGND_M1017_d N_VGND_M1024_d
+ N_VGND_M1028_d N_VGND_M1032_d N_VGND_M1035_d N_VGND_M1041_d VGND
+ N_VGND_c_1254_n N_VGND_c_1256_n N_VGND_c_1258_n N_VGND_c_1260_n
+ N_VGND_c_1262_n N_VGND_c_1264_n N_VGND_c_1266_n N_VGND_c_1268_n
+ N_VGND_c_1270_n N_VGND_c_1272_n N_VGND_c_1274_n N_VGND_c_1276_n
+ N_VGND_c_1278_n PM_SKY130_FD_SC_HVL__BUF_16%VGND
cc_1 N_VNB_M1006_b N_A_c_227_n 0.0468242f $X=-0.33 $Y=-0.265 $X2=0.665 $Y2=1.565
cc_2 N_VNB_c_2_p N_A_c_227_n 0.00104452f $X=17.52 $Y=0 $X2=0.665 $Y2=1.565
cc_3 N_VNB_M1006_b N_A_c_229_n 0.0390915f $X=-0.33 $Y=-0.265 $X2=1.445 $Y2=1.565
cc_4 N_VNB_c_2_p N_A_c_229_n 5.62728e-19 $X=17.52 $Y=0 $X2=1.445 $Y2=1.565
cc_5 N_VNB_M1006_b N_A_c_231_n 0.0405965f $X=-0.33 $Y=-0.265 $X2=2.225 $Y2=1.565
cc_6 N_VNB_c_2_p N_A_c_231_n 9.48159e-19 $X=17.52 $Y=0 $X2=2.225 $Y2=1.565
cc_7 N_VNB_M1006_b N_A_c_233_n 0.0400608f $X=-0.33 $Y=-0.265 $X2=3.005 $Y2=1.565
cc_8 N_VNB_c_2_p N_A_c_233_n 7.93986e-19 $X=17.52 $Y=0 $X2=3.005 $Y2=1.565
cc_9 N_VNB_M1006_b N_A_c_235_n 0.0397162f $X=-0.33 $Y=-0.265 $X2=3.785 $Y2=1.565
cc_10 N_VNB_c_2_p N_A_c_235_n 6.97629e-19 $X=17.52 $Y=0 $X2=3.785 $Y2=1.565
cc_11 N_VNB_M1006_b N_A_c_237_n 0.0382604f $X=-0.33 $Y=-0.265 $X2=4.565
+ $Y2=1.565
cc_12 N_VNB_c_2_p N_A_c_237_n 4.85642e-19 $X=17.52 $Y=0 $X2=4.565 $Y2=1.565
cc_13 N_VNB_M1006_b N_A_c_239_n 0.0094895f $X=-0.33 $Y=-0.265 $X2=4.465 $Y2=1.73
cc_14 N_VNB_M1006_b N_A_c_240_n 0.18914f $X=-0.33 $Y=-0.265 $X2=4.565 $Y2=1.815
cc_15 N_VNB_M1006_b N_A_183_141#_c_359_n 0.0404132f $X=-0.33 $Y=-0.265 $X2=2.225
+ $Y2=2.965
cc_16 N_VNB_c_2_p N_A_183_141#_c_359_n 0.00102524f $X=17.52 $Y=0 $X2=2.225
+ $Y2=2.965
cc_17 N_VNB_M1006_b N_A_183_141#_c_361_n 0.0395228f $X=-0.33 $Y=-0.265 $X2=3.005
+ $Y2=2.965
cc_18 N_VNB_c_2_p N_A_183_141#_c_361_n 7.55443e-19 $X=17.52 $Y=0 $X2=3.005
+ $Y2=2.965
cc_19 N_VNB_M1006_b N_A_183_141#_c_363_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=3.785
+ $Y2=2.965
cc_20 N_VNB_c_2_p N_A_183_141#_c_363_n 7.55443e-19 $X=17.52 $Y=0 $X2=3.785
+ $Y2=2.965
cc_21 N_VNB_M1006_b N_A_183_141#_c_365_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=4.565
+ $Y2=2.965
cc_22 N_VNB_c_2_p N_A_183_141#_c_365_n 7.55443e-19 $X=17.52 $Y=0 $X2=4.565
+ $Y2=2.965
cc_23 N_VNB_M1006_b N_A_183_141#_c_367_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=2.555
+ $Y2=1.58
cc_24 N_VNB_c_2_p N_A_183_141#_c_367_n 7.55443e-19 $X=17.52 $Y=0 $X2=2.555
+ $Y2=1.58
cc_25 N_VNB_M1006_b N_A_183_141#_c_369_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_26 N_VNB_c_2_p N_A_183_141#_c_369_n 7.55443e-19 $X=17.52 $Y=0 $X2=0 $Y2=0
cc_27 N_VNB_M1006_b N_A_183_141#_c_371_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0.665
+ $Y2=1.815
cc_28 N_VNB_c_2_p N_A_183_141#_c_371_n 7.55443e-19 $X=17.52 $Y=0 $X2=0.665
+ $Y2=1.815
cc_29 N_VNB_M1006_b N_A_183_141#_c_373_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=4.465
+ $Y2=1.73
cc_30 N_VNB_c_2_p N_A_183_141#_c_373_n 7.55443e-19 $X=17.52 $Y=0 $X2=4.465
+ $Y2=1.73
cc_31 N_VNB_M1006_b N_A_183_141#_c_375_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=1.2
+ $Y2=1.697
cc_32 N_VNB_c_2_p N_A_183_141#_c_375_n 7.55443e-19 $X=17.52 $Y=0 $X2=1.2
+ $Y2=1.697
cc_33 N_VNB_M1006_b N_A_183_141#_c_377_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_34 N_VNB_c_2_p N_A_183_141#_c_377_n 7.55443e-19 $X=17.52 $Y=0 $X2=0 $Y2=0
cc_35 N_VNB_M1006_b N_A_183_141#_c_379_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_36 N_VNB_c_2_p N_A_183_141#_c_379_n 7.55443e-19 $X=17.52 $Y=0 $X2=0 $Y2=0
cc_37 N_VNB_M1006_b N_A_183_141#_c_381_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_38 N_VNB_c_2_p N_A_183_141#_c_381_n 7.55443e-19 $X=17.52 $Y=0 $X2=0 $Y2=0
cc_39 N_VNB_M1006_b N_A_183_141#_c_383_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_40 N_VNB_c_2_p N_A_183_141#_c_383_n 7.55443e-19 $X=17.52 $Y=0 $X2=0 $Y2=0
cc_41 N_VNB_M1006_b N_A_183_141#_c_385_n 0.0395213f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_42 N_VNB_c_2_p N_A_183_141#_c_385_n 7.55443e-19 $X=17.52 $Y=0 $X2=0 $Y2=0
cc_43 N_VNB_M1006_b N_A_183_141#_c_387_n 0.0395229f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_44 N_VNB_c_2_p N_A_183_141#_c_387_n 7.55443e-19 $X=17.52 $Y=0 $X2=0 $Y2=0
cc_45 N_VNB_M1006_b N_A_183_141#_c_389_n 0.525041f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_46 N_VNB_c_2_p N_A_183_141#_c_389_n 0.00106379f $X=17.52 $Y=0 $X2=0 $Y2=0
cc_47 N_VNB_M1006_b N_A_183_141#_c_391_n 0.00340102f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_48 N_VNB_M1006_b N_A_183_141#_c_392_n 0.00388959f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_49 N_VNB_M1006_b N_A_183_141#_c_393_n 0.00250789f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_50 N_VNB_M1006_b N_A_183_141#_c_394_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_51 N_VNB_M1006_b N_A_183_141#_c_395_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_52 N_VNB_M1006_b N_A_183_141#_c_396_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_53 N_VNB_M1006_b N_A_183_141#_c_397_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_54 N_VNB_M1006_b N_A_183_141#_c_398_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_55 N_VNB_M1006_b N_A_183_141#_c_399_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_56 N_VNB_M1006_b N_A_183_141#_c_400_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_57 N_VNB_M1006_b N_A_183_141#_c_401_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_58 N_VNB_M1006_b N_A_183_141#_c_402_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_59 N_VNB_M1006_b N_A_183_141#_c_403_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_60 N_VNB_M1006_b N_A_183_141#_c_404_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_61 N_VNB_M1006_b N_A_183_141#_c_405_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_62 N_VNB_M1006_b N_A_183_141#_c_406_n 0.00198224f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_63 N_VNB_M1006_b N_A_183_141#_c_407_n 3.38774e-19 $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_64 N_VNB_M1006_b N_VGND_c_1254_n 0.0613833f $X=-0.33 $Y=-0.265 $X2=4.565
+ $Y2=2.965
cc_65 N_VNB_c_2_p N_VGND_c_1254_n 0.00138265f $X=17.52 $Y=0 $X2=4.565 $Y2=2.965
cc_66 N_VNB_M1006_b N_VGND_c_1256_n 0.0415829f $X=-0.33 $Y=-0.265 $X2=2.555
+ $Y2=1.58
cc_67 N_VNB_c_2_p N_VGND_c_1256_n 0.00234213f $X=17.52 $Y=0 $X2=2.555 $Y2=1.58
cc_68 N_VNB_M1006_b N_VGND_c_1258_n 0.0399392f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_69 N_VNB_c_2_p N_VGND_c_1258_n 0.0023214f $X=17.52 $Y=0 $X2=0 $Y2=0
cc_70 N_VNB_M1006_b N_VGND_c_1260_n 0.0397337f $X=-0.33 $Y=-0.265 $X2=3.785
+ $Y2=1.815
cc_71 N_VNB_c_2_p N_VGND_c_1260_n 0.00230841f $X=17.52 $Y=0 $X2=3.785 $Y2=1.815
cc_72 N_VNB_M1006_b N_VGND_c_1262_n 0.039901f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_73 N_VNB_c_2_p N_VGND_c_1262_n 0.00230355f $X=17.52 $Y=0 $X2=0 $Y2=0
cc_74 N_VNB_M1006_b N_VGND_c_1264_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=3.12
+ $Y2=1.697
cc_75 N_VNB_c_2_p N_VGND_c_1264_n 0.00230355f $X=17.52 $Y=0 $X2=3.12 $Y2=1.697
cc_76 N_VNB_M1006_b N_VGND_c_1266_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_77 N_VNB_c_2_p N_VGND_c_1266_n 0.00230355f $X=17.52 $Y=0 $X2=0 $Y2=0
cc_78 N_VNB_M1006_b N_VGND_c_1268_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_79 N_VNB_c_2_p N_VGND_c_1268_n 0.00230355f $X=17.52 $Y=0 $X2=0 $Y2=0
cc_80 N_VNB_M1006_b N_VGND_c_1270_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_81 N_VNB_c_2_p N_VGND_c_1270_n 0.00230355f $X=17.52 $Y=0 $X2=0 $Y2=0
cc_82 N_VNB_M1006_b N_VGND_c_1272_n 0.0393532f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_83 N_VNB_c_2_p N_VGND_c_1272_n 0.00230355f $X=17.52 $Y=0 $X2=0 $Y2=0
cc_84 N_VNB_M1006_b N_VGND_c_1274_n 0.039901f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_85 N_VNB_c_2_p N_VGND_c_1274_n 0.00230355f $X=17.52 $Y=0 $X2=0 $Y2=0
cc_86 N_VNB_M1006_b N_VGND_c_1276_n 0.0684821f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_87 N_VNB_c_2_p N_VGND_c_1276_n 0.00136968f $X=17.52 $Y=0 $X2=0 $Y2=0
cc_88 N_VNB_M1006_b N_VGND_c_1278_n 0.263558f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_89 N_VNB_c_2_p N_VGND_c_1278_n 1.9002f $X=17.52 $Y=0 $X2=0 $Y2=0
cc_90 N_VPB_M1000_b N_A_M1000_g 0.0430944f $X=-0.33 $Y=1.885 $X2=0.665 $Y2=2.965
cc_91 N_VPB_c_91_p N_A_M1000_g 0.0157621f $X=17.52 $Y=4.07 $X2=0.665 $Y2=2.965
cc_92 N_VPB_c_92_p N_A_M1000_g 0.00970178f $X=17.52 $Y=4.07 $X2=0.665 $Y2=2.965
cc_93 N_VPB_M1000_b N_A_M1005_g 0.0352958f $X=-0.33 $Y=1.885 $X2=1.445 $Y2=2.965
cc_94 N_VPB_c_91_p N_A_M1005_g 0.0157169f $X=17.52 $Y=4.07 $X2=1.445 $Y2=2.965
cc_95 N_VPB_c_92_p N_A_M1005_g 0.00970178f $X=17.52 $Y=4.07 $X2=1.445 $Y2=2.965
cc_96 N_VPB_M1000_b N_A_M1011_g 0.0352691f $X=-0.33 $Y=1.885 $X2=2.225 $Y2=2.965
cc_97 N_VPB_c_91_p N_A_M1011_g 0.0159522f $X=17.52 $Y=4.07 $X2=2.225 $Y2=2.965
cc_98 N_VPB_c_92_p N_A_M1011_g 0.00970178f $X=17.52 $Y=4.07 $X2=2.225 $Y2=2.965
cc_99 N_VPB_M1000_b N_A_M1023_g 0.0352958f $X=-0.33 $Y=1.885 $X2=3.005 $Y2=2.965
cc_100 N_VPB_c_91_p N_A_M1023_g 0.0154933f $X=17.52 $Y=4.07 $X2=3.005 $Y2=2.965
cc_101 N_VPB_c_92_p N_A_M1023_g 0.00970178f $X=17.52 $Y=4.07 $X2=3.005 $Y2=2.965
cc_102 N_VPB_M1000_b N_A_M1029_g 0.0352669f $X=-0.33 $Y=1.885 $X2=3.785
+ $Y2=2.965
cc_103 N_VPB_c_91_p N_A_M1029_g 0.0159373f $X=17.52 $Y=4.07 $X2=3.785 $Y2=2.965
cc_104 N_VPB_c_92_p N_A_M1029_g 0.00970178f $X=17.52 $Y=4.07 $X2=3.785 $Y2=2.965
cc_105 N_VPB_M1000_b N_A_M1036_g 0.0354096f $X=-0.33 $Y=1.885 $X2=4.565
+ $Y2=2.965
cc_106 N_VPB_c_91_p N_A_M1036_g 0.0157169f $X=17.52 $Y=4.07 $X2=4.565 $Y2=2.965
cc_107 N_VPB_c_92_p N_A_M1036_g 0.00970178f $X=17.52 $Y=4.07 $X2=4.565 $Y2=2.965
cc_108 N_VPB_M1000_b N_A_c_240_n 0.119162f $X=-0.33 $Y=1.885 $X2=4.565 $Y2=1.815
cc_109 N_VPB_M1000_b N_A_183_141#_M1001_g 0.0401913f $X=-0.33 $Y=1.885 $X2=3.005
+ $Y2=1.08
cc_110 N_VPB_c_91_p N_A_183_141#_M1001_g 0.0165487f $X=17.52 $Y=4.07 $X2=3.005
+ $Y2=1.08
cc_111 N_VPB_c_92_p N_A_183_141#_M1001_g 0.00970178f $X=17.52 $Y=4.07 $X2=3.005
+ $Y2=1.08
cc_112 N_VPB_M1000_b N_A_183_141#_M1003_g 0.040726f $X=-0.33 $Y=1.885 $X2=3.785
+ $Y2=1.08
cc_113 N_VPB_c_91_p N_A_183_141#_M1003_g 0.0157621f $X=17.52 $Y=4.07 $X2=3.785
+ $Y2=1.08
cc_114 N_VPB_c_92_p N_A_183_141#_M1003_g 0.00970178f $X=17.52 $Y=4.07 $X2=3.785
+ $Y2=1.08
cc_115 N_VPB_M1000_b N_A_183_141#_M1008_g 0.040726f $X=-0.33 $Y=1.885 $X2=4.565
+ $Y2=1.08
cc_116 N_VPB_c_91_p N_A_183_141#_M1008_g 0.0157621f $X=17.52 $Y=4.07 $X2=4.565
+ $Y2=1.08
cc_117 N_VPB_c_92_p N_A_183_141#_M1008_g 0.00970178f $X=17.52 $Y=4.07 $X2=4.565
+ $Y2=1.08
cc_118 N_VPB_M1000_b N_A_183_141#_M1010_g 0.040726f $X=-0.33 $Y=1.885 $X2=1.595
+ $Y2=1.58
cc_119 N_VPB_c_91_p N_A_183_141#_M1010_g 0.0157621f $X=17.52 $Y=4.07 $X2=1.595
+ $Y2=1.58
cc_120 N_VPB_c_92_p N_A_183_141#_M1010_g 0.00970178f $X=17.52 $Y=4.07 $X2=1.595
+ $Y2=1.58
cc_121 N_VPB_M1000_b N_A_183_141#_M1012_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_122 N_VPB_c_91_p N_A_183_141#_M1012_g 0.0157621f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_123 N_VPB_c_92_p N_A_183_141#_M1012_g 0.00970178f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_124 N_VPB_M1000_b N_A_183_141#_M1013_g 0.040726f $X=-0.33 $Y=1.885 $X2=0.385
+ $Y2=1.73
cc_125 N_VPB_c_91_p N_A_183_141#_M1013_g 0.0157621f $X=17.52 $Y=4.07 $X2=0.385
+ $Y2=1.73
cc_126 N_VPB_c_92_p N_A_183_141#_M1013_g 0.00970178f $X=17.52 $Y=4.07 $X2=0.385
+ $Y2=1.73
cc_127 N_VPB_M1000_b N_A_183_141#_M1015_g 0.040726f $X=-0.33 $Y=1.885 $X2=4.465
+ $Y2=1.815
cc_128 N_VPB_c_91_p N_A_183_141#_M1015_g 0.0157621f $X=17.52 $Y=4.07 $X2=4.465
+ $Y2=1.815
cc_129 N_VPB_c_92_p N_A_183_141#_M1015_g 0.00970178f $X=17.52 $Y=4.07 $X2=4.465
+ $Y2=1.815
cc_130 N_VPB_M1000_b N_A_183_141#_M1018_g 0.040726f $X=-0.33 $Y=1.885 $X2=0.72
+ $Y2=1.697
cc_131 N_VPB_c_91_p N_A_183_141#_M1018_g 0.0157621f $X=17.52 $Y=4.07 $X2=0.72
+ $Y2=1.697
cc_132 N_VPB_c_92_p N_A_183_141#_M1018_g 0.00970178f $X=17.52 $Y=4.07 $X2=0.72
+ $Y2=1.697
cc_133 N_VPB_M1000_b N_A_183_141#_M1021_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_134 N_VPB_c_91_p N_A_183_141#_M1021_g 0.0157621f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_135 N_VPB_c_92_p N_A_183_141#_M1021_g 0.00970178f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_136 N_VPB_M1000_b N_A_183_141#_M1022_g 0.040726f $X=-0.33 $Y=1.885 $X2=4.465
+ $Y2=1.697
cc_137 N_VPB_c_91_p N_A_183_141#_M1022_g 0.0157621f $X=17.52 $Y=4.07 $X2=4.465
+ $Y2=1.697
cc_138 N_VPB_c_92_p N_A_183_141#_M1022_g 0.00970178f $X=17.52 $Y=4.07 $X2=4.465
+ $Y2=1.697
cc_139 N_VPB_M1000_b N_A_183_141#_M1025_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_140 N_VPB_c_91_p N_A_183_141#_M1025_g 0.0157621f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_141 N_VPB_c_92_p N_A_183_141#_M1025_g 0.00970178f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_142 N_VPB_M1000_b N_A_183_141#_M1031_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_143 N_VPB_c_91_p N_A_183_141#_M1031_g 0.0157621f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_144 N_VPB_c_92_p N_A_183_141#_M1031_g 0.00970178f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_145 N_VPB_M1000_b N_A_183_141#_M1033_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_146 N_VPB_c_91_p N_A_183_141#_M1033_g 0.0157621f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_147 N_VPB_c_92_p N_A_183_141#_M1033_g 0.00970178f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_148 N_VPB_M1000_b N_A_183_141#_M1038_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_149 N_VPB_c_91_p N_A_183_141#_M1038_g 0.0157621f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_150 N_VPB_c_92_p N_A_183_141#_M1038_g 0.00970178f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_151 N_VPB_M1000_b N_A_183_141#_M1039_g 0.040726f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_152 N_VPB_c_91_p N_A_183_141#_M1039_g 0.0157621f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_153 N_VPB_c_92_p N_A_183_141#_M1039_g 0.00970178f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_154 N_VPB_M1000_b N_A_183_141#_c_389_n 0.203856f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_155 N_VPB_M1000_b N_A_183_141#_M1042_g 0.0502706f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_156 N_VPB_c_91_p N_A_183_141#_M1042_g 0.0157621f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_157 N_VPB_c_92_p N_A_183_141#_M1042_g 0.00970178f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_158 N_VPB_M1000_b N_A_183_141#_c_457_n 0.00168525f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_159 N_VPB_c_91_p N_A_183_141#_c_457_n 0.0160222f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_160 N_VPB_c_92_p N_A_183_141#_c_457_n 0.00105499f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_161 N_VPB_M1000_b N_A_183_141#_c_460_n 0.00161463f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_162 N_VPB_c_91_p N_A_183_141#_c_460_n 0.0159826f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_163 N_VPB_c_92_p N_A_183_141#_c_460_n 0.00107233f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_164 N_VPB_M1000_b N_A_183_141#_c_463_n 0.00173328f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_165 N_VPB_c_91_p N_A_183_141#_c_463_n 0.0180171f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_166 N_VPB_c_92_p N_A_183_141#_c_463_n 0.00122962f $X=17.52 $Y=4.07 $X2=0
+ $Y2=0
cc_167 N_VPB_M1000_b N_VPWR_c_841_n 0.0644578f $X=-0.33 $Y=1.885 $X2=4.565
+ $Y2=2.965
cc_168 N_VPB_c_91_p N_VPWR_c_841_n 0.0289697f $X=17.52 $Y=4.07 $X2=4.565
+ $Y2=2.965
cc_169 N_VPB_c_92_p N_VPWR_c_841_n 0.00219871f $X=17.52 $Y=4.07 $X2=4.565
+ $Y2=2.965
cc_170 N_VPB_c_91_p N_VPWR_c_844_n 0.0306445f $X=17.52 $Y=4.07 $X2=3.515
+ $Y2=1.58
cc_171 N_VPB_c_92_p N_VPWR_c_844_n 0.00361083f $X=17.52 $Y=4.07 $X2=3.515
+ $Y2=1.58
cc_172 N_VPB_c_91_p N_VPWR_c_846_n 0.0306445f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_173 N_VPB_c_92_p N_VPWR_c_846_n 0.00361083f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_174 N_VPB_c_91_p N_VPWR_c_848_n 0.0306445f $X=17.52 $Y=4.07 $X2=0.385
+ $Y2=1.697
cc_175 N_VPB_c_92_p N_VPWR_c_848_n 0.00361083f $X=17.52 $Y=4.07 $X2=0.385
+ $Y2=1.697
cc_176 N_VPB_M1000_b N_VPWR_c_850_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_177 N_VPB_c_91_p N_VPWR_c_850_n 0.0445179f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_178 N_VPB_c_92_p N_VPWR_c_850_n 0.00377602f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_179 N_VPB_M1000_b N_VPWR_c_853_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_180 N_VPB_c_91_p N_VPWR_c_853_n 0.0445179f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_181 N_VPB_c_92_p N_VPWR_c_853_n 0.00377602f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_182 N_VPB_M1000_b N_VPWR_c_856_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_183 N_VPB_c_91_p N_VPWR_c_856_n 0.0445179f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_184 N_VPB_c_92_p N_VPWR_c_856_n 0.00377602f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_185 N_VPB_M1000_b N_VPWR_c_859_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_186 N_VPB_c_91_p N_VPWR_c_859_n 0.0445179f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_187 N_VPB_c_92_p N_VPWR_c_859_n 0.00377602f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_188 N_VPB_M1000_b N_VPWR_c_862_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_189 N_VPB_c_91_p N_VPWR_c_862_n 0.0445179f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_190 N_VPB_c_92_p N_VPWR_c_862_n 0.00377602f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_191 N_VPB_M1000_b N_VPWR_c_865_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_192 N_VPB_c_91_p N_VPWR_c_865_n 0.0445179f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_193 N_VPB_c_92_p N_VPWR_c_865_n 0.00377602f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_194 N_VPB_M1000_b N_VPWR_c_868_n 0.00369605f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_195 N_VPB_c_91_p N_VPWR_c_868_n 0.0445179f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_196 N_VPB_c_92_p N_VPWR_c_868_n 0.00377602f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_197 N_VPB_M1000_b N_VPWR_c_871_n 0.0633596f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_198 N_VPB_c_91_p N_VPWR_c_871_n 0.0270143f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_199 N_VPB_c_92_p N_VPWR_c_871_n 0.00200674f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_200 N_VPB_M1000_b N_VPWR_c_874_n 0.0647268f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_201 N_VPB_c_91_p N_VPWR_c_874_n 0.0770278f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_202 N_VPB_c_92_p N_VPWR_c_874_n 1.88095f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_203 N_VPB_M1000_b N_X_c_1046_n 0.00125033f $X=-0.33 $Y=1.885 $X2=4.465
+ $Y2=1.815
cc_204 N_VPB_c_91_p N_X_c_1046_n 0.0171423f $X=17.52 $Y=4.07 $X2=4.465 $Y2=1.815
cc_205 N_VPB_c_92_p N_X_c_1046_n 0.00108855f $X=17.52 $Y=4.07 $X2=4.465
+ $Y2=1.815
cc_206 N_VPB_M1000_b N_X_c_1049_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_207 N_VPB_c_91_p N_X_c_1049_n 0.0171423f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_208 N_VPB_c_92_p N_X_c_1049_n 0.00108855f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_209 N_VPB_M1000_b N_X_c_1052_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_210 N_VPB_c_91_p N_X_c_1052_n 0.0171423f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_211 N_VPB_c_92_p N_X_c_1052_n 0.00108855f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_212 N_VPB_M1000_b N_X_c_1055_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_213 N_VPB_c_91_p N_X_c_1055_n 0.0171423f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_214 N_VPB_c_92_p N_X_c_1055_n 0.00108855f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_215 N_VPB_M1000_b N_X_c_1058_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_216 N_VPB_c_91_p N_X_c_1058_n 0.0171423f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_217 N_VPB_c_92_p N_X_c_1058_n 0.00108855f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_218 N_VPB_M1000_b N_X_c_1061_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_219 N_VPB_c_91_p N_X_c_1061_n 0.0171423f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_220 N_VPB_c_92_p N_X_c_1061_n 0.00108855f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_221 N_VPB_M1000_b N_X_c_1064_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_222 N_VPB_c_91_p N_X_c_1064_n 0.0171423f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_223 N_VPB_c_92_p N_X_c_1064_n 0.00108855f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_224 N_VPB_M1000_b N_X_c_1067_n 0.00125033f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_225 N_VPB_c_91_p N_X_c_1067_n 0.0210531f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_226 N_VPB_c_92_p N_X_c_1067_n 0.00147247f $X=17.52 $Y=4.07 $X2=0 $Y2=0
cc_227 N_A_c_237_n N_A_183_141#_c_359_n 0.0243468f $X=4.565 $Y=1.565 $X2=0 $Y2=0
cc_228 N_A_M1036_g N_A_183_141#_M1001_g 0.0243468f $X=4.565 $Y=2.965 $X2=0 $Y2=0
cc_229 N_A_c_240_n N_A_183_141#_c_389_n 0.0243468f $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_230 N_A_c_227_n N_A_183_141#_c_391_n 0.012066f $X=0.665 $Y=1.565 $X2=0 $Y2=0
cc_231 N_A_M1000_g N_A_183_141#_c_457_n 0.0293976f $X=0.665 $Y=2.965 $X2=0 $Y2=0
cc_232 N_A_M1005_g N_A_183_141#_c_457_n 0.0022192f $X=1.445 $Y=2.965 $X2=0 $Y2=0
cc_233 N_A_M1005_g N_A_183_141#_c_472_n 0.0253301f $X=1.445 $Y=2.965 $X2=0 $Y2=0
cc_234 N_A_M1011_g N_A_183_141#_c_472_n 0.0218849f $X=2.225 $Y=2.965 $X2=0 $Y2=0
cc_235 N_A_c_239_n N_A_183_141#_c_472_n 0.0894665f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_236 N_A_c_240_n N_A_183_141#_c_472_n 0.0283643f $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_237 N_A_M1000_g N_A_183_141#_c_476_n 0.00954688f $X=0.665 $Y=2.965 $X2=0
+ $Y2=0
cc_238 N_A_c_239_n N_A_183_141#_c_476_n 0.024153f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_239 N_A_c_240_n N_A_183_141#_c_476_n 0.013297f $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_240 N_A_c_229_n N_A_183_141#_c_479_n 0.0276926f $X=1.445 $Y=1.565 $X2=0 $Y2=0
cc_241 N_A_c_231_n N_A_183_141#_c_479_n 0.0243589f $X=2.225 $Y=1.565 $X2=0 $Y2=0
cc_242 N_A_c_239_n N_A_183_141#_c_479_n 0.0824875f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_243 N_A_c_240_n N_A_183_141#_c_479_n 0.0024988f $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_244 N_A_c_227_n N_A_183_141#_c_483_n 0.00653924f $X=0.665 $Y=1.565 $X2=0
+ $Y2=0
cc_245 N_A_c_239_n N_A_183_141#_c_483_n 0.0242608f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_246 N_A_c_240_n N_A_183_141#_c_483_n 0.0025699f $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_247 N_A_c_231_n N_A_183_141#_c_392_n 0.0163015f $X=2.225 $Y=1.565 $X2=0 $Y2=0
cc_248 N_A_c_233_n N_A_183_141#_c_392_n 0.0139077f $X=3.005 $Y=1.565 $X2=0 $Y2=0
cc_249 N_A_M1011_g N_A_183_141#_c_460_n 0.0373895f $X=2.225 $Y=2.965 $X2=0 $Y2=0
cc_250 N_A_M1023_g N_A_183_141#_c_460_n 0.00215741f $X=3.005 $Y=2.965 $X2=0
+ $Y2=0
cc_251 N_A_M1023_g N_A_183_141#_c_490_n 0.0246803f $X=3.005 $Y=2.965 $X2=0 $Y2=0
cc_252 N_A_M1029_g N_A_183_141#_c_490_n 0.0212247f $X=3.785 $Y=2.965 $X2=0 $Y2=0
cc_253 N_A_c_239_n N_A_183_141#_c_490_n 0.0887444f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_254 N_A_c_240_n N_A_183_141#_c_490_n 0.02815f $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_255 N_A_c_233_n N_A_183_141#_c_494_n 0.026264f $X=3.005 $Y=1.565 $X2=0 $Y2=0
cc_256 N_A_c_235_n N_A_183_141#_c_494_n 0.0274546f $X=3.785 $Y=1.565 $X2=0 $Y2=0
cc_257 N_A_c_239_n N_A_183_141#_c_494_n 0.0837197f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_258 N_A_c_240_n N_A_183_141#_c_494_n 0.0024988f $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_259 N_A_M1023_g N_A_183_141#_c_463_n 8.05117e-19 $X=3.005 $Y=2.965 $X2=0
+ $Y2=0
cc_260 N_A_M1029_g N_A_183_141#_c_463_n 0.0361085f $X=3.785 $Y=2.965 $X2=0 $Y2=0
cc_261 N_A_M1036_g N_A_183_141#_c_463_n 0.00227089f $X=4.565 $Y=2.965 $X2=0
+ $Y2=0
cc_262 N_A_c_235_n N_A_183_141#_c_393_n 0.0119333f $X=3.785 $Y=1.565 $X2=0 $Y2=0
cc_263 N_A_c_237_n N_A_183_141#_c_502_n 0.0291623f $X=4.565 $Y=1.565 $X2=0 $Y2=0
cc_264 N_A_c_239_n N_A_183_141#_c_502_n 0.0238559f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_265 N_A_M1036_g N_A_183_141#_c_504_n 0.0253075f $X=4.565 $Y=2.965 $X2=0 $Y2=0
cc_266 N_A_c_239_n N_A_183_141#_c_504_n 0.0245146f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_267 N_A_c_240_n N_A_183_141#_c_504_n 0.0138465f $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_268 N_A_c_231_n N_A_183_141#_c_507_n 0.00255636f $X=2.225 $Y=1.565 $X2=0
+ $Y2=0
cc_269 N_A_c_233_n N_A_183_141#_c_507_n 0.00116671f $X=3.005 $Y=1.565 $X2=0
+ $Y2=0
cc_270 N_A_c_239_n N_A_183_141#_c_507_n 0.0259572f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_271 N_A_c_240_n N_A_183_141#_c_507_n 0.00257254f $X=4.565 $Y=1.815 $X2=0
+ $Y2=0
cc_272 N_A_M1011_g N_A_183_141#_c_511_n 0.00316841f $X=2.225 $Y=2.965 $X2=0
+ $Y2=0
cc_273 N_A_c_239_n N_A_183_141#_c_511_n 0.024153f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_274 N_A_c_240_n N_A_183_141#_c_511_n 0.00931804f $X=4.565 $Y=1.815 $X2=0
+ $Y2=0
cc_275 N_A_M1029_g N_A_183_141#_c_514_n 0.00354318f $X=3.785 $Y=2.965 $X2=0
+ $Y2=0
cc_276 N_A_c_239_n N_A_183_141#_c_514_n 0.0272695f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_277 N_A_c_240_n N_A_183_141#_c_514_n 0.0101992f $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_278 N_A_c_235_n N_A_183_141#_c_517_n 2.98176e-19 $X=3.785 $Y=1.565 $X2=0
+ $Y2=0
cc_279 N_A_c_239_n N_A_183_141#_c_517_n 0.0165976f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_280 N_A_c_240_n N_A_183_141#_c_517_n 0.00257254f $X=4.565 $Y=1.815 $X2=0
+ $Y2=0
cc_281 N_A_c_237_n N_A_183_141#_c_520_n 0.00112921f $X=4.565 $Y=1.565 $X2=0
+ $Y2=0
cc_282 N_A_c_239_n N_A_183_141#_c_520_n 0.00634454f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_283 N_A_c_240_n N_A_183_141#_c_520_n 0.00320764f $X=4.565 $Y=1.815 $X2=0
+ $Y2=0
cc_284 N_A_c_237_n N_A_183_141#_c_523_n 0.00894719f $X=4.565 $Y=1.565 $X2=0
+ $Y2=0
cc_285 N_A_c_239_n N_A_183_141#_c_523_n 0.0160237f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_286 N_A_c_240_n N_A_183_141#_c_523_n 0.0165299f $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_287 N_A_M1000_g N_VPWR_c_841_n 0.0688276f $X=0.665 $Y=2.965 $X2=0 $Y2=0
cc_288 N_A_c_239_n N_VPWR_c_841_n 0.0204297f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_289 N_A_c_240_n N_VPWR_c_841_n 0.00594552f $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_290 N_A_M1000_g N_VPWR_c_844_n 4.82782e-19 $X=0.665 $Y=2.965 $X2=0 $Y2=0
cc_291 N_A_M1005_g N_VPWR_c_844_n 0.0590539f $X=1.445 $Y=2.965 $X2=0 $Y2=0
cc_292 N_A_M1011_g N_VPWR_c_844_n 0.050844f $X=2.225 $Y=2.965 $X2=0 $Y2=0
cc_293 N_A_c_240_n N_VPWR_c_844_n 4.98839e-19 $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_294 N_A_M1011_g N_VPWR_c_846_n 4.84763e-19 $X=2.225 $Y=2.965 $X2=0 $Y2=0
cc_295 N_A_M1023_g N_VPWR_c_846_n 0.0609199f $X=3.005 $Y=2.965 $X2=0 $Y2=0
cc_296 N_A_M1029_g N_VPWR_c_846_n 0.0481049f $X=3.785 $Y=2.965 $X2=0 $Y2=0
cc_297 N_A_c_240_n N_VPWR_c_846_n 4.98839e-19 $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_298 N_A_M1029_g N_VPWR_c_848_n 4.5995e-19 $X=3.785 $Y=2.965 $X2=0 $Y2=0
cc_299 N_A_M1036_g N_VPWR_c_848_n 0.058787f $X=4.565 $Y=2.965 $X2=0 $Y2=0
cc_300 N_A_M1000_g N_VPWR_c_874_n 0.0100933f $X=0.665 $Y=2.965 $X2=0 $Y2=0
cc_301 N_A_M1005_g N_VPWR_c_874_n 0.00971346f $X=1.445 $Y=2.965 $X2=0 $Y2=0
cc_302 N_A_M1011_g N_VPWR_c_874_n 0.0104855f $X=2.225 $Y=2.965 $X2=0 $Y2=0
cc_303 N_A_M1023_g N_VPWR_c_874_n 0.00883212f $X=3.005 $Y=2.965 $X2=0 $Y2=0
cc_304 N_A_M1029_g N_VPWR_c_874_n 0.0104497f $X=3.785 $Y=2.965 $X2=0 $Y2=0
cc_305 N_A_M1036_g N_VPWR_c_874_n 0.00972336f $X=4.565 $Y=2.965 $X2=0 $Y2=0
cc_306 N_A_c_227_n N_VGND_c_1254_n 0.0413536f $X=0.665 $Y=1.565 $X2=0 $Y2=0
cc_307 N_A_c_229_n N_VGND_c_1254_n 8.88499e-19 $X=1.445 $Y=1.565 $X2=0 $Y2=0
cc_308 N_A_c_239_n N_VGND_c_1254_n 0.0309722f $X=4.465 $Y=1.73 $X2=0 $Y2=0
cc_309 N_A_c_240_n N_VGND_c_1254_n 0.0048454f $X=4.565 $Y=1.815 $X2=0 $Y2=0
cc_310 N_A_c_227_n N_VGND_c_1256_n 0.00101241f $X=0.665 $Y=1.565 $X2=0 $Y2=0
cc_311 N_A_c_229_n N_VGND_c_1256_n 0.0339149f $X=1.445 $Y=1.565 $X2=0 $Y2=0
cc_312 N_A_c_231_n N_VGND_c_1256_n 0.0281515f $X=2.225 $Y=1.565 $X2=0 $Y2=0
cc_313 N_A_c_233_n N_VGND_c_1256_n 7.4453e-19 $X=3.005 $Y=1.565 $X2=0 $Y2=0
cc_314 N_A_c_231_n N_VGND_c_1258_n 7.99935e-19 $X=2.225 $Y=1.565 $X2=0 $Y2=0
cc_315 N_A_c_233_n N_VGND_c_1258_n 0.0309163f $X=3.005 $Y=1.565 $X2=0 $Y2=0
cc_316 N_A_c_235_n N_VGND_c_1258_n 0.032189f $X=3.785 $Y=1.565 $X2=0 $Y2=0
cc_317 N_A_c_237_n N_VGND_c_1258_n 5.19551e-19 $X=4.565 $Y=1.565 $X2=0 $Y2=0
cc_318 N_A_c_235_n N_VGND_c_1260_n 5.04771e-19 $X=3.785 $Y=1.565 $X2=0 $Y2=0
cc_319 N_A_c_237_n N_VGND_c_1260_n 0.034076f $X=4.565 $Y=1.565 $X2=0 $Y2=0
cc_320 N_A_c_227_n N_VGND_c_1278_n 0.0127777f $X=0.665 $Y=1.565 $X2=0 $Y2=0
cc_321 N_A_c_229_n N_VGND_c_1278_n 0.00454157f $X=1.445 $Y=1.565 $X2=0 $Y2=0
cc_322 N_A_c_231_n N_VGND_c_1278_n 0.00710298f $X=2.225 $Y=1.565 $X2=0 $Y2=0
cc_323 N_A_c_233_n N_VGND_c_1278_n 0.00613925f $X=3.005 $Y=1.565 $X2=0 $Y2=0
cc_324 N_A_c_235_n N_VGND_c_1278_n 0.00553692f $X=3.785 $Y=1.565 $X2=0 $Y2=0
cc_325 N_A_c_237_n N_VGND_c_1278_n 0.00393066f $X=4.565 $Y=1.565 $X2=0 $Y2=0
cc_326 N_A_183_141#_c_472_n N_VPWR_M1005_d 0.00183555f $X=2.4 $Y=2.125 $X2=0
+ $Y2=0
cc_327 N_A_183_141#_c_490_n N_VPWR_M1023_d 0.00183555f $X=3.94 $Y=2.125 $X2=0
+ $Y2=0
cc_328 N_A_183_141#_c_504_n N_VPWR_M1036_d 0.00188202f $X=4.8 $Y=2.125 $X2=0
+ $Y2=0
cc_329 N_A_183_141#_c_457_n N_VPWR_c_841_n 0.112221f $X=1.055 $Y=2.34 $X2=0
+ $Y2=0
cc_330 N_A_183_141#_c_476_n N_VPWR_c_841_n 0.00747993f $X=1.16 $Y=2.125 $X2=0
+ $Y2=0
cc_331 N_A_183_141#_c_457_n N_VPWR_c_844_n 0.0510355f $X=1.055 $Y=2.34 $X2=0
+ $Y2=0
cc_332 N_A_183_141#_c_472_n N_VPWR_c_844_n 0.0591121f $X=2.4 $Y=2.125 $X2=0
+ $Y2=0
cc_333 N_A_183_141#_c_460_n N_VPWR_c_844_n 0.0941391f $X=2.615 $Y=2.34 $X2=0
+ $Y2=0
cc_334 N_A_183_141#_c_460_n N_VPWR_c_846_n 0.0536079f $X=2.615 $Y=2.34 $X2=0
+ $Y2=0
cc_335 N_A_183_141#_c_490_n N_VPWR_c_846_n 0.0591121f $X=3.94 $Y=2.125 $X2=0
+ $Y2=0
cc_336 N_A_183_141#_c_463_n N_VPWR_c_846_n 0.0948437f $X=4.175 $Y=2.34 $X2=0
+ $Y2=0
cc_337 N_A_183_141#_M1001_g N_VPWR_c_848_n 0.0532403f $X=5.345 $Y=2.965 $X2=0
+ $Y2=0
cc_338 N_A_183_141#_M1003_g N_VPWR_c_848_n 4.38254e-19 $X=6.125 $Y=2.965 $X2=0
+ $Y2=0
cc_339 N_A_183_141#_c_463_n N_VPWR_c_848_n 0.0536237f $X=4.175 $Y=2.34 $X2=0
+ $Y2=0
cc_340 N_A_183_141#_c_504_n N_VPWR_c_848_n 0.0614975f $X=4.8 $Y=2.125 $X2=0
+ $Y2=0
cc_341 N_A_183_141#_M1001_g N_VPWR_c_850_n 5.95094e-19 $X=5.345 $Y=2.965 $X2=0
+ $Y2=0
cc_342 N_A_183_141#_M1003_g N_VPWR_c_850_n 0.0732563f $X=6.125 $Y=2.965 $X2=0
+ $Y2=0
cc_343 N_A_183_141#_M1008_g N_VPWR_c_850_n 0.0734744f $X=6.905 $Y=2.965 $X2=0
+ $Y2=0
cc_344 N_A_183_141#_M1010_g N_VPWR_c_850_n 5.95094e-19 $X=7.685 $Y=2.965 $X2=0
+ $Y2=0
cc_345 N_A_183_141#_c_389_n N_VPWR_c_850_n 0.00264079f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_346 N_A_183_141#_c_546_p N_VPWR_c_850_n 0.0031325f $X=6.17 $Y=1.665 $X2=0
+ $Y2=0
cc_347 N_A_183_141#_c_547_p N_VPWR_c_850_n 0.00287695f $X=6.285 $Y=1.665 $X2=0
+ $Y2=0
cc_348 N_A_183_141#_c_395_n N_VPWR_c_850_n 0.0282532f $X=6.675 $Y=1.665 $X2=0
+ $Y2=0
cc_349 N_A_183_141#_c_549_p N_VPWR_c_850_n 0.0045029f $X=7.73 $Y=1.665 $X2=0
+ $Y2=0
cc_350 N_A_183_141#_M1008_g N_VPWR_c_853_n 5.95094e-19 $X=6.905 $Y=2.965 $X2=0
+ $Y2=0
cc_351 N_A_183_141#_M1010_g N_VPWR_c_853_n 0.0732563f $X=7.685 $Y=2.965 $X2=0
+ $Y2=0
cc_352 N_A_183_141#_M1012_g N_VPWR_c_853_n 0.0734744f $X=8.465 $Y=2.965 $X2=0
+ $Y2=0
cc_353 N_A_183_141#_M1013_g N_VPWR_c_853_n 5.95094e-19 $X=9.245 $Y=2.965 $X2=0
+ $Y2=0
cc_354 N_A_183_141#_c_389_n N_VPWR_c_853_n 0.00264079f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_355 N_A_183_141#_c_549_p N_VPWR_c_853_n 0.0031325f $X=7.73 $Y=1.665 $X2=0
+ $Y2=0
cc_356 N_A_183_141#_c_556_p N_VPWR_c_853_n 0.00287695f $X=7.845 $Y=1.665 $X2=0
+ $Y2=0
cc_357 N_A_183_141#_c_397_n N_VPWR_c_853_n 0.0282532f $X=8.235 $Y=1.665 $X2=0
+ $Y2=0
cc_358 N_A_183_141#_c_558_p N_VPWR_c_853_n 0.0045029f $X=9.29 $Y=1.665 $X2=0
+ $Y2=0
cc_359 N_A_183_141#_M1012_g N_VPWR_c_856_n 5.95094e-19 $X=8.465 $Y=2.965 $X2=0
+ $Y2=0
cc_360 N_A_183_141#_M1013_g N_VPWR_c_856_n 0.0732563f $X=9.245 $Y=2.965 $X2=0
+ $Y2=0
cc_361 N_A_183_141#_M1015_g N_VPWR_c_856_n 0.0734744f $X=10.025 $Y=2.965 $X2=0
+ $Y2=0
cc_362 N_A_183_141#_M1018_g N_VPWR_c_856_n 5.95094e-19 $X=10.805 $Y=2.965 $X2=0
+ $Y2=0
cc_363 N_A_183_141#_c_389_n N_VPWR_c_856_n 0.00264079f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_364 N_A_183_141#_c_558_p N_VPWR_c_856_n 0.0031325f $X=9.29 $Y=1.665 $X2=0
+ $Y2=0
cc_365 N_A_183_141#_c_565_p N_VPWR_c_856_n 0.00287695f $X=9.405 $Y=1.665 $X2=0
+ $Y2=0
cc_366 N_A_183_141#_c_399_n N_VPWR_c_856_n 0.0282532f $X=9.795 $Y=1.665 $X2=0
+ $Y2=0
cc_367 N_A_183_141#_c_567_p N_VPWR_c_856_n 0.0045029f $X=10.85 $Y=1.665 $X2=0
+ $Y2=0
cc_368 N_A_183_141#_M1015_g N_VPWR_c_859_n 5.95094e-19 $X=10.025 $Y=2.965 $X2=0
+ $Y2=0
cc_369 N_A_183_141#_M1018_g N_VPWR_c_859_n 0.0732563f $X=10.805 $Y=2.965 $X2=0
+ $Y2=0
cc_370 N_A_183_141#_M1021_g N_VPWR_c_859_n 0.0734744f $X=11.585 $Y=2.965 $X2=0
+ $Y2=0
cc_371 N_A_183_141#_M1022_g N_VPWR_c_859_n 5.95094e-19 $X=12.365 $Y=2.965 $X2=0
+ $Y2=0
cc_372 N_A_183_141#_c_389_n N_VPWR_c_859_n 0.00264079f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_373 N_A_183_141#_c_567_p N_VPWR_c_859_n 0.0031325f $X=10.85 $Y=1.665 $X2=0
+ $Y2=0
cc_374 N_A_183_141#_c_574_p N_VPWR_c_859_n 0.00287695f $X=10.965 $Y=1.665 $X2=0
+ $Y2=0
cc_375 N_A_183_141#_c_401_n N_VPWR_c_859_n 0.0282532f $X=11.355 $Y=1.665 $X2=0
+ $Y2=0
cc_376 N_A_183_141#_c_576_p N_VPWR_c_859_n 0.0045029f $X=12.41 $Y=1.665 $X2=0
+ $Y2=0
cc_377 N_A_183_141#_M1021_g N_VPWR_c_862_n 5.95094e-19 $X=11.585 $Y=2.965 $X2=0
+ $Y2=0
cc_378 N_A_183_141#_M1022_g N_VPWR_c_862_n 0.0732563f $X=12.365 $Y=2.965 $X2=0
+ $Y2=0
cc_379 N_A_183_141#_M1025_g N_VPWR_c_862_n 0.0734744f $X=13.145 $Y=2.965 $X2=0
+ $Y2=0
cc_380 N_A_183_141#_M1031_g N_VPWR_c_862_n 5.95094e-19 $X=13.925 $Y=2.965 $X2=0
+ $Y2=0
cc_381 N_A_183_141#_c_389_n N_VPWR_c_862_n 0.00264079f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_382 N_A_183_141#_c_576_p N_VPWR_c_862_n 0.0031325f $X=12.41 $Y=1.665 $X2=0
+ $Y2=0
cc_383 N_A_183_141#_c_583_p N_VPWR_c_862_n 0.00287695f $X=12.525 $Y=1.665 $X2=0
+ $Y2=0
cc_384 N_A_183_141#_c_403_n N_VPWR_c_862_n 0.0282532f $X=12.915 $Y=1.665 $X2=0
+ $Y2=0
cc_385 N_A_183_141#_c_585_p N_VPWR_c_862_n 0.0045029f $X=13.97 $Y=1.665 $X2=0
+ $Y2=0
cc_386 N_A_183_141#_M1025_g N_VPWR_c_865_n 5.95094e-19 $X=13.145 $Y=2.965 $X2=0
+ $Y2=0
cc_387 N_A_183_141#_M1031_g N_VPWR_c_865_n 0.0732563f $X=13.925 $Y=2.965 $X2=0
+ $Y2=0
cc_388 N_A_183_141#_M1033_g N_VPWR_c_865_n 0.0734744f $X=14.705 $Y=2.965 $X2=0
+ $Y2=0
cc_389 N_A_183_141#_M1038_g N_VPWR_c_865_n 5.95094e-19 $X=15.485 $Y=2.965 $X2=0
+ $Y2=0
cc_390 N_A_183_141#_c_389_n N_VPWR_c_865_n 0.00264079f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_391 N_A_183_141#_c_585_p N_VPWR_c_865_n 0.0031325f $X=13.97 $Y=1.665 $X2=0
+ $Y2=0
cc_392 N_A_183_141#_c_592_p N_VPWR_c_865_n 0.00287695f $X=14.085 $Y=1.665 $X2=0
+ $Y2=0
cc_393 N_A_183_141#_c_405_n N_VPWR_c_865_n 0.0282532f $X=14.475 $Y=1.665 $X2=0
+ $Y2=0
cc_394 N_A_183_141#_c_594_p N_VPWR_c_865_n 0.0045029f $X=15.53 $Y=1.665 $X2=0
+ $Y2=0
cc_395 N_A_183_141#_M1033_g N_VPWR_c_868_n 5.95094e-19 $X=14.705 $Y=2.965 $X2=0
+ $Y2=0
cc_396 N_A_183_141#_M1038_g N_VPWR_c_868_n 0.0732563f $X=15.485 $Y=2.965 $X2=0
+ $Y2=0
cc_397 N_A_183_141#_M1039_g N_VPWR_c_868_n 0.0753959f $X=16.265 $Y=2.965 $X2=0
+ $Y2=0
cc_398 N_A_183_141#_c_389_n N_VPWR_c_868_n 0.00264079f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_399 N_A_183_141#_M1042_g N_VPWR_c_868_n 5.95094e-19 $X=17.045 $Y=2.965 $X2=0
+ $Y2=0
cc_400 N_A_183_141#_c_594_p N_VPWR_c_868_n 0.0031325f $X=15.53 $Y=1.665 $X2=0
+ $Y2=0
cc_401 N_A_183_141#_c_601_p N_VPWR_c_868_n 0.00287695f $X=15.645 $Y=1.665 $X2=0
+ $Y2=0
cc_402 N_A_183_141#_c_406_n N_VPWR_c_868_n 0.0021415f $X=16.035 $Y=1.665 $X2=0
+ $Y2=0
cc_403 N_A_183_141#_c_407_n N_VPWR_c_868_n 0.0282532f $X=16.035 $Y=1.665 $X2=0
+ $Y2=0
cc_404 N_A_183_141#_M1039_g N_VPWR_c_871_n 4.37802e-19 $X=16.265 $Y=2.965 $X2=0
+ $Y2=0
cc_405 N_A_183_141#_M1042_g N_VPWR_c_871_n 0.0636473f $X=17.045 $Y=2.965 $X2=0
+ $Y2=0
cc_406 N_A_183_141#_M1000_s N_VPWR_c_874_n 0.00137624f $X=0.915 $Y=2.215 $X2=0
+ $Y2=0
cc_407 N_A_183_141#_M1011_s N_VPWR_c_874_n 0.00179328f $X=2.475 $Y=2.215 $X2=0
+ $Y2=0
cc_408 N_A_183_141#_M1029_s N_VPWR_c_874_n 9.59196e-19 $X=4.035 $Y=2.215 $X2=0
+ $Y2=0
cc_409 N_A_183_141#_M1001_g N_VPWR_c_874_n 0.0131764f $X=5.345 $Y=2.965 $X2=0
+ $Y2=0
cc_410 N_A_183_141#_M1003_g N_VPWR_c_874_n 0.00965647f $X=6.125 $Y=2.965 $X2=0
+ $Y2=0
cc_411 N_A_183_141#_M1008_g N_VPWR_c_874_n 0.00965647f $X=6.905 $Y=2.965 $X2=0
+ $Y2=0
cc_412 N_A_183_141#_M1010_g N_VPWR_c_874_n 0.00965647f $X=7.685 $Y=2.965 $X2=0
+ $Y2=0
cc_413 N_A_183_141#_M1012_g N_VPWR_c_874_n 0.00965647f $X=8.465 $Y=2.965 $X2=0
+ $Y2=0
cc_414 N_A_183_141#_M1013_g N_VPWR_c_874_n 0.00965647f $X=9.245 $Y=2.965 $X2=0
+ $Y2=0
cc_415 N_A_183_141#_M1015_g N_VPWR_c_874_n 0.00965647f $X=10.025 $Y=2.965 $X2=0
+ $Y2=0
cc_416 N_A_183_141#_M1018_g N_VPWR_c_874_n 0.00965647f $X=10.805 $Y=2.965 $X2=0
+ $Y2=0
cc_417 N_A_183_141#_M1021_g N_VPWR_c_874_n 0.00965647f $X=11.585 $Y=2.965 $X2=0
+ $Y2=0
cc_418 N_A_183_141#_M1022_g N_VPWR_c_874_n 0.00965647f $X=12.365 $Y=2.965 $X2=0
+ $Y2=0
cc_419 N_A_183_141#_M1025_g N_VPWR_c_874_n 0.00965647f $X=13.145 $Y=2.965 $X2=0
+ $Y2=0
cc_420 N_A_183_141#_M1031_g N_VPWR_c_874_n 0.00965647f $X=13.925 $Y=2.965 $X2=0
+ $Y2=0
cc_421 N_A_183_141#_M1033_g N_VPWR_c_874_n 0.00965647f $X=14.705 $Y=2.965 $X2=0
+ $Y2=0
cc_422 N_A_183_141#_M1038_g N_VPWR_c_874_n 0.00965647f $X=15.485 $Y=2.965 $X2=0
+ $Y2=0
cc_423 N_A_183_141#_M1039_g N_VPWR_c_874_n 0.00965647f $X=16.265 $Y=2.965 $X2=0
+ $Y2=0
cc_424 N_A_183_141#_M1042_g N_VPWR_c_874_n 0.0101127f $X=17.045 $Y=2.965 $X2=0
+ $Y2=0
cc_425 N_A_183_141#_c_457_n N_VPWR_c_874_n 0.0381773f $X=1.055 $Y=2.34 $X2=0
+ $Y2=0
cc_426 N_A_183_141#_c_460_n N_VPWR_c_874_n 0.0394745f $X=2.615 $Y=2.34 $X2=0
+ $Y2=0
cc_427 N_A_183_141#_c_463_n N_VPWR_c_874_n 0.043412f $X=4.175 $Y=2.34 $X2=0
+ $Y2=0
cc_428 N_A_183_141#_c_359_n N_X_c_1046_n 0.0208809f $X=5.345 $Y=1.565 $X2=0
+ $Y2=0
cc_429 N_A_183_141#_M1001_g N_X_c_1046_n 0.0402736f $X=5.345 $Y=2.965 $X2=0
+ $Y2=0
cc_430 N_A_183_141#_c_361_n N_X_c_1046_n 0.0190601f $X=6.125 $Y=1.565 $X2=0
+ $Y2=0
cc_431 N_A_183_141#_M1003_g N_X_c_1046_n 0.0345177f $X=6.125 $Y=2.965 $X2=0
+ $Y2=0
cc_432 N_A_183_141#_c_389_n N_X_c_1046_n 0.0345088f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_433 N_A_183_141#_c_502_n N_X_c_1046_n 0.01395f $X=4.8 $Y=1.302 $X2=0 $Y2=0
cc_434 N_A_183_141#_c_504_n N_X_c_1046_n 0.0181025f $X=4.8 $Y=2.125 $X2=0 $Y2=0
cc_435 N_A_183_141#_c_546_p N_X_c_1046_n 0.0387052f $X=6.17 $Y=1.665 $X2=0 $Y2=0
cc_436 N_A_183_141#_c_636_p N_X_c_1046_n 0.00164429f $X=5.36 $Y=1.665 $X2=0
+ $Y2=0
cc_437 N_A_183_141#_c_547_p N_X_c_1046_n 9.02799e-19 $X=6.285 $Y=1.665 $X2=0
+ $Y2=0
cc_438 N_A_183_141#_c_395_n N_X_c_1046_n 0.0155872f $X=6.675 $Y=1.665 $X2=0
+ $Y2=0
cc_439 N_A_183_141#_c_523_n N_X_c_1046_n 0.0330205f $X=5.245 $Y=1.665 $X2=0
+ $Y2=0
cc_440 N_A_183_141#_c_363_n N_X_c_1049_n 0.0190713f $X=6.905 $Y=1.565 $X2=0
+ $Y2=0
cc_441 N_A_183_141#_M1008_g N_X_c_1049_n 0.0345177f $X=6.905 $Y=2.965 $X2=0
+ $Y2=0
cc_442 N_A_183_141#_c_365_n N_X_c_1049_n 0.0190601f $X=7.685 $Y=1.565 $X2=0
+ $Y2=0
cc_443 N_A_183_141#_M1010_g N_X_c_1049_n 0.0345177f $X=7.685 $Y=2.965 $X2=0
+ $Y2=0
cc_444 N_A_183_141#_c_389_n N_X_c_1049_n 0.0389693f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_445 N_A_183_141#_c_395_n N_X_c_1049_n 0.0135035f $X=6.675 $Y=1.665 $X2=0
+ $Y2=0
cc_446 N_A_183_141#_c_549_p N_X_c_1049_n 0.0392608f $X=7.73 $Y=1.665 $X2=0 $Y2=0
cc_447 N_A_183_141#_c_647_p N_X_c_1049_n 8.70571e-19 $X=6.82 $Y=1.665 $X2=0
+ $Y2=0
cc_448 N_A_183_141#_c_556_p N_X_c_1049_n 9.02799e-19 $X=7.845 $Y=1.665 $X2=0
+ $Y2=0
cc_449 N_A_183_141#_c_397_n N_X_c_1049_n 0.0155872f $X=8.235 $Y=1.665 $X2=0
+ $Y2=0
cc_450 N_A_183_141#_c_367_n N_X_c_1052_n 0.0190713f $X=8.465 $Y=1.565 $X2=0
+ $Y2=0
cc_451 N_A_183_141#_M1012_g N_X_c_1052_n 0.0345177f $X=8.465 $Y=2.965 $X2=0
+ $Y2=0
cc_452 N_A_183_141#_c_369_n N_X_c_1052_n 0.0190601f $X=9.245 $Y=1.565 $X2=0
+ $Y2=0
cc_453 N_A_183_141#_M1013_g N_X_c_1052_n 0.0345177f $X=9.245 $Y=2.965 $X2=0
+ $Y2=0
cc_454 N_A_183_141#_c_389_n N_X_c_1052_n 0.0389693f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_455 N_A_183_141#_c_397_n N_X_c_1052_n 0.0135035f $X=8.235 $Y=1.665 $X2=0
+ $Y2=0
cc_456 N_A_183_141#_c_558_p N_X_c_1052_n 0.0392608f $X=9.29 $Y=1.665 $X2=0 $Y2=0
cc_457 N_A_183_141#_c_657_p N_X_c_1052_n 8.70571e-19 $X=8.38 $Y=1.665 $X2=0
+ $Y2=0
cc_458 N_A_183_141#_c_565_p N_X_c_1052_n 9.02799e-19 $X=9.405 $Y=1.665 $X2=0
+ $Y2=0
cc_459 N_A_183_141#_c_399_n N_X_c_1052_n 0.0155872f $X=9.795 $Y=1.665 $X2=0
+ $Y2=0
cc_460 N_A_183_141#_c_371_n N_X_c_1055_n 0.0190713f $X=10.025 $Y=1.565 $X2=0
+ $Y2=0
cc_461 N_A_183_141#_M1015_g N_X_c_1055_n 0.0345177f $X=10.025 $Y=2.965 $X2=0
+ $Y2=0
cc_462 N_A_183_141#_c_373_n N_X_c_1055_n 0.0190601f $X=10.805 $Y=1.565 $X2=0
+ $Y2=0
cc_463 N_A_183_141#_M1018_g N_X_c_1055_n 0.0345177f $X=10.805 $Y=2.965 $X2=0
+ $Y2=0
cc_464 N_A_183_141#_c_389_n N_X_c_1055_n 0.0389693f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_465 N_A_183_141#_c_399_n N_X_c_1055_n 0.0135035f $X=9.795 $Y=1.665 $X2=0
+ $Y2=0
cc_466 N_A_183_141#_c_567_p N_X_c_1055_n 0.0392608f $X=10.85 $Y=1.665 $X2=0
+ $Y2=0
cc_467 N_A_183_141#_c_667_p N_X_c_1055_n 8.70571e-19 $X=9.94 $Y=1.665 $X2=0
+ $Y2=0
cc_468 N_A_183_141#_c_574_p N_X_c_1055_n 9.02799e-19 $X=10.965 $Y=1.665 $X2=0
+ $Y2=0
cc_469 N_A_183_141#_c_401_n N_X_c_1055_n 0.0155872f $X=11.355 $Y=1.665 $X2=0
+ $Y2=0
cc_470 N_A_183_141#_c_375_n N_X_c_1058_n 0.0190713f $X=11.585 $Y=1.565 $X2=0
+ $Y2=0
cc_471 N_A_183_141#_M1021_g N_X_c_1058_n 0.0345177f $X=11.585 $Y=2.965 $X2=0
+ $Y2=0
cc_472 N_A_183_141#_c_377_n N_X_c_1058_n 0.0190601f $X=12.365 $Y=1.565 $X2=0
+ $Y2=0
cc_473 N_A_183_141#_M1022_g N_X_c_1058_n 0.0345177f $X=12.365 $Y=2.965 $X2=0
+ $Y2=0
cc_474 N_A_183_141#_c_389_n N_X_c_1058_n 0.0389693f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_475 N_A_183_141#_c_401_n N_X_c_1058_n 0.0135035f $X=11.355 $Y=1.665 $X2=0
+ $Y2=0
cc_476 N_A_183_141#_c_576_p N_X_c_1058_n 0.0392608f $X=12.41 $Y=1.665 $X2=0
+ $Y2=0
cc_477 N_A_183_141#_c_677_p N_X_c_1058_n 8.70571e-19 $X=11.5 $Y=1.665 $X2=0
+ $Y2=0
cc_478 N_A_183_141#_c_583_p N_X_c_1058_n 9.02799e-19 $X=12.525 $Y=1.665 $X2=0
+ $Y2=0
cc_479 N_A_183_141#_c_403_n N_X_c_1058_n 0.0155872f $X=12.915 $Y=1.665 $X2=0
+ $Y2=0
cc_480 N_A_183_141#_c_379_n N_X_c_1061_n 0.0190713f $X=13.145 $Y=1.565 $X2=0
+ $Y2=0
cc_481 N_A_183_141#_M1025_g N_X_c_1061_n 0.0345177f $X=13.145 $Y=2.965 $X2=0
+ $Y2=0
cc_482 N_A_183_141#_c_381_n N_X_c_1061_n 0.0190601f $X=13.925 $Y=1.565 $X2=0
+ $Y2=0
cc_483 N_A_183_141#_M1031_g N_X_c_1061_n 0.0345177f $X=13.925 $Y=2.965 $X2=0
+ $Y2=0
cc_484 N_A_183_141#_c_389_n N_X_c_1061_n 0.0389693f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_485 N_A_183_141#_c_403_n N_X_c_1061_n 0.0135035f $X=12.915 $Y=1.665 $X2=0
+ $Y2=0
cc_486 N_A_183_141#_c_585_p N_X_c_1061_n 0.0392608f $X=13.97 $Y=1.665 $X2=0
+ $Y2=0
cc_487 N_A_183_141#_c_687_p N_X_c_1061_n 8.70571e-19 $X=13.06 $Y=1.665 $X2=0
+ $Y2=0
cc_488 N_A_183_141#_c_592_p N_X_c_1061_n 9.02799e-19 $X=14.085 $Y=1.665 $X2=0
+ $Y2=0
cc_489 N_A_183_141#_c_405_n N_X_c_1061_n 0.0155872f $X=14.475 $Y=1.665 $X2=0
+ $Y2=0
cc_490 N_A_183_141#_c_383_n N_X_c_1064_n 0.0190713f $X=14.705 $Y=1.565 $X2=0
+ $Y2=0
cc_491 N_A_183_141#_M1033_g N_X_c_1064_n 0.0345177f $X=14.705 $Y=2.965 $X2=0
+ $Y2=0
cc_492 N_A_183_141#_c_385_n N_X_c_1064_n 0.0190601f $X=15.485 $Y=1.565 $X2=0
+ $Y2=0
cc_493 N_A_183_141#_M1038_g N_X_c_1064_n 0.0345177f $X=15.485 $Y=2.965 $X2=0
+ $Y2=0
cc_494 N_A_183_141#_c_389_n N_X_c_1064_n 0.0389693f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_495 N_A_183_141#_c_405_n N_X_c_1064_n 0.0135035f $X=14.475 $Y=1.665 $X2=0
+ $Y2=0
cc_496 N_A_183_141#_c_594_p N_X_c_1064_n 0.0392608f $X=15.53 $Y=1.665 $X2=0
+ $Y2=0
cc_497 N_A_183_141#_c_697_p N_X_c_1064_n 8.70571e-19 $X=14.62 $Y=1.665 $X2=0
+ $Y2=0
cc_498 N_A_183_141#_c_601_p N_X_c_1064_n 9.02799e-19 $X=15.645 $Y=1.665 $X2=0
+ $Y2=0
cc_499 N_A_183_141#_c_407_n N_X_c_1064_n 0.0155872f $X=16.035 $Y=1.665 $X2=0
+ $Y2=0
cc_500 N_A_183_141#_c_387_n N_X_c_1067_n 0.01933f $X=16.265 $Y=1.565 $X2=0 $Y2=0
cc_501 N_A_183_141#_M1039_g N_X_c_1067_n 0.0348483f $X=16.265 $Y=2.965 $X2=0
+ $Y2=0
cc_502 N_A_183_141#_c_389_n N_X_c_1067_n 0.0769778f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_503 N_A_183_141#_M1042_g N_X_c_1067_n 0.0494075f $X=17.045 $Y=2.965 $X2=0
+ $Y2=0
cc_504 N_A_183_141#_c_406_n N_X_c_1067_n 0.00574079f $X=16.035 $Y=1.665 $X2=0
+ $Y2=0
cc_505 N_A_183_141#_c_407_n N_X_c_1067_n 0.0134415f $X=16.035 $Y=1.665 $X2=0
+ $Y2=0
cc_506 N_A_183_141#_M1003_g N_X_c_1148_n 0.014391f $X=6.125 $Y=2.965 $X2=0 $Y2=0
cc_507 N_A_183_141#_M1008_g N_X_c_1148_n 0.014391f $X=6.905 $Y=2.965 $X2=0 $Y2=0
cc_508 N_A_183_141#_c_547_p N_X_c_1148_n 0.0256666f $X=6.285 $Y=1.665 $X2=0
+ $Y2=0
cc_509 N_A_183_141#_c_395_n N_X_c_1148_n 0.00234231f $X=6.675 $Y=1.665 $X2=0
+ $Y2=0
cc_510 N_A_183_141#_c_546_p N_X_c_1152_n 0.0114767f $X=6.17 $Y=1.665 $X2=0 $Y2=0
cc_511 N_A_183_141#_M1010_g N_X_c_1153_n 0.014391f $X=7.685 $Y=2.965 $X2=0 $Y2=0
cc_512 N_A_183_141#_M1012_g N_X_c_1153_n 0.014391f $X=8.465 $Y=2.965 $X2=0 $Y2=0
cc_513 N_A_183_141#_c_556_p N_X_c_1153_n 0.0256666f $X=7.845 $Y=1.665 $X2=0
+ $Y2=0
cc_514 N_A_183_141#_c_397_n N_X_c_1153_n 0.00234231f $X=8.235 $Y=1.665 $X2=0
+ $Y2=0
cc_515 N_A_183_141#_c_549_p N_X_c_1157_n 0.0114767f $X=7.73 $Y=1.665 $X2=0 $Y2=0
cc_516 N_A_183_141#_M1013_g N_X_c_1158_n 0.014391f $X=9.245 $Y=2.965 $X2=0 $Y2=0
cc_517 N_A_183_141#_M1015_g N_X_c_1158_n 0.014391f $X=10.025 $Y=2.965 $X2=0
+ $Y2=0
cc_518 N_A_183_141#_c_565_p N_X_c_1158_n 0.0256666f $X=9.405 $Y=1.665 $X2=0
+ $Y2=0
cc_519 N_A_183_141#_c_399_n N_X_c_1158_n 0.00234231f $X=9.795 $Y=1.665 $X2=0
+ $Y2=0
cc_520 N_A_183_141#_c_558_p N_X_c_1162_n 0.0114767f $X=9.29 $Y=1.665 $X2=0 $Y2=0
cc_521 N_A_183_141#_M1018_g N_X_c_1163_n 0.014391f $X=10.805 $Y=2.965 $X2=0
+ $Y2=0
cc_522 N_A_183_141#_M1021_g N_X_c_1163_n 0.014391f $X=11.585 $Y=2.965 $X2=0
+ $Y2=0
cc_523 N_A_183_141#_c_574_p N_X_c_1163_n 0.0256666f $X=10.965 $Y=1.665 $X2=0
+ $Y2=0
cc_524 N_A_183_141#_c_401_n N_X_c_1163_n 0.00234231f $X=11.355 $Y=1.665 $X2=0
+ $Y2=0
cc_525 N_A_183_141#_c_567_p N_X_c_1167_n 0.0114767f $X=10.85 $Y=1.665 $X2=0
+ $Y2=0
cc_526 N_A_183_141#_M1022_g N_X_c_1168_n 0.014391f $X=12.365 $Y=2.965 $X2=0
+ $Y2=0
cc_527 N_A_183_141#_M1025_g N_X_c_1168_n 0.014391f $X=13.145 $Y=2.965 $X2=0
+ $Y2=0
cc_528 N_A_183_141#_c_583_p N_X_c_1168_n 0.0256666f $X=12.525 $Y=1.665 $X2=0
+ $Y2=0
cc_529 N_A_183_141#_c_403_n N_X_c_1168_n 0.00234231f $X=12.915 $Y=1.665 $X2=0
+ $Y2=0
cc_530 N_A_183_141#_c_576_p N_X_c_1172_n 0.0114767f $X=12.41 $Y=1.665 $X2=0
+ $Y2=0
cc_531 N_A_183_141#_M1031_g N_X_c_1173_n 0.014391f $X=13.925 $Y=2.965 $X2=0
+ $Y2=0
cc_532 N_A_183_141#_M1033_g N_X_c_1173_n 0.014391f $X=14.705 $Y=2.965 $X2=0
+ $Y2=0
cc_533 N_A_183_141#_c_592_p N_X_c_1173_n 0.0256666f $X=14.085 $Y=1.665 $X2=0
+ $Y2=0
cc_534 N_A_183_141#_c_405_n N_X_c_1173_n 0.00234231f $X=14.475 $Y=1.665 $X2=0
+ $Y2=0
cc_535 N_A_183_141#_c_585_p N_X_c_1177_n 0.0114767f $X=13.97 $Y=1.665 $X2=0
+ $Y2=0
cc_536 N_A_183_141#_M1038_g N_X_c_1178_n 0.014391f $X=15.485 $Y=2.965 $X2=0
+ $Y2=0
cc_537 N_A_183_141#_M1039_g N_X_c_1178_n 0.014391f $X=16.265 $Y=2.965 $X2=0
+ $Y2=0
cc_538 N_A_183_141#_c_601_p N_X_c_1178_n 0.0256666f $X=15.645 $Y=1.665 $X2=0
+ $Y2=0
cc_539 N_A_183_141#_c_407_n N_X_c_1178_n 0.00234231f $X=16.035 $Y=1.665 $X2=0
+ $Y2=0
cc_540 N_A_183_141#_c_594_p N_X_c_1182_n 0.0114767f $X=15.53 $Y=1.665 $X2=0
+ $Y2=0
cc_541 N_A_183_141#_c_479_n N_VGND_M1016_d 0.00329714f $X=2.4 $Y=1.302 $X2=0
+ $Y2=0
cc_542 N_A_183_141#_c_494_n N_VGND_M1026_d 0.00329714f $X=4.025 $Y=1.302 $X2=0
+ $Y2=0
cc_543 N_A_183_141#_c_502_n N_VGND_M1043_d 0.00180843f $X=4.8 $Y=1.302 $X2=0
+ $Y2=0
cc_544 N_A_183_141#_c_391_n N_VGND_c_1254_n 0.0344333f $X=1.055 $Y=0.92 $X2=0
+ $Y2=0
cc_545 N_A_183_141#_c_483_n N_VGND_c_1254_n 0.0177838f $X=1.17 $Y=1.302 $X2=0
+ $Y2=0
cc_546 N_A_183_141#_c_479_n N_VGND_c_1256_n 0.058686f $X=2.4 $Y=1.302 $X2=0
+ $Y2=0
cc_547 N_A_183_141#_c_392_n N_VGND_c_1256_n 0.0237236f $X=2.615 $Y=0.895 $X2=0
+ $Y2=0
cc_548 N_A_183_141#_c_392_n N_VGND_c_1258_n 0.0237236f $X=2.615 $Y=0.895 $X2=0
+ $Y2=0
cc_549 N_A_183_141#_c_494_n N_VGND_c_1258_n 0.0589786f $X=4.025 $Y=1.302 $X2=0
+ $Y2=0
cc_550 N_A_183_141#_c_393_n N_VGND_c_1258_n 0.0229431f $X=4.175 $Y=0.895 $X2=0
+ $Y2=0
cc_551 N_A_183_141#_c_359_n N_VGND_c_1260_n 0.027438f $X=5.345 $Y=1.565 $X2=0
+ $Y2=0
cc_552 N_A_183_141#_c_361_n N_VGND_c_1260_n 9.65869e-19 $X=6.125 $Y=1.565 $X2=0
+ $Y2=0
cc_553 N_A_183_141#_c_502_n N_VGND_c_1260_n 0.0602028f $X=4.8 $Y=1.302 $X2=0
+ $Y2=0
cc_554 N_A_183_141#_c_520_n N_VGND_c_1260_n 0.00218255f $X=5.245 $Y=1.665 $X2=0
+ $Y2=0
cc_555 N_A_183_141#_c_359_n N_VGND_c_1262_n 0.00109327f $X=5.345 $Y=1.565 $X2=0
+ $Y2=0
cc_556 N_A_183_141#_c_361_n N_VGND_c_1262_n 0.0476133f $X=6.125 $Y=1.565 $X2=0
+ $Y2=0
cc_557 N_A_183_141#_c_363_n N_VGND_c_1262_n 0.04751f $X=6.905 $Y=1.565 $X2=0
+ $Y2=0
cc_558 N_A_183_141#_c_365_n N_VGND_c_1262_n 6.39245e-19 $X=7.685 $Y=1.565 $X2=0
+ $Y2=0
cc_559 N_A_183_141#_c_389_n N_VGND_c_1262_n 7.87968e-19 $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_560 N_A_183_141#_c_546_p N_VGND_c_1262_n 0.00410965f $X=6.17 $Y=1.665 $X2=0
+ $Y2=0
cc_561 N_A_183_141#_c_547_p N_VGND_c_1262_n 0.0171054f $X=6.285 $Y=1.665 $X2=0
+ $Y2=0
cc_562 N_A_183_141#_c_395_n N_VGND_c_1262_n 0.041453f $X=6.675 $Y=1.665 $X2=0
+ $Y2=0
cc_563 N_A_183_141#_c_549_p N_VGND_c_1262_n 0.00590701f $X=7.73 $Y=1.665 $X2=0
+ $Y2=0
cc_564 N_A_183_141#_c_363_n N_VGND_c_1264_n 6.39245e-19 $X=6.905 $Y=1.565 $X2=0
+ $Y2=0
cc_565 N_A_183_141#_c_365_n N_VGND_c_1264_n 0.0473216f $X=7.685 $Y=1.565 $X2=0
+ $Y2=0
cc_566 N_A_183_141#_c_367_n N_VGND_c_1264_n 0.04751f $X=8.465 $Y=1.565 $X2=0
+ $Y2=0
cc_567 N_A_183_141#_c_369_n N_VGND_c_1264_n 6.39245e-19 $X=9.245 $Y=1.565 $X2=0
+ $Y2=0
cc_568 N_A_183_141#_c_389_n N_VGND_c_1264_n 7.87968e-19 $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_569 N_A_183_141#_c_549_p N_VGND_c_1264_n 0.00410965f $X=7.73 $Y=1.665 $X2=0
+ $Y2=0
cc_570 N_A_183_141#_c_556_p N_VGND_c_1264_n 0.0171054f $X=7.845 $Y=1.665 $X2=0
+ $Y2=0
cc_571 N_A_183_141#_c_397_n N_VGND_c_1264_n 0.041453f $X=8.235 $Y=1.665 $X2=0
+ $Y2=0
cc_572 N_A_183_141#_c_558_p N_VGND_c_1264_n 0.00590701f $X=9.29 $Y=1.665 $X2=0
+ $Y2=0
cc_573 N_A_183_141#_c_367_n N_VGND_c_1266_n 6.39245e-19 $X=8.465 $Y=1.565 $X2=0
+ $Y2=0
cc_574 N_A_183_141#_c_369_n N_VGND_c_1266_n 0.0473216f $X=9.245 $Y=1.565 $X2=0
+ $Y2=0
cc_575 N_A_183_141#_c_371_n N_VGND_c_1266_n 0.04751f $X=10.025 $Y=1.565 $X2=0
+ $Y2=0
cc_576 N_A_183_141#_c_373_n N_VGND_c_1266_n 6.39245e-19 $X=10.805 $Y=1.565 $X2=0
+ $Y2=0
cc_577 N_A_183_141#_c_389_n N_VGND_c_1266_n 7.87968e-19 $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_578 N_A_183_141#_c_558_p N_VGND_c_1266_n 0.00410965f $X=9.29 $Y=1.665 $X2=0
+ $Y2=0
cc_579 N_A_183_141#_c_565_p N_VGND_c_1266_n 0.0171054f $X=9.405 $Y=1.665 $X2=0
+ $Y2=0
cc_580 N_A_183_141#_c_399_n N_VGND_c_1266_n 0.041453f $X=9.795 $Y=1.665 $X2=0
+ $Y2=0
cc_581 N_A_183_141#_c_567_p N_VGND_c_1266_n 0.00590701f $X=10.85 $Y=1.665 $X2=0
+ $Y2=0
cc_582 N_A_183_141#_c_371_n N_VGND_c_1268_n 6.39245e-19 $X=10.025 $Y=1.565 $X2=0
+ $Y2=0
cc_583 N_A_183_141#_c_373_n N_VGND_c_1268_n 0.0473216f $X=10.805 $Y=1.565 $X2=0
+ $Y2=0
cc_584 N_A_183_141#_c_375_n N_VGND_c_1268_n 0.04751f $X=11.585 $Y=1.565 $X2=0
+ $Y2=0
cc_585 N_A_183_141#_c_377_n N_VGND_c_1268_n 6.39245e-19 $X=12.365 $Y=1.565 $X2=0
+ $Y2=0
cc_586 N_A_183_141#_c_389_n N_VGND_c_1268_n 7.87968e-19 $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_587 N_A_183_141#_c_567_p N_VGND_c_1268_n 0.00410965f $X=10.85 $Y=1.665 $X2=0
+ $Y2=0
cc_588 N_A_183_141#_c_574_p N_VGND_c_1268_n 0.0171054f $X=10.965 $Y=1.665 $X2=0
+ $Y2=0
cc_589 N_A_183_141#_c_401_n N_VGND_c_1268_n 0.041453f $X=11.355 $Y=1.665 $X2=0
+ $Y2=0
cc_590 N_A_183_141#_c_576_p N_VGND_c_1268_n 0.00590701f $X=12.41 $Y=1.665 $X2=0
+ $Y2=0
cc_591 N_A_183_141#_c_375_n N_VGND_c_1270_n 6.39245e-19 $X=11.585 $Y=1.565 $X2=0
+ $Y2=0
cc_592 N_A_183_141#_c_377_n N_VGND_c_1270_n 0.0473216f $X=12.365 $Y=1.565 $X2=0
+ $Y2=0
cc_593 N_A_183_141#_c_379_n N_VGND_c_1270_n 0.04751f $X=13.145 $Y=1.565 $X2=0
+ $Y2=0
cc_594 N_A_183_141#_c_381_n N_VGND_c_1270_n 6.39245e-19 $X=13.925 $Y=1.565 $X2=0
+ $Y2=0
cc_595 N_A_183_141#_c_389_n N_VGND_c_1270_n 7.87968e-19 $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_596 N_A_183_141#_c_576_p N_VGND_c_1270_n 0.00410965f $X=12.41 $Y=1.665 $X2=0
+ $Y2=0
cc_597 N_A_183_141#_c_583_p N_VGND_c_1270_n 0.0171054f $X=12.525 $Y=1.665 $X2=0
+ $Y2=0
cc_598 N_A_183_141#_c_403_n N_VGND_c_1270_n 0.041453f $X=12.915 $Y=1.665 $X2=0
+ $Y2=0
cc_599 N_A_183_141#_c_585_p N_VGND_c_1270_n 0.00590701f $X=13.97 $Y=1.665 $X2=0
+ $Y2=0
cc_600 N_A_183_141#_c_379_n N_VGND_c_1272_n 6.39245e-19 $X=13.145 $Y=1.565 $X2=0
+ $Y2=0
cc_601 N_A_183_141#_c_381_n N_VGND_c_1272_n 0.0473216f $X=13.925 $Y=1.565 $X2=0
+ $Y2=0
cc_602 N_A_183_141#_c_383_n N_VGND_c_1272_n 0.04751f $X=14.705 $Y=1.565 $X2=0
+ $Y2=0
cc_603 N_A_183_141#_c_385_n N_VGND_c_1272_n 6.39245e-19 $X=15.485 $Y=1.565 $X2=0
+ $Y2=0
cc_604 N_A_183_141#_c_389_n N_VGND_c_1272_n 7.87968e-19 $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_605 N_A_183_141#_c_585_p N_VGND_c_1272_n 0.00410965f $X=13.97 $Y=1.665 $X2=0
+ $Y2=0
cc_606 N_A_183_141#_c_592_p N_VGND_c_1272_n 0.0171054f $X=14.085 $Y=1.665 $X2=0
+ $Y2=0
cc_607 N_A_183_141#_c_405_n N_VGND_c_1272_n 0.041453f $X=14.475 $Y=1.665 $X2=0
+ $Y2=0
cc_608 N_A_183_141#_c_594_p N_VGND_c_1272_n 0.00590701f $X=15.53 $Y=1.665 $X2=0
+ $Y2=0
cc_609 N_A_183_141#_c_383_n N_VGND_c_1274_n 6.39245e-19 $X=14.705 $Y=1.565 $X2=0
+ $Y2=0
cc_610 N_A_183_141#_c_385_n N_VGND_c_1274_n 0.0473216f $X=15.485 $Y=1.565 $X2=0
+ $Y2=0
cc_611 N_A_183_141#_c_387_n N_VGND_c_1274_n 0.050102f $X=16.265 $Y=1.565 $X2=0
+ $Y2=0
cc_612 N_A_183_141#_c_389_n N_VGND_c_1274_n 0.00188124f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_613 N_A_183_141#_c_594_p N_VGND_c_1274_n 0.00410965f $X=15.53 $Y=1.665 $X2=0
+ $Y2=0
cc_614 N_A_183_141#_c_601_p N_VGND_c_1274_n 0.0171054f $X=15.645 $Y=1.665 $X2=0
+ $Y2=0
cc_615 N_A_183_141#_c_406_n N_VGND_c_1274_n 0.00281117f $X=16.035 $Y=1.665 $X2=0
+ $Y2=0
cc_616 N_A_183_141#_c_407_n N_VGND_c_1274_n 0.041453f $X=16.035 $Y=1.665 $X2=0
+ $Y2=0
cc_617 N_A_183_141#_c_387_n N_VGND_c_1276_n 0.00109203f $X=16.265 $Y=1.565 $X2=0
+ $Y2=0
cc_618 N_A_183_141#_c_389_n N_VGND_c_1276_n 0.0488451f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_619 N_A_183_141#_c_359_n N_VGND_c_1278_n 0.0145374f $X=5.345 $Y=1.565 $X2=0
+ $Y2=0
cc_620 N_A_183_141#_c_361_n N_VGND_c_1278_n 0.0109642f $X=6.125 $Y=1.565 $X2=0
+ $Y2=0
cc_621 N_A_183_141#_c_363_n N_VGND_c_1278_n 0.0109642f $X=6.905 $Y=1.565 $X2=0
+ $Y2=0
cc_622 N_A_183_141#_c_365_n N_VGND_c_1278_n 0.0109642f $X=7.685 $Y=1.565 $X2=0
+ $Y2=0
cc_623 N_A_183_141#_c_367_n N_VGND_c_1278_n 0.0109642f $X=8.465 $Y=1.565 $X2=0
+ $Y2=0
cc_624 N_A_183_141#_c_369_n N_VGND_c_1278_n 0.0109642f $X=9.245 $Y=1.565 $X2=0
+ $Y2=0
cc_625 N_A_183_141#_c_371_n N_VGND_c_1278_n 0.0109642f $X=10.025 $Y=1.565 $X2=0
+ $Y2=0
cc_626 N_A_183_141#_c_373_n N_VGND_c_1278_n 0.0109642f $X=10.805 $Y=1.565 $X2=0
+ $Y2=0
cc_627 N_A_183_141#_c_375_n N_VGND_c_1278_n 0.0109642f $X=11.585 $Y=1.565 $X2=0
+ $Y2=0
cc_628 N_A_183_141#_c_377_n N_VGND_c_1278_n 0.0109642f $X=12.365 $Y=1.565 $X2=0
+ $Y2=0
cc_629 N_A_183_141#_c_379_n N_VGND_c_1278_n 0.0109642f $X=13.145 $Y=1.565 $X2=0
+ $Y2=0
cc_630 N_A_183_141#_c_381_n N_VGND_c_1278_n 0.0109642f $X=13.925 $Y=1.565 $X2=0
+ $Y2=0
cc_631 N_A_183_141#_c_383_n N_VGND_c_1278_n 0.0109642f $X=14.705 $Y=1.565 $X2=0
+ $Y2=0
cc_632 N_A_183_141#_c_385_n N_VGND_c_1278_n 0.0109642f $X=15.485 $Y=1.565 $X2=0
+ $Y2=0
cc_633 N_A_183_141#_c_387_n N_VGND_c_1278_n 0.0109642f $X=16.265 $Y=1.565 $X2=0
+ $Y2=0
cc_634 N_A_183_141#_c_389_n N_VGND_c_1278_n 0.0129321f $X=17.045 $Y=1.565 $X2=0
+ $Y2=0
cc_635 N_A_183_141#_c_391_n N_VGND_c_1278_n 0.0140143f $X=1.055 $Y=0.92 $X2=0
+ $Y2=0
cc_636 N_A_183_141#_c_479_n N_VGND_c_1278_n 0.0124959f $X=2.4 $Y=1.302 $X2=0
+ $Y2=0
cc_637 N_A_183_141#_c_392_n N_VGND_c_1278_n 0.0157921f $X=2.615 $Y=0.895 $X2=0
+ $Y2=0
cc_638 N_A_183_141#_c_494_n N_VGND_c_1278_n 0.0123648f $X=4.025 $Y=1.302 $X2=0
+ $Y2=0
cc_639 N_A_183_141#_c_393_n N_VGND_c_1278_n 0.0102287f $X=4.175 $Y=0.895 $X2=0
+ $Y2=0
cc_640 N_A_183_141#_c_502_n N_VGND_c_1278_n 0.00874732f $X=4.8 $Y=1.302 $X2=0
+ $Y2=0
cc_641 N_VPWR_c_868_n X 4.51816e-19 $X=15.875 $Y=2.34 $X2=0 $Y2=0
cc_642 N_VPWR_c_871_n X 0.00134284f $X=17.435 $Y=2.36 $X2=0 $Y2=0
cc_643 N_VPWR_c_848_n N_X_c_1046_n 0.0753269f $X=4.955 $Y=2.55 $X2=0 $Y2=0
cc_644 N_VPWR_c_850_n N_X_c_1046_n 0.11835f $X=6.515 $Y=2.34 $X2=0 $Y2=0
cc_645 N_VPWR_c_874_n N_X_c_1046_n 0.0397803f $X=17.515 $Y=3.56 $X2=0 $Y2=0
cc_646 N_VPWR_c_850_n N_X_c_1049_n 0.11835f $X=6.515 $Y=2.34 $X2=0 $Y2=0
cc_647 N_VPWR_c_853_n N_X_c_1049_n 0.11835f $X=8.075 $Y=2.34 $X2=0 $Y2=0
cc_648 N_VPWR_c_874_n N_X_c_1049_n 0.037804f $X=17.515 $Y=3.56 $X2=0 $Y2=0
cc_649 N_VPWR_c_853_n N_X_c_1052_n 0.11835f $X=8.075 $Y=2.34 $X2=0 $Y2=0
cc_650 N_VPWR_c_856_n N_X_c_1052_n 0.11835f $X=9.635 $Y=2.34 $X2=0 $Y2=0
cc_651 N_VPWR_c_874_n N_X_c_1052_n 0.037804f $X=17.515 $Y=3.56 $X2=0 $Y2=0
cc_652 N_VPWR_c_856_n N_X_c_1055_n 0.11835f $X=9.635 $Y=2.34 $X2=0 $Y2=0
cc_653 N_VPWR_c_859_n N_X_c_1055_n 0.11835f $X=11.195 $Y=2.34 $X2=0 $Y2=0
cc_654 N_VPWR_c_874_n N_X_c_1055_n 0.037804f $X=17.515 $Y=3.56 $X2=0 $Y2=0
cc_655 N_VPWR_c_859_n N_X_c_1058_n 0.11835f $X=11.195 $Y=2.34 $X2=0 $Y2=0
cc_656 N_VPWR_c_862_n N_X_c_1058_n 0.11835f $X=12.755 $Y=2.34 $X2=0 $Y2=0
cc_657 N_VPWR_c_874_n N_X_c_1058_n 0.037804f $X=17.515 $Y=3.56 $X2=0 $Y2=0
cc_658 N_VPWR_c_862_n N_X_c_1061_n 0.11835f $X=12.755 $Y=2.34 $X2=0 $Y2=0
cc_659 N_VPWR_c_865_n N_X_c_1061_n 0.11835f $X=14.315 $Y=2.34 $X2=0 $Y2=0
cc_660 N_VPWR_c_874_n N_X_c_1061_n 0.037804f $X=17.515 $Y=3.56 $X2=0 $Y2=0
cc_661 N_VPWR_c_865_n N_X_c_1064_n 0.11835f $X=14.315 $Y=2.34 $X2=0 $Y2=0
cc_662 N_VPWR_c_868_n N_X_c_1064_n 0.11835f $X=15.875 $Y=2.34 $X2=0 $Y2=0
cc_663 N_VPWR_c_874_n N_X_c_1064_n 0.037804f $X=17.515 $Y=3.56 $X2=0 $Y2=0
cc_664 N_VPWR_c_868_n N_X_c_1067_n 0.119772f $X=15.875 $Y=2.34 $X2=0 $Y2=0
cc_665 N_VPWR_c_871_n N_X_c_1067_n 0.119397f $X=17.435 $Y=2.36 $X2=0 $Y2=0
cc_666 N_VPWR_c_874_n N_X_c_1067_n 0.0456596f $X=17.515 $Y=3.56 $X2=0 $Y2=0
cc_667 N_VPWR_c_850_n N_X_c_1148_n 0.0903983f $X=6.515 $Y=2.34 $X2=0 $Y2=0
cc_668 N_VPWR_c_848_n N_X_c_1152_n 5.42233e-19 $X=4.955 $Y=2.55 $X2=0 $Y2=0
cc_669 N_VPWR_c_850_n N_X_c_1152_n 4.51816e-19 $X=6.515 $Y=2.34 $X2=0 $Y2=0
cc_670 N_VPWR_c_853_n N_X_c_1153_n 0.0903983f $X=8.075 $Y=2.34 $X2=0 $Y2=0
cc_671 N_VPWR_c_850_n N_X_c_1157_n 4.51816e-19 $X=6.515 $Y=2.34 $X2=0 $Y2=0
cc_672 N_VPWR_c_853_n N_X_c_1157_n 4.51816e-19 $X=8.075 $Y=2.34 $X2=0 $Y2=0
cc_673 N_VPWR_c_856_n N_X_c_1158_n 0.0903983f $X=9.635 $Y=2.34 $X2=0 $Y2=0
cc_674 N_VPWR_c_853_n N_X_c_1162_n 4.51816e-19 $X=8.075 $Y=2.34 $X2=0 $Y2=0
cc_675 N_VPWR_c_856_n N_X_c_1162_n 4.51816e-19 $X=9.635 $Y=2.34 $X2=0 $Y2=0
cc_676 N_VPWR_c_859_n N_X_c_1163_n 0.0903983f $X=11.195 $Y=2.34 $X2=0 $Y2=0
cc_677 N_VPWR_c_856_n N_X_c_1167_n 4.51816e-19 $X=9.635 $Y=2.34 $X2=0 $Y2=0
cc_678 N_VPWR_c_859_n N_X_c_1167_n 4.51816e-19 $X=11.195 $Y=2.34 $X2=0 $Y2=0
cc_679 N_VPWR_c_862_n N_X_c_1168_n 0.0903983f $X=12.755 $Y=2.34 $X2=0 $Y2=0
cc_680 N_VPWR_c_859_n N_X_c_1172_n 4.51816e-19 $X=11.195 $Y=2.34 $X2=0 $Y2=0
cc_681 N_VPWR_c_862_n N_X_c_1172_n 4.51816e-19 $X=12.755 $Y=2.34 $X2=0 $Y2=0
cc_682 N_VPWR_c_865_n N_X_c_1173_n 0.0903983f $X=14.315 $Y=2.34 $X2=0 $Y2=0
cc_683 N_VPWR_c_862_n N_X_c_1177_n 4.51816e-19 $X=12.755 $Y=2.34 $X2=0 $Y2=0
cc_684 N_VPWR_c_865_n N_X_c_1177_n 4.51816e-19 $X=14.315 $Y=2.34 $X2=0 $Y2=0
cc_685 N_VPWR_c_868_n N_X_c_1178_n 0.0903983f $X=15.875 $Y=2.34 $X2=0 $Y2=0
cc_686 N_VPWR_c_865_n N_X_c_1182_n 4.51816e-19 $X=14.315 $Y=2.34 $X2=0 $Y2=0
cc_687 N_VPWR_c_868_n N_X_c_1182_n 4.51816e-19 $X=15.875 $Y=2.34 $X2=0 $Y2=0
cc_688 N_VPWR_c_871_n N_VGND_c_1276_n 0.0166422f $X=17.435 $Y=2.36 $X2=0 $Y2=0
cc_689 N_X_c_1046_n N_VGND_c_1260_n 0.0141738f $X=5.735 $Y=0.955 $X2=0 $Y2=0
cc_690 N_X_c_1046_n N_VGND_c_1262_n 0.0480657f $X=5.735 $Y=0.955 $X2=0 $Y2=0
cc_691 N_X_c_1049_n N_VGND_c_1262_n 0.0480657f $X=7.295 $Y=0.955 $X2=0 $Y2=0
cc_692 N_X_c_1049_n N_VGND_c_1264_n 0.0480657f $X=7.295 $Y=0.955 $X2=0 $Y2=0
cc_693 N_X_c_1052_n N_VGND_c_1264_n 0.0480657f $X=8.855 $Y=0.955 $X2=0 $Y2=0
cc_694 N_X_c_1052_n N_VGND_c_1266_n 0.0480657f $X=8.855 $Y=0.955 $X2=0 $Y2=0
cc_695 N_X_c_1055_n N_VGND_c_1266_n 0.0480657f $X=10.415 $Y=0.955 $X2=0 $Y2=0
cc_696 N_X_c_1055_n N_VGND_c_1268_n 0.0480657f $X=10.415 $Y=0.955 $X2=0 $Y2=0
cc_697 N_X_c_1058_n N_VGND_c_1268_n 0.0480657f $X=11.975 $Y=0.955 $X2=0 $Y2=0
cc_698 N_X_c_1058_n N_VGND_c_1270_n 0.0480657f $X=11.975 $Y=0.955 $X2=0 $Y2=0
cc_699 N_X_c_1061_n N_VGND_c_1270_n 0.0480657f $X=13.535 $Y=0.955 $X2=0 $Y2=0
cc_700 N_X_c_1061_n N_VGND_c_1272_n 0.0480657f $X=13.535 $Y=0.955 $X2=0 $Y2=0
cc_701 N_X_c_1064_n N_VGND_c_1272_n 0.0480657f $X=15.095 $Y=0.955 $X2=0 $Y2=0
cc_702 N_X_c_1064_n N_VGND_c_1274_n 0.0480657f $X=15.095 $Y=0.955 $X2=0 $Y2=0
cc_703 N_X_c_1067_n N_VGND_c_1274_n 0.0488323f $X=16.655 $Y=0.955 $X2=0 $Y2=0
cc_704 N_X_c_1067_n N_VGND_c_1276_n 0.0557875f $X=16.655 $Y=0.955 $X2=0 $Y2=0
cc_705 N_X_c_1046_n N_VGND_c_1278_n 0.0184011f $X=5.735 $Y=0.955 $X2=0 $Y2=0
cc_706 N_X_c_1049_n N_VGND_c_1278_n 0.0184011f $X=7.295 $Y=0.955 $X2=0 $Y2=0
cc_707 N_X_c_1052_n N_VGND_c_1278_n 0.0184011f $X=8.855 $Y=0.955 $X2=0 $Y2=0
cc_708 N_X_c_1055_n N_VGND_c_1278_n 0.0184011f $X=10.415 $Y=0.955 $X2=0 $Y2=0
cc_709 N_X_c_1058_n N_VGND_c_1278_n 0.0184011f $X=11.975 $Y=0.955 $X2=0 $Y2=0
cc_710 N_X_c_1061_n N_VGND_c_1278_n 0.0184011f $X=13.535 $Y=0.955 $X2=0 $Y2=0
cc_711 N_X_c_1064_n N_VGND_c_1278_n 0.0184011f $X=15.095 $Y=0.955 $X2=0 $Y2=0
cc_712 N_X_c_1067_n N_VGND_c_1278_n 0.0223691f $X=16.655 $Y=0.955 $X2=0 $Y2=0
