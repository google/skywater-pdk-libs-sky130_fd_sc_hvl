* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__buf_2 A VGND VNB VPB VPWR X
M1000 a_129_279# A VPWR VPB phv w=750000u l=500000u
+  ad=2.1375e+11p pd=2.07e+06u as=1.01625e+12p ps=7.57e+06u
M1001 X a_129_279# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=4.2e+11p pd=3.56e+06u as=0p ps=0u
M1002 X a_129_279# VGND VNB nhv w=750000u l=500000u
+  ad=2.1e+11p pd=2.06e+06u as=5.178e+11p ps=4.57e+06u
M1003 VPWR a_129_279# X VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_129_279# A VGND VNB nhv w=420000u l=500000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 VGND a_129_279# X VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
