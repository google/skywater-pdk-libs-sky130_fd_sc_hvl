* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__and3_1 A B C VGND VNB VPB VPWR X
M1000 a_30_517# B VPWR VPB phv w=420000u l=500000u
+  ad=2.373e+11p pd=2.81e+06u as=5.913e+11p ps=5.19e+06u
M1001 X a_30_517# VGND VNB nhv w=750000u l=500000u
+  ad=1.9875e+11p pd=2.03e+06u as=3.0405e+11p ps=2.5e+06u
M1002 a_201_173# A a_30_517# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=1.302e+11p ps=1.46e+06u
M1003 a_343_173# B a_201_173# VNB nhv w=420000u l=500000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 VGND C a_343_173# VNB nhv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_30_517# VPWR VPB phv w=1.5e+06u l=500000u
+  ad=4.275e+11p pd=3.57e+06u as=0p ps=0u
M1006 VPWR C a_30_517# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_30_517# VPB phv w=420000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
.ends
