* File: sky130_fd_sc_hvl__inv_4.pxi.spice
* Created: Wed Sep  2 09:07:00 2020
* 
x_PM_SKY130_FD_SC_HVL__INV_4%VNB N_VNB_M1001_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__INV_4%VNB
x_PM_SKY130_FD_SC_HVL__INV_4%VPB N_VPB_M1000_b VPB N_VPB_c_29_p VPB
+ PM_SKY130_FD_SC_HVL__INV_4%VPB
x_PM_SKY130_FD_SC_HVL__INV_4%A N_A_M1001_g N_A_M1000_g N_A_M1003_g N_A_M1002_g
+ N_A_M1005_g N_A_M1004_g N_A_M1007_g N_A_M1006_g A A A A A A N_A_c_68_n
+ N_A_c_69_n PM_SKY130_FD_SC_HVL__INV_4%A
x_PM_SKY130_FD_SC_HVL__INV_4%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_M1006_d
+ VPWR N_VPWR_c_142_n N_VPWR_c_145_n N_VPWR_c_148_n N_VPWR_c_151_n
+ PM_SKY130_FD_SC_HVL__INV_4%VPWR
x_PM_SKY130_FD_SC_HVL__INV_4%Y N_Y_M1001_d N_Y_M1005_d N_Y_M1000_s N_Y_M1004_s
+ N_Y_c_177_n N_Y_c_185_n N_Y_c_179_n N_Y_c_180_n N_Y_c_188_n N_Y_c_208_n
+ N_Y_c_181_n N_Y_c_189_n N_Y_c_216_n N_Y_c_183_n Y Y
+ PM_SKY130_FD_SC_HVL__INV_4%Y
x_PM_SKY130_FD_SC_HVL__INV_4%VGND N_VGND_M1001_s N_VGND_M1003_s N_VGND_M1007_s
+ VGND N_VGND_c_247_n N_VGND_c_249_n N_VGND_c_251_n N_VGND_c_253_n
+ PM_SKY130_FD_SC_HVL__INV_4%VGND
cc_1 N_VNB_M1001_b N_A_M1001_g 0.0523828f $X=-0.33 $Y=-0.265 $X2=0.815 $Y2=0.91
cc_2 N_VNB_c_2_p N_A_M1001_g 0.00179668f $X=0.24 $Y=0 $X2=0.815 $Y2=0.91
cc_3 N_VNB_M1001_b N_A_M1003_g 0.0403708f $X=-0.33 $Y=-0.265 $X2=1.595 $Y2=0.91
cc_4 N_VNB_c_2_p N_A_M1003_g 5.86481e-19 $X=0.24 $Y=0 $X2=1.595 $Y2=0.91
cc_5 N_VNB_M1001_b N_A_M1005_g 0.0420403f $X=-0.33 $Y=-0.265 $X2=2.375 $Y2=0.91
cc_6 N_VNB_c_2_p N_A_M1005_g 9.58849e-19 $X=0.24 $Y=0 $X2=2.375 $Y2=0.91
cc_7 N_VNB_M1001_b N_A_M1007_g 0.0524448f $X=-0.33 $Y=-0.265 $X2=3.155 $Y2=0.91
cc_8 N_VNB_c_2_p N_A_M1007_g 0.00221559f $X=0.24 $Y=0 $X2=3.155 $Y2=0.91
cc_9 N_VNB_M1001_b N_A_c_68_n 0.0709068f $X=-0.33 $Y=-0.265 $X2=0.565 $Y2=1.75
cc_10 N_VNB_M1001_b N_A_c_69_n 0.166907f $X=-0.33 $Y=-0.265 $X2=3.155 $Y2=1.75
cc_11 N_VNB_M1001_b N_Y_c_177_n 0.00864253f $X=-0.33 $Y=-0.265 $X2=1.595
+ $Y2=2.965
cc_12 N_VNB_c_2_p N_Y_c_177_n 6.32535e-19 $X=0.24 $Y=0 $X2=1.595 $Y2=2.965
cc_13 N_VNB_M1001_b N_Y_c_179_n 0.00277761f $X=-0.33 $Y=-0.265 $X2=2.375
+ $Y2=2.965
cc_14 N_VNB_M1001_b N_Y_c_180_n 0.00179631f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_15 N_VNB_M1001_b N_Y_c_181_n 0.0171253f $X=-0.33 $Y=-0.265 $X2=3.155
+ $Y2=2.085
cc_16 N_VNB_c_2_p N_Y_c_181_n 0.00201444f $X=0.24 $Y=0 $X2=3.155 $Y2=2.085
cc_17 N_VNB_M1001_b N_Y_c_183_n 0.00256618f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_18 N_VNB_M1001_b Y 0.0186833f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_19 N_VNB_M1001_b N_VGND_c_247_n 0.071716f $X=-0.33 $Y=-0.265 $X2=1.595
+ $Y2=2.085
cc_20 N_VNB_c_2_p N_VGND_c_247_n 0.00166879f $X=0.24 $Y=0 $X2=1.595 $Y2=2.085
cc_21 N_VNB_M1001_b N_VGND_c_249_n 0.0470168f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_22 N_VNB_c_2_p N_VGND_c_249_n 0.00269018f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_23 N_VNB_M1001_b N_VGND_c_251_n 0.0505015f $X=-0.33 $Y=-0.265 $X2=3.155
+ $Y2=2.085
cc_24 N_VNB_c_2_p N_VGND_c_251_n 9.30887e-19 $X=0.24 $Y=0 $X2=3.155 $Y2=2.085
cc_25 N_VNB_M1001_b N_VGND_c_253_n 0.0757686f $X=-0.33 $Y=-0.265 $X2=3.155
+ $Y2=2.965
cc_26 N_VNB_c_2_p N_VGND_c_253_n 0.410695f $X=0.24 $Y=0 $X2=3.155 $Y2=2.965
cc_27 N_VPB_M1000_b N_A_M1000_g 0.0407294f $X=-0.33 $Y=1.885 $X2=0.815 $Y2=2.965
cc_28 VPB N_A_M1000_g 0.00970178f $X=0 $Y=3.955 $X2=0.815 $Y2=2.965
cc_29 N_VPB_c_29_p N_A_M1000_g 0.0180287f $X=3.6 $Y=4.07 $X2=0.815 $Y2=2.965
cc_30 N_VPB_M1000_b N_A_M1002_g 0.0341668f $X=-0.33 $Y=1.885 $X2=1.595 $Y2=2.965
cc_31 VPB N_A_M1002_g 0.00970178f $X=0 $Y=3.955 $X2=1.595 $Y2=2.965
cc_32 N_VPB_c_29_p N_A_M1002_g 0.0158814f $X=3.6 $Y=4.07 $X2=1.595 $Y2=2.965
cc_33 N_VPB_M1000_b N_A_M1004_g 0.0346403f $X=-0.33 $Y=1.885 $X2=2.375 $Y2=2.965
cc_34 VPB N_A_M1004_g 0.00970178f $X=0 $Y=3.955 $X2=2.375 $Y2=2.965
cc_35 N_VPB_c_29_p N_A_M1004_g 0.0152133f $X=3.6 $Y=4.07 $X2=2.375 $Y2=2.965
cc_36 N_VPB_M1000_b N_A_M1006_g 0.0413942f $X=-0.33 $Y=1.885 $X2=3.155 $Y2=2.965
cc_37 VPB N_A_M1006_g 0.00970178f $X=0 $Y=3.955 $X2=3.155 $Y2=2.965
cc_38 N_VPB_c_29_p N_A_M1006_g 0.0160007f $X=3.6 $Y=4.07 $X2=3.155 $Y2=2.965
cc_39 N_VPB_M1000_b N_A_c_69_n 0.0856065f $X=-0.33 $Y=1.885 $X2=3.155 $Y2=1.75
cc_40 N_VPB_M1000_b N_VPWR_c_142_n 0.0731649f $X=-0.33 $Y=1.885 $X2=1.595
+ $Y2=2.085
cc_41 VPB N_VPWR_c_142_n 0.00199989f $X=0 $Y=3.955 $X2=1.595 $Y2=2.085
cc_42 N_VPB_c_29_p N_VPWR_c_142_n 0.0306202f $X=3.6 $Y=4.07 $X2=1.595 $Y2=2.085
cc_43 N_VPB_M1000_b N_VPWR_c_145_n 0.00125033f $X=-0.33 $Y=1.885 $X2=2.375
+ $Y2=2.085
cc_44 VPB N_VPWR_c_145_n 0.00406397f $X=0 $Y=3.955 $X2=2.375 $Y2=2.085
cc_45 N_VPB_c_29_p N_VPWR_c_145_n 0.047451f $X=3.6 $Y=4.07 $X2=2.375 $Y2=2.085
cc_46 N_VPB_M1000_b N_VPWR_c_148_n 0.0533552f $X=-0.33 $Y=1.885 $X2=3.155
+ $Y2=2.965
cc_47 VPB N_VPWR_c_148_n 0.00229469f $X=0 $Y=3.955 $X2=3.155 $Y2=2.965
cc_48 N_VPB_c_29_p N_VPWR_c_148_n 0.0299474f $X=3.6 $Y=4.07 $X2=3.155 $Y2=2.965
cc_49 N_VPB_M1000_b N_VPWR_c_151_n 0.0453415f $X=-0.33 $Y=1.885 $X2=1.595
+ $Y2=1.58
cc_50 VPB N_VPWR_c_151_n 0.407271f $X=0 $Y=3.955 $X2=1.595 $Y2=1.58
cc_51 N_VPB_c_29_p N_VPWR_c_151_n 0.0176808f $X=3.6 $Y=4.07 $X2=1.595 $Y2=1.58
cc_52 N_VPB_M1000_b N_Y_c_185_n 0.00125033f $X=-0.33 $Y=1.885 $X2=2.375 $Y2=0.91
cc_53 VPB N_Y_c_185_n 0.00108855f $X=0 $Y=3.955 $X2=2.375 $Y2=0.91
cc_54 N_VPB_c_29_p N_Y_c_185_n 0.0171423f $X=3.6 $Y=4.07 $X2=2.375 $Y2=0.91
cc_55 N_VPB_M1000_b N_Y_c_188_n 0.00447242f $X=-0.33 $Y=1.885 $X2=3.155
+ $Y2=1.415
cc_56 N_VPB_M1000_b N_Y_c_189_n 0.00228189f $X=-0.33 $Y=1.885 $X2=0.155 $Y2=1.58
cc_57 VPB N_Y_c_189_n 8.01732e-19 $X=0 $Y=3.955 $X2=0.155 $Y2=1.58
cc_58 N_VPB_c_29_p N_Y_c_189_n 0.0130099f $X=3.6 $Y=4.07 $X2=0.155 $Y2=1.58
cc_59 N_VPB_M1000_b Y 0.0129296f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_60 N_A_M1000_g N_VPWR_c_142_n 0.0546482f $X=0.815 $Y=2.965 $X2=0 $Y2=0
cc_61 N_A_M1002_g N_VPWR_c_142_n 6.45057e-19 $X=1.595 $Y=2.965 $X2=0 $Y2=0
cc_62 A N_VPWR_c_142_n 0.0220896f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_63 N_A_c_68_n N_VPWR_c_142_n 0.0114394f $X=0.565 $Y=1.75 $X2=0 $Y2=0
cc_64 N_A_M1000_g N_VPWR_c_145_n 5.07605e-19 $X=0.815 $Y=2.965 $X2=1.92 $Y2=0
cc_65 N_A_M1002_g N_VPWR_c_145_n 0.066565f $X=1.595 $Y=2.965 $X2=1.92 $Y2=0
cc_66 N_A_M1004_g N_VPWR_c_145_n 0.0712227f $X=2.375 $Y=2.965 $X2=1.92 $Y2=0
cc_67 N_A_M1006_g N_VPWR_c_145_n 6.22801e-19 $X=3.155 $Y=2.965 $X2=1.92 $Y2=0
cc_68 N_A_c_69_n N_VPWR_c_145_n 7.47936e-19 $X=3.155 $Y=1.75 $X2=1.92 $Y2=0
cc_69 N_A_M1006_g N_VPWR_c_148_n 0.0662647f $X=3.155 $Y=2.965 $X2=0 $Y2=0
cc_70 N_A_M1000_g N_VPWR_c_151_n 0.0213723f $X=0.815 $Y=2.965 $X2=0 $Y2=0
cc_71 N_A_M1002_g N_VPWR_c_151_n 0.0101061f $X=1.595 $Y=2.965 $X2=0 $Y2=0
cc_72 N_A_M1004_g N_VPWR_c_151_n 0.00778801f $X=2.375 $Y=2.965 $X2=0 $Y2=0
cc_73 N_A_M1006_g N_VPWR_c_151_n 0.0110007f $X=3.155 $Y=2.965 $X2=0 $Y2=0
cc_74 N_A_M1001_g N_Y_c_177_n 0.0176991f $X=0.815 $Y=0.91 $X2=0 $Y2=0
cc_75 N_A_M1003_g N_Y_c_177_n 9.97785e-19 $X=1.595 $Y=0.91 $X2=0 $Y2=0
cc_76 N_A_M1000_g N_Y_c_185_n 0.0412678f $X=0.815 $Y=2.965 $X2=0 $Y2=0
cc_77 N_A_M1002_g N_Y_c_185_n 0.033886f $X=1.595 $Y=2.965 $X2=0 $Y2=0
cc_78 N_A_M1003_g N_Y_c_179_n 0.0265845f $X=1.595 $Y=0.91 $X2=1.92 $Y2=0.057
cc_79 N_A_M1005_g N_Y_c_179_n 0.024675f $X=2.375 $Y=0.91 $X2=1.92 $Y2=0.057
cc_80 A N_Y_c_179_n 0.086013f $X=2.555 $Y=1.58 $X2=1.92 $Y2=0.057
cc_81 N_A_c_69_n N_Y_c_179_n 0.00313555f $X=3.155 $Y=1.75 $X2=1.92 $Y2=0.057
cc_82 N_A_M1001_g N_Y_c_180_n 0.00785763f $X=0.815 $Y=0.91 $X2=1.92 $Y2=0.058
cc_83 A N_Y_c_180_n 0.0192109f $X=2.555 $Y=1.58 $X2=1.92 $Y2=0.058
cc_84 N_A_c_69_n N_Y_c_180_n 0.00326295f $X=3.155 $Y=1.75 $X2=1.92 $Y2=0.058
cc_85 N_A_M1002_g N_Y_c_188_n 0.0128294f $X=1.595 $Y=2.965 $X2=1.92 $Y2=0.058
cc_86 N_A_M1004_g N_Y_c_188_n 0.0117526f $X=2.375 $Y=2.965 $X2=1.92 $Y2=0.058
cc_87 A N_Y_c_188_n 0.0847495f $X=2.555 $Y=1.58 $X2=1.92 $Y2=0.058
cc_88 N_A_c_69_n N_Y_c_188_n 0.0388162f $X=3.155 $Y=1.75 $X2=1.92 $Y2=0.058
cc_89 N_A_M1000_g N_Y_c_208_n 8.80685e-19 $X=0.815 $Y=2.965 $X2=0 $Y2=0
cc_90 N_A_M1002_g N_Y_c_208_n 2.00174e-19 $X=1.595 $Y=2.965 $X2=0 $Y2=0
cc_91 A N_Y_c_208_n 0.024005f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_92 N_A_c_69_n N_Y_c_208_n 0.0197872f $X=3.155 $Y=1.75 $X2=0 $Y2=0
cc_93 N_A_M1005_g N_Y_c_181_n 0.0194835f $X=2.375 $Y=0.91 $X2=0 $Y2=0
cc_94 N_A_M1007_g N_Y_c_181_n 0.0336881f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_95 N_A_M1004_g N_Y_c_189_n 0.00413112f $X=2.375 $Y=2.965 $X2=0 $Y2=0
cc_96 N_A_M1006_g N_Y_c_189_n 0.033388f $X=3.155 $Y=2.965 $X2=0 $Y2=0
cc_97 N_A_M1007_g N_Y_c_216_n 9.05608e-19 $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_98 N_A_c_69_n N_Y_c_216_n 0.013301f $X=3.155 $Y=1.75 $X2=0 $Y2=0
cc_99 N_A_M1005_g N_Y_c_183_n 0.00212994f $X=2.375 $Y=0.91 $X2=0 $Y2=0
cc_100 N_A_M1007_g N_Y_c_183_n 0.0134952f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_101 A N_Y_c_183_n 0.0180512f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A_c_69_n N_Y_c_183_n 0.00326295f $X=3.155 $Y=1.75 $X2=0 $Y2=0
cc_103 N_A_M1006_g Y 0.0145764f $X=3.155 $Y=2.965 $X2=0 $Y2=0
cc_104 A Y 0.0248818f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_105 N_A_c_69_n Y 0.0685439f $X=3.155 $Y=1.75 $X2=0 $Y2=0
cc_106 N_A_M1001_g N_VGND_c_247_n 0.0382519f $X=0.815 $Y=0.91 $X2=0 $Y2=0
cc_107 N_A_M1003_g N_VGND_c_247_n 7.71762e-19 $X=1.595 $Y=0.91 $X2=0 $Y2=0
cc_108 A N_VGND_c_247_n 0.0324963f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_109 N_A_c_68_n N_VGND_c_247_n 0.0137184f $X=0.565 $Y=1.75 $X2=0 $Y2=0
cc_110 N_A_M1001_g N_VGND_c_249_n 0.00104383f $X=0.815 $Y=0.91 $X2=0 $Y2=0
cc_111 N_A_M1003_g N_VGND_c_249_n 0.0426782f $X=1.595 $Y=0.91 $X2=0 $Y2=0
cc_112 N_A_M1005_g N_VGND_c_249_n 0.0385262f $X=2.375 $Y=0.91 $X2=0 $Y2=0
cc_113 N_A_M1007_g N_VGND_c_249_n 8.83219e-19 $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_114 N_A_M1007_g N_VGND_c_251_n 0.0221583f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_115 N_A_M1001_g N_VGND_c_253_n 0.0225077f $X=0.815 $Y=0.91 $X2=0 $Y2=0
cc_116 N_A_M1003_g N_VGND_c_253_n 0.00415827f $X=1.595 $Y=0.91 $X2=0 $Y2=0
cc_117 N_A_M1005_g N_VGND_c_253_n 0.00566915f $X=2.375 $Y=0.91 $X2=0 $Y2=0
cc_118 N_A_M1007_g N_VGND_c_253_n 0.0144441f $X=3.155 $Y=0.91 $X2=0 $Y2=0
cc_119 N_VPWR_c_151_n N_Y_M1004_s 0.00221032f $X=3.595 $Y=3.59 $X2=-0.33
+ $Y2=1.885
cc_120 N_VPWR_c_142_n N_Y_c_185_n 0.0628567f $X=0.425 $Y=2.34 $X2=0 $Y2=0
cc_121 N_VPWR_c_145_n N_Y_c_185_n 0.107449f $X=1.985 $Y=2.365 $X2=0 $Y2=0
cc_122 N_VPWR_c_151_n N_Y_c_185_n 0.0403613f $X=3.595 $Y=3.59 $X2=0 $Y2=0
cc_123 N_VPWR_c_145_n N_Y_c_188_n 0.0658156f $X=1.985 $Y=2.365 $X2=0 $Y2=0
cc_124 N_VPWR_c_145_n N_Y_c_189_n 0.0620876f $X=1.985 $Y=2.365 $X2=0 $Y2=0
cc_125 N_VPWR_c_148_n N_Y_c_189_n 0.0999238f $X=3.545 $Y=2.365 $X2=0 $Y2=0
cc_126 N_VPWR_c_151_n N_Y_c_189_n 0.0306945f $X=3.595 $Y=3.59 $X2=0 $Y2=0
cc_127 N_VPWR_c_148_n Y 0.046572f $X=3.545 $Y=2.365 $X2=0 $Y2=0
cc_128 N_Y_c_179_n N_VGND_M1003_s 0.00178343f $X=2.6 $Y=1.315 $X2=0 $Y2=0
cc_129 N_Y_c_177_n N_VGND_c_247_n 0.0289319f $X=1.205 $Y=0.66 $X2=0 $Y2=0
cc_130 N_Y_c_180_n N_VGND_c_247_n 0.00432383f $X=1.29 $Y=1.315 $X2=0 $Y2=0
cc_131 N_Y_c_177_n N_VGND_c_249_n 0.0238737f $X=1.205 $Y=0.66 $X2=0 $Y2=0
cc_132 N_Y_c_179_n N_VGND_c_249_n 0.0600374f $X=2.6 $Y=1.315 $X2=0 $Y2=0
cc_133 N_Y_c_181_n N_VGND_c_249_n 0.0416488f $X=2.765 $Y=0.66 $X2=0 $Y2=0
cc_134 N_Y_c_181_n N_VGND_c_251_n 0.0498041f $X=2.765 $Y=0.66 $X2=0 $Y2=0
cc_135 N_Y_c_183_n N_VGND_c_251_n 0.00679007f $X=2.892 $Y=1.315 $X2=0 $Y2=0
cc_136 Y N_VGND_c_251_n 0.0245923f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_137 N_Y_M1001_d N_VGND_c_253_n 7.65036e-19 $X=1.065 $Y=0.535 $X2=0 $Y2=0
cc_138 N_Y_c_177_n N_VGND_c_253_n 0.0252438f $X=1.205 $Y=0.66 $X2=0 $Y2=0
cc_139 N_Y_c_179_n N_VGND_c_253_n 0.0126589f $X=2.6 $Y=1.315 $X2=0 $Y2=0
cc_140 N_Y_c_181_n N_VGND_c_253_n 0.0534736f $X=2.765 $Y=0.66 $X2=0 $Y2=0
