* File: sky130_fd_sc_hvl__lsbufhv2lv_simple_1.spice
* Created: Fri Aug 28 09:36:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__lsbufhv2lv_simple_1.pex.spice"
.subckt sky130_fd_sc_hvl__lsbufhv2lv_simple_1  VNB VPB LVPWR A X VGND VPWR
* 
* VGND	VGND
* X	X
* A	A
* LVPWR	LVPWR
* VPB	VPB
* VNB	VNB
MM0_noxref N_VGND_M0_noxref_d N_A_662_81#_M0_noxref_g N_X_M0_noxref_s
+ N_VNB_M0_noxref_b NHV L=0.5 W=0.75 AD=0.194904 AS=0.19875 PD=1.60256 PS=2.03
+ NRD=0 NRS=0 M=1 R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1_noxref N_A_662_81#_M1_noxref_d N_A_M1_noxref_g N_VGND_M0_noxref_d
+ N_VNB_M0_noxref_b NHV L=0.5 W=0.42 AD=0.1197 AS=0.109146 PD=1.41 PS=0.897436
+ NRD=0 NRS=59.7132 M=1 R=0.84 SA=250001 SB=250000 A=0.21 P=1.84 MULT=1
MM1001 N_LVPWR_M1001_d N_A_662_81#_M1001_g N_X_M1001_s N_LVPWR_M1001_b PHV L=0.5
+ W=1.5 AD=0.34 AS=0.4275 PD=2.52667 PS=3.57 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
MM1003 N_A_662_81#_M1003_d N_A_M1003_g N_LVPWR_M1001_d N_LVPWR_M1001_b PHV L=0.5
+ W=0.75 AD=0.21375 AS=0.17 PD=2.07 PS=1.26333 NRD=0 NRS=29.2803 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
DX4_noxref N_VNB_M0_noxref_b N_VPB_X4_noxref_D1 NWDIODE A=4.9381 P=11
DX5_noxref N_VNB_M0_noxref_b N_LVPWR_M1001_b NWDIODE A=7.7175 P=11.13
DX6_noxref N_VNB_M0_noxref_b N_VPB_X6_noxref_D1 NWDIODE A=6.75165 P=11.83
*
.include "sky130_fd_sc_hvl__lsbufhv2lv_simple_1.pxi.spice"
*
.ends
*
*
