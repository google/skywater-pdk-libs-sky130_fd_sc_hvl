# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__nor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__nor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.775000 1.315000 2.120000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 1.775000 1.825000 2.120000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.637500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.200000 0.495000 1.530000 1.425000 ;
        RECT 1.200000 1.425000 2.275000 1.595000 ;
        RECT 2.020000 1.595000 2.275000 3.755000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 2.400000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 2.400000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 2.400000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 2.400000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 2.730000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 2.400000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.985000 2.400000 4.155000 ;
      RECT 0.090000  0.365000 1.020000 1.325000 ;
      RECT 0.090000  2.300000 1.760000 3.755000 ;
      RECT 1.720000  0.365000 2.310000 1.245000 ;
    LAYER mcon ;
      RECT 0.110000  0.395000 0.280000 0.565000 ;
      RECT 0.120000  3.505000 0.290000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.470000  0.395000 0.640000 0.565000 ;
      RECT 0.480000  3.505000 0.650000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.830000  0.395000 1.000000 0.565000 ;
      RECT 0.840000  3.505000 1.010000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.200000  3.505000 1.370000 3.675000 ;
      RECT 1.560000  3.505000 1.730000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.750000  0.395000 1.920000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.110000  0.395000 2.280000 0.565000 ;
  END
END sky130_fd_sc_hvl__nor2_1
END LIBRARY
