* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hvl__xor2_1 A B VGND VNB VPB VPWR X
M1000 a_531_443# a_30_443# X VPB phv w=1.5e+06u l=500000u
+  ad=8.475e+11p pd=7.13e+06u as=4.275e+11p ps=3.57e+06u
M1001 VPWR B a_531_443# VPB phv w=1.5e+06u l=500000u
+  ad=1.1925e+12p pd=7.59e+06u as=0p ps=0u
M1002 VGND a_30_443# X VNB nhv w=750000u l=500000u
+  ad=1.08e+12p pd=7.38e+06u as=2.1e+11p ps=2.06e+06u
M1003 a_617_107# A VGND VNB nhv w=750000u l=500000u
+  ad=1.575e+11p pd=1.92e+06u as=0p ps=0u
M1004 X B a_617_107# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_30_443# B VGND VNB nhv w=750000u l=500000u
+  ad=2.1e+11p pd=2.06e+06u as=0p ps=0u
M1006 a_531_443# A VPWR VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_187_443# VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=3.15e+11p ps=3.42e+06u
M1008 VGND A a_30_443# VNB nhv w=750000u l=500000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_187_443# B a_30_443# VPB phv w=1.5e+06u l=500000u
+  ad=0p pd=0u as=4.275e+11p ps=3.57e+06u
.ends
