* File: sky130_fd_sc_hvl__inv_2.pex.spice
* Created: Fri Aug 28 09:36:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__INV_2%VNB 5 7 11 25
r14 7 25 5.20833e-05 $w=2.4e-06 $l=1e-09 $layer=MET1_cond $X=1.2 $Y=0.057
+ $X2=1.2 $Y2=0.058
r15 7 11 0.00296875 $w=2.4e-06 $l=5.7e-08 $layer=MET1_cond $X=1.2 $Y=0.057
+ $X2=1.2 $Y2=0
r16 5 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r17 5 11 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_2%VPB 4 6 14 21
r19 10 21 0.00296875 $w=2.4e-06 $l=5.7e-08 $layer=MET1_cond $X=1.2 $Y=4.07
+ $X2=1.2 $Y2=4.013
r20 10 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=4.07
+ $X2=2.16 $Y2=4.07
r21 9 14 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=4.07
+ $X2=2.16 $Y2=4.07
r22 9 10 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r23 6 21 5.20833e-05 $w=2.4e-06 $l=1e-09 $layer=MET1_cond $X=1.2 $Y=4.012
+ $X2=1.2 $Y2=4.013
r24 4 14 72.8 $w=1.7e-07 $l=2.20209e-06 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=2.16 $Y2=4.07
r25 4 9 72.8 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=2 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_2%A 3 7 11 15 17 18 23 25
r40 24 25 65.8424 $w=5.71e-07 $l=7.8e-07 $layer=POLY_cond $X=0.935 $Y=1.772
+ $X2=1.715 $Y2=1.772
r41 22 24 2.5324 $w=5.71e-07 $l=3e-08 $layer=POLY_cond $X=0.905 $Y=1.772
+ $X2=0.935 $Y2=1.772
r42 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.905
+ $Y=1.715 $X2=0.905 $Y2=1.715
r43 18 23 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.72 $Y=1.715
+ $X2=0.905 $Y2=1.715
r44 17 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.715
+ $X2=0.72 $Y2=1.715
r45 13 25 5.98163 $w=5e-07 $l=3.13e-07 $layer=POLY_cond $X=1.715 $Y=2.085
+ $X2=1.715 $Y2=1.772
r46 13 15 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.715 $Y=2.085
+ $X2=1.715 $Y2=2.965
r47 9 25 5.98163 $w=5e-07 $l=3.12e-07 $layer=POLY_cond $X=1.715 $Y=1.46
+ $X2=1.715 $Y2=1.772
r48 9 11 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.715 $Y=1.46 $X2=1.715
+ $Y2=0.955
r49 5 24 5.98163 $w=5e-07 $l=3.13e-07 $layer=POLY_cond $X=0.935 $Y=2.085
+ $X2=0.935 $Y2=1.772
r50 5 7 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.935 $Y=2.085 $X2=0.935
+ $Y2=2.965
r51 1 24 5.98163 $w=5e-07 $l=3.12e-07 $layer=POLY_cond $X=0.935 $Y=1.46
+ $X2=0.935 $Y2=1.772
r52 1 3 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.935 $Y=1.46 $X2=0.935
+ $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_2%VPWR 1 2 7 10 20 25
r21 23 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.155 $Y=3.59
+ $X2=2.155 $Y2=3.59
r22 20 23 25.3406 $w=5.88e-07 $l=1.25e-06 $layer=LI1_cond $X=1.975 $Y=2.34
+ $X2=1.975 $Y2=3.59
r23 14 17 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.225 $Y=3.63
+ $X2=0.945 $Y2=3.63
r24 13 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.945 $Y=3.59
+ $X2=0.945 $Y2=3.59
r25 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.225 $Y=3.59
+ $X2=0.225 $Y2=3.59
r26 10 13 16.0526 $w=9.48e-07 $l=1.25e-06 $layer=LI1_cond $X=0.585 $Y=2.34
+ $X2=0.585 $Y2=3.59
r27 7 25 0.36663 $w=3.7e-07 $l=9.55e-07 $layer=MET1_cond $X=1.2 $Y=3.63
+ $X2=2.155 $Y2=3.63
r28 7 17 0.0978959 $w=3.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.2 $Y=3.63
+ $X2=0.945 $Y2=3.63
r29 2 23 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.965
+ $Y=2.215 $X2=2.105 $Y2=3.59
r30 2 20 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.965
+ $Y=2.215 $X2=2.105 $Y2=2.34
r31 1 13 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.4
+ $Y=2.215 $X2=0.545 $Y2=3.59
r32 1 10 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.4
+ $Y=2.215 $X2=0.545 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_2%Y 1 2 9 13 14 15 26 32
r27 32 33 6.18884 $w=5.93e-07 $l=7.5e-08 $layer=LI1_cond $X=1.497 $Y=1.295
+ $X2=1.497 $Y2=1.37
r28 14 32 0.100511 $w=5.93e-07 $l=5e-09 $layer=LI1_cond $X=1.497 $Y=1.29
+ $X2=1.497 $Y2=1.295
r29 14 15 11.0234 $w=2.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.68 $Y=1.375
+ $X2=1.68 $Y2=1.595
r30 14 33 0.250531 $w=2.28e-07 $l=5e-09 $layer=LI1_cond $X=1.68 $Y=1.375
+ $X2=1.68 $Y2=1.37
r31 13 14 7.33729 $w=5.93e-07 $l=3.65e-07 $layer=LI1_cond $X=1.497 $Y=0.925
+ $X2=1.497 $Y2=1.29
r32 13 26 4.42247 $w=5.93e-07 $l=2.2e-07 $layer=LI1_cond $X=1.497 $Y=0.925
+ $X2=1.497 $Y2=0.705
r33 9 11 57.6222 $w=2.48e-07 $l=1.25e-06 $layer=LI1_cond $X=1.365 $Y=2.34
+ $X2=1.365 $Y2=3.59
r34 7 15 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.365 $Y=1.695
+ $X2=1.68 $Y2=1.695
r35 7 9 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=1.365 $Y=1.78
+ $X2=1.365 $Y2=2.34
r36 2 11 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.185
+ $Y=2.215 $X2=1.325 $Y2=3.59
r37 2 9 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.185
+ $Y=2.215 $X2=1.325 $Y2=2.34
r38 1 26 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.185
+ $Y=0.58 $X2=1.325 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_2%VGND 1 2 7 10 19 20
r17 19 23 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=2.145 $Y=0.48
+ $X2=2.145 $Y2=0.705
r18 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.095 $Y=0.48
+ $X2=2.095 $Y2=0.48
r19 11 14 0.276412 $w=3.7e-07 $l=7.2e-07 $layer=MET1_cond $X=0.195 $Y=0.44
+ $X2=0.915 $Y2=0.44
r20 10 16 2.95161 $w=9.28e-07 $l=2.25e-07 $layer=LI1_cond $X=0.555 $Y=0.48
+ $X2=0.555 $Y2=0.705
r21 10 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.915 $Y=0.48
+ $X2=0.915 $Y2=0.48
r22 10 11 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.195 $Y=0.48
+ $X2=0.195 $Y2=0.48
r23 7 20 0.343595 $w=3.7e-07 $l=8.95e-07 $layer=MET1_cond $X=1.2 $Y=0.44
+ $X2=2.095 $Y2=0.44
r24 7 14 0.109413 $w=3.7e-07 $l=2.85e-07 $layer=MET1_cond $X=1.2 $Y=0.44
+ $X2=0.915 $Y2=0.44
r25 2 23 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.965
+ $Y=0.58 $X2=2.105 $Y2=0.705
r26 1 16 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.4
+ $Y=0.58 $X2=0.545 $Y2=0.705
.ends

