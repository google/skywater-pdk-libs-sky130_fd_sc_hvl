* File: sky130_fd_sc_hvl__inv_4.pex.spice
* Created: Wed Sep  2 09:07:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__INV_4%VNB 5 7 11 25
r26 7 25 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=0.057
+ $X2=1.92 $Y2=0.058
r27 7 11 0.00185547 $w=3.84e-06 $l=5.7e-08 $layer=MET1_cond $X=1.92 $Y=0.057
+ $X2=1.92 $Y2=0
r28 5 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r29 5 11 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_4%VPB 4 6 14 21
r33 10 21 0.00185547 $w=3.84e-06 $l=5.7e-08 $layer=MET1_cond $X=1.92 $Y=4.07
+ $X2=1.92 $Y2=4.013
r34 10 14 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=4.07
+ $X2=3.6 $Y2=4.07
r35 9 14 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=4.07 $X2=3.6
+ $Y2=4.07
r36 9 10 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r37 6 21 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=4.012
+ $X2=1.92 $Y2=4.013
r38 4 14 45.5 $w=1.7e-07 $l=3.64225e-06 $layer=licon1_NTAP_notbjt $count=4 $X=0
+ $Y=3.985 $X2=3.6 $Y2=4.07
r39 4 9 45.5 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=4 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_4%A 3 7 11 15 19 23 27 31 33 34 35 36 37 38 51
+ 57
c82 19 0 7.78561e-20 $X=2.375 $Y=0.91
r83 55 57 38.7297 $w=6.7e-07 $l=4.85e-07 $layer=POLY_cond $X=2.67 $Y=1.75
+ $X2=3.155 $Y2=1.75
r84 53 55 23.5573 $w=6.7e-07 $l=2.95e-07 $layer=POLY_cond $X=2.375 $Y=1.75
+ $X2=2.67 $Y2=1.75
r85 52 53 62.287 $w=6.7e-07 $l=7.8e-07 $layer=POLY_cond $X=1.595 $Y=1.75
+ $X2=2.375 $Y2=1.75
r86 50 52 62.287 $w=6.7e-07 $l=7.8e-07 $layer=POLY_cond $X=0.815 $Y=1.75
+ $X2=1.595 $Y2=1.75
r87 50 51 25.5047 $w=6.7e-07 $l=2.5e-07 $layer=POLY_cond $X=0.815 $Y=1.75
+ $X2=0.565 $Y2=1.75
r88 47 51 33.6137 $w=4.55e-07 $l=2.75e-07 $layer=POLY_cond $X=0.29 $Y=1.642
+ $X2=0.565 $Y2=1.642
r89 38 55 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=2.67
+ $Y=1.665 $X2=2.67 $Y2=1.665
r90 37 38 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.64 $Y2=1.665
r91 36 37 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=2.16 $Y2=1.665
r92 35 36 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.665
+ $X2=1.68 $Y2=1.665
r93 34 35 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=1.2 $Y2=1.665
r94 33 34 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.72 $Y2=1.665
r95 33 47 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=0.29
+ $Y=1.665 $X2=0.29 $Y2=1.665
r96 29 57 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.155 $Y=2.085
+ $X2=3.155 $Y2=1.75
r97 29 31 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.155 $Y=2.085
+ $X2=3.155 $Y2=2.965
r98 25 57 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.155 $Y=1.415
+ $X2=3.155 $Y2=1.75
r99 25 27 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.155 $Y=1.415
+ $X2=3.155 $Y2=0.91
r100 21 53 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.375 $Y=2.085
+ $X2=2.375 $Y2=1.75
r101 21 23 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.375 $Y=2.085
+ $X2=2.375 $Y2=2.965
r102 17 53 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.375 $Y=1.415
+ $X2=2.375 $Y2=1.75
r103 17 19 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.375 $Y=1.415
+ $X2=2.375 $Y2=0.91
r104 13 52 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.595 $Y=2.085
+ $X2=1.595 $Y2=1.75
r105 13 15 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.595 $Y=2.085
+ $X2=1.595 $Y2=2.965
r106 9 52 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.595 $Y=1.415
+ $X2=1.595 $Y2=1.75
r107 9 11 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.595 $Y=1.415
+ $X2=1.595 $Y2=0.91
r108 5 50 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.815 $Y=2.085
+ $X2=0.815 $Y2=1.75
r109 5 7 94.1652 $w=5e-07 $l=8.8e-07 $layer=POLY_cond $X=0.815 $Y=2.085
+ $X2=0.815 $Y2=2.965
r110 1 50 9.69179 $w=5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.815 $Y=1.415
+ $X2=0.815 $Y2=1.75
r111 1 3 54.038 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.815 $Y=1.415
+ $X2=0.815 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_4%VPWR 1 2 3 10 13 21 31 36
r35 34 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.595 $Y=3.59
+ $X2=3.595 $Y2=3.59
r36 31 34 24.8338 $w=5.88e-07 $l=1.225e-06 $layer=LI1_cond $X=3.415 $Y=2.365
+ $X2=3.415 $Y2=3.59
r37 28 36 0.464526 $w=3.7e-07 $l=1.21e-06 $layer=MET1_cond $X=2.385 $Y=3.63
+ $X2=3.595 $Y2=3.63
r38 24 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.385 $Y=3.59
+ $X2=2.385 $Y2=3.59
r39 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.665 $Y=3.59
+ $X2=1.665 $Y2=3.59
r40 21 24 15.7316 $w=9.48e-07 $l=1.225e-06 $layer=LI1_cond $X=2.025 $Y=2.365
+ $X2=2.025 $Y2=3.59
r41 18 25 0.422296 $w=3.7e-07 $l=1.1e-06 $layer=MET1_cond $X=0.565 $Y=3.63
+ $X2=1.665 $Y2=3.63
r42 16 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.565 $Y=3.59
+ $X2=0.565 $Y2=3.59
r43 13 16 25.3406 $w=5.88e-07 $l=1.25e-06 $layer=LI1_cond $X=0.385 $Y=2.34
+ $X2=0.385 $Y2=3.59
r44 10 28 0.178516 $w=3.7e-07 $l=4.65e-07 $layer=MET1_cond $X=1.92 $Y=3.63
+ $X2=2.385 $Y2=3.63
r45 10 25 0.0978959 $w=3.7e-07 $l=2.55e-07 $layer=MET1_cond $X=1.92 $Y=3.63
+ $X2=1.665 $Y2=3.63
r46 3 34 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=2.215 $X2=3.545 $Y2=3.59
r47 3 31 300 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=2.215 $X2=3.545 $Y2=2.365
r48 2 24 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.845
+ $Y=2.215 $X2=1.985 $Y2=3.59
r49 2 21 300 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=2 $X=1.845
+ $Y=2.215 $X2=1.985 $Y2=2.365
r50 1 16 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=0.28
+ $Y=2.215 $X2=0.425 $Y2=3.59
r51 1 13 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.28
+ $Y=2.215 $X2=0.425 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_4%Y 1 2 3 4 15 19 23 24 25 26 29 33 38 39 40 41
c70 38 0 7.78561e-20 $X=3.1 $Y=1.55
r71 40 41 13.7143 $w=4.27e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.825
+ $X2=3.6 $Y2=1.825
r72 40 45 0.571429 $w=4.27e-07 $l=2e-08 $layer=LI1_cond $X=3.12 $Y=1.825 $X2=3.1
+ $Y2=1.825
r73 38 45 6.17726 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.1 $Y=1.55 $X2=3.1
+ $Y2=1.825
r74 37 39 2.55177 $w=3.77e-07 $l=2.46868e-07 $layer=LI1_cond $X=3.1 $Y=1.4
+ $X2=2.892 $Y2=1.315
r75 37 38 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.1 $Y=1.4 $X2=3.1
+ $Y2=1.55
r76 33 35 57.6222 $w=2.48e-07 $l=1.25e-06 $layer=LI1_cond $X=2.805 $Y=2.34
+ $X2=2.805 $Y2=3.59
r77 31 45 8.42857 $w=4.27e-07 $l=4.10061e-07 $layer=LI1_cond $X=2.805 $Y=2.1
+ $X2=3.1 $Y2=1.825
r78 31 33 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=2.805 $Y=2.1
+ $X2=2.805 $Y2=2.34
r79 27 39 2.55177 $w=3.77e-07 $l=8.5e-08 $layer=LI1_cond $X=2.892 $Y=1.23
+ $X2=2.892 $Y2=1.315
r80 27 29 11.6541 $w=5.83e-07 $l=5.7e-07 $layer=LI1_cond $X=2.892 $Y=1.23
+ $X2=2.892 $Y2=0.66
r81 25 31 8.14142 $w=4.27e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.68 $Y=2.015
+ $X2=2.805 $Y2=2.1
r82 25 26 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=2.68 $Y=2.015
+ $X2=1.37 $Y2=2.015
r83 23 39 4.32201 $w=1.7e-07 $l=2.92e-07 $layer=LI1_cond $X=2.6 $Y=1.315
+ $X2=2.892 $Y2=1.315
r84 23 24 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=2.6 $Y=1.315
+ $X2=1.29 $Y2=1.315
r85 19 21 43.6531 $w=3.28e-07 $l=1.25e-06 $layer=LI1_cond $X=1.205 $Y=2.34
+ $X2=1.205 $Y2=3.59
r86 17 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.205 $Y=2.1
+ $X2=1.37 $Y2=2.015
r87 17 19 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.205 $Y=2.1
+ $X2=1.205 $Y2=2.34
r88 13 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.165 $Y=1.23
+ $X2=1.29 $Y2=1.315
r89 13 15 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=1.165 $Y=1.23
+ $X2=1.165 $Y2=0.66
r90 4 35 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=2.625
+ $Y=2.215 $X2=2.765 $Y2=3.59
r91 4 33 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.625
+ $Y=2.215 $X2=2.765 $Y2=2.34
r92 3 21 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=1.065
+ $Y=2.215 $X2=1.205 $Y2=3.59
r93 3 19 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.065
+ $Y=2.215 $X2=1.205 $Y2=2.34
r94 2 29 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.625
+ $Y=0.535 $X2=2.765 $Y2=0.66
r95 1 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.535 $X2=1.205 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HVL__INV_4%VGND 1 2 3 10 13 20 29 30
r34 29 33 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.545 $Y=0.48
+ $X2=3.545 $Y2=0.66
r35 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.495 $Y=0.48
+ $X2=3.495 $Y2=0.48
r36 24 30 0.456847 $w=3.7e-07 $l=1.19e-06 $layer=MET1_cond $X=2.305 $Y=0.44
+ $X2=3.495 $Y2=0.44
r37 20 26 4.23789 $w=9.48e-07 $l=3.3e-07 $layer=LI1_cond $X=1.945 $Y=0.48
+ $X2=1.945 $Y2=0.81
r38 20 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.305 $Y=0.48
+ $X2=2.305 $Y2=0.48
r39 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.585 $Y=0.48
+ $X2=1.585 $Y2=0.48
r40 14 21 0.391584 $w=3.7e-07 $l=1.02e-06 $layer=MET1_cond $X=0.565 $Y=0.44
+ $X2=1.585 $Y2=0.44
r41 13 17 3.64905 $w=5.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.385 $Y=0.48
+ $X2=0.385 $Y2=0.66
r42 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.565 $Y=0.48
+ $X2=0.565 $Y2=0.48
r43 10 24 0.147804 $w=3.7e-07 $l=3.85e-07 $layer=MET1_cond $X=1.92 $Y=0.44
+ $X2=2.305 $Y2=0.44
r44 10 21 0.128608 $w=3.7e-07 $l=3.35e-07 $layer=MET1_cond $X=1.92 $Y=0.44
+ $X2=1.585 $Y2=0.44
r45 3 33 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.535 $X2=3.545 $Y2=0.66
r46 2 26 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.535 $X2=1.985 $Y2=0.81
r47 1 17 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.28
+ $Y=0.535 $X2=0.425 $Y2=0.66
.ends

