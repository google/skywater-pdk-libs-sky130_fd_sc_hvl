* File: sky130_fd_sc_hvl__or2_1.pxi.spice
* Created: Fri Aug 28 09:39:02 2020
* 
x_PM_SKY130_FD_SC_HVL__OR2_1%VNB N_VNB_M1005_b VNB N_VNB_c_2_p VNB
+ PM_SKY130_FD_SC_HVL__OR2_1%VNB
x_PM_SKY130_FD_SC_HVL__OR2_1%VPB N_VPB_M1001_b VPB N_VPB_c_32_p VPB
+ PM_SKY130_FD_SC_HVL__OR2_1%VPB
x_PM_SKY130_FD_SC_HVL__OR2_1%B N_B_M1005_g N_B_M1001_g B N_B_c_45_n
+ PM_SKY130_FD_SC_HVL__OR2_1%B
x_PM_SKY130_FD_SC_HVL__OR2_1%A N_A_M1002_g N_A_M1003_g A N_A_c_73_n
+ PM_SKY130_FD_SC_HVL__OR2_1%A
x_PM_SKY130_FD_SC_HVL__OR2_1%A_84_443# N_A_84_443#_M1005_d N_A_84_443#_M1001_s
+ N_A_84_443#_c_105_n N_A_84_443#_c_106_n N_A_84_443#_c_107_n N_A_84_443#_c_99_n
+ N_A_84_443#_c_101_n N_A_84_443#_c_108_n N_A_84_443#_c_102_n
+ N_A_84_443#_c_109_n N_A_84_443#_c_135_n N_A_84_443#_M1004_g
+ N_A_84_443#_M1000_g PM_SKY130_FD_SC_HVL__OR2_1%A_84_443#
x_PM_SKY130_FD_SC_HVL__OR2_1%VPWR N_VPWR_M1002_d VPWR N_VPWR_c_157_n
+ N_VPWR_c_160_n PM_SKY130_FD_SC_HVL__OR2_1%VPWR
x_PM_SKY130_FD_SC_HVL__OR2_1%X N_X_M1004_d N_X_M1000_d X X X X X X X N_X_c_176_n
+ PM_SKY130_FD_SC_HVL__OR2_1%X
x_PM_SKY130_FD_SC_HVL__OR2_1%VGND N_VGND_M1005_s N_VGND_M1003_d VGND
+ N_VGND_c_189_n N_VGND_c_191_n N_VGND_c_193_n PM_SKY130_FD_SC_HVL__OR2_1%VGND
cc_1 N_VNB_M1005_b N_B_M1005_g 0.0480878f $X=-0.33 $Y=-0.265 $X2=0.955 $Y2=0.745
cc_2 N_VNB_c_2_p N_B_M1005_g 9.58849e-19 $X=0.24 $Y=0 $X2=0.955 $Y2=0.745
cc_3 N_VNB_M1005_b N_B_M1001_g 0.00920168f $X=-0.33 $Y=-0.265 $X2=0.955
+ $Y2=2.425
cc_4 N_VNB_M1005_b N_B_c_45_n 0.0999422f $X=-0.33 $Y=-0.265 $X2=0.77 $Y2=1.28
cc_5 N_VNB_M1005_b N_A_M1002_g 0.0076917f $X=-0.33 $Y=-0.265 $X2=0.955 $Y2=0.745
cc_6 N_VNB_M1005_b N_A_M1003_g 0.0517762f $X=-0.33 $Y=-0.265 $X2=0.955 $Y2=2.425
cc_7 N_VNB_c_2_p N_A_M1003_g 0.0023273f $X=0.24 $Y=0 $X2=0.955 $Y2=2.425
cc_8 N_VNB_M1005_b N_A_c_73_n 0.0774524f $X=-0.33 $Y=-0.265 $X2=0.77 $Y2=1.28
cc_9 N_VNB_M1005_b N_A_84_443#_c_99_n 0.0109585f $X=-0.33 $Y=-0.265 $X2=0.895
+ $Y2=1.805
cc_10 N_VNB_c_2_p N_A_84_443#_c_99_n 8.6949e-19 $X=0.24 $Y=0 $X2=0.895 $Y2=1.805
cc_11 N_VNB_M1005_b N_A_84_443#_c_101_n 0.00635686f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_12 N_VNB_M1005_b N_A_84_443#_c_102_n 0.00328414f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_13 N_VNB_M1005_b N_A_84_443#_M1004_g 0.0988747f $X=-0.33 $Y=-0.265 $X2=0
+ $Y2=0
cc_14 N_VNB_c_2_p N_A_84_443#_M1004_g 0.00137776f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_15 N_VNB_M1005_b N_X_c_176_n 0.068038f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_16 N_VNB_c_2_p N_X_c_176_n 5.92913e-19 $X=0.24 $Y=0 $X2=0 $Y2=0
cc_17 N_VNB_M1005_b N_VGND_c_189_n 0.0921789f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_18 N_VNB_c_2_p N_VGND_c_189_n 0.00258007f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_19 N_VNB_M1005_b N_VGND_c_191_n 0.0431647f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_20 N_VNB_c_2_p N_VGND_c_191_n 0.00166879f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_21 N_VNB_M1005_b N_VGND_c_193_n 0.0708262f $X=-0.33 $Y=-0.265 $X2=0 $Y2=0
cc_22 N_VNB_c_2_p N_VGND_c_193_n 0.359393f $X=0.24 $Y=0 $X2=0 $Y2=0
cc_23 N_VPB_M1001_b N_B_M1001_g 0.0626493f $X=-0.33 $Y=1.885 $X2=0.955 $Y2=2.425
cc_24 N_VPB_M1001_b N_A_M1002_g 0.054919f $X=-0.33 $Y=1.885 $X2=0.955 $Y2=0.745
cc_25 N_VPB_M1001_b N_A_84_443#_c_105_n 0.0345221f $X=-0.33 $Y=1.885 $X2=0.635
+ $Y2=1.21
cc_26 N_VPB_M1001_b N_A_84_443#_c_106_n 0.00217592f $X=-0.33 $Y=1.885 $X2=0.895
+ $Y2=1.28
cc_27 N_VPB_M1001_b N_A_84_443#_c_107_n 0.0157411f $X=-0.33 $Y=1.885 $X2=0.77
+ $Y2=1.28
cc_28 N_VPB_M1001_b N_A_84_443#_c_108_n 0.017055f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_29 N_VPB_M1001_b N_A_84_443#_c_109_n 0.00137622f $X=-0.33 $Y=1.885 $X2=0
+ $Y2=0
cc_30 N_VPB_M1001_b N_A_84_443#_M1004_g 0.062857f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_31 VPB N_A_84_443#_M1004_g 0.00970178f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_32 N_VPB_c_32_p N_A_84_443#_M1004_g 0.0152133f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_33 N_VPB_M1001_b N_VPWR_c_157_n 0.078714f $X=-0.33 $Y=1.885 $X2=0.955
+ $Y2=2.425
cc_34 VPB N_VPWR_c_157_n 0.00668042f $X=0 $Y=3.955 $X2=0.955 $Y2=2.425
cc_35 N_VPB_c_32_p N_VPWR_c_157_n 0.102514f $X=3.12 $Y=4.07 $X2=0.955 $Y2=2.425
cc_36 N_VPB_M1001_b N_VPWR_c_160_n 0.0844432f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_160_n 0.358324f $X=0 $Y=3.955 $X2=0 $Y2=0
cc_38 N_VPB_c_32_p N_VPWR_c_160_n 0.016558f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_39 N_VPB_M1001_b N_X_c_176_n 0.0688705f $X=-0.33 $Y=1.885 $X2=0 $Y2=0
cc_40 VPB N_X_c_176_n 7.75439e-19 $X=0 $Y=3.955 $X2=0 $Y2=0
cc_41 N_VPB_c_32_p N_X_c_176_n 0.0133691f $X=3.12 $Y=4.07 $X2=0 $Y2=0
cc_42 N_B_M1001_g N_A_M1002_g 0.0556707f $X=0.955 $Y=2.425 $X2=0 $Y2=0
cc_43 N_B_M1005_g N_A_M1003_g 0.0136537f $X=0.955 $Y=0.745 $X2=0 $Y2=0
cc_44 N_B_c_45_n A 4.38031e-19 $X=0.77 $Y=1.28 $X2=0 $Y2=0
cc_45 N_B_c_45_n N_A_c_73_n 0.0556707f $X=0.77 $Y=1.28 $X2=0 $Y2=0
cc_46 N_B_M1001_g N_A_84_443#_c_105_n 0.0083834f $X=0.955 $Y=2.425 $X2=0 $Y2=0
cc_47 N_B_M1001_g N_A_84_443#_c_106_n 0.0354123f $X=0.955 $Y=2.425 $X2=0.24
+ $Y2=0
cc_48 B N_A_84_443#_c_106_n 0.0204667f $X=0.635 $Y=1.21 $X2=0.24 $Y2=0
cc_49 N_B_c_45_n N_A_84_443#_c_106_n 0.00157739f $X=0.77 $Y=1.28 $X2=0.24 $Y2=0
cc_50 B N_A_84_443#_c_107_n 0.00369903f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_51 N_B_c_45_n N_A_84_443#_c_107_n 0.00240714f $X=0.77 $Y=1.28 $X2=0 $Y2=0
cc_52 N_B_M1005_g N_A_84_443#_c_99_n 0.00557052f $X=0.955 $Y=0.745 $X2=0 $Y2=0
cc_53 N_B_M1005_g N_A_84_443#_c_101_n 0.00449815f $X=0.955 $Y=0.745 $X2=0 $Y2=0
cc_54 N_B_M1001_g N_A_84_443#_c_101_n 0.00483648f $X=0.955 $Y=2.425 $X2=0 $Y2=0
cc_55 B N_A_84_443#_c_101_n 0.0293312f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_56 N_B_c_45_n N_A_84_443#_c_101_n 0.0219548f $X=0.77 $Y=1.28 $X2=0 $Y2=0
cc_57 N_B_M1005_g N_A_84_443#_c_102_n 0.00341076f $X=0.955 $Y=0.745 $X2=1.68
+ $Y2=0
cc_58 N_B_M1001_g N_A_84_443#_c_109_n 0.00230908f $X=0.955 $Y=2.425 $X2=0 $Y2=0
cc_59 N_B_M1001_g N_VPWR_c_157_n 0.0452934f $X=0.955 $Y=2.425 $X2=0 $Y2=0
cc_60 N_B_M1005_g N_VGND_c_189_n 0.0401989f $X=0.955 $Y=0.745 $X2=0.24 $Y2=0
cc_61 B N_VGND_c_189_n 0.025517f $X=0.635 $Y=1.21 $X2=0.24 $Y2=0
cc_62 N_B_c_45_n N_VGND_c_189_n 0.00406586f $X=0.77 $Y=1.28 $X2=0.24 $Y2=0
cc_63 N_B_M1005_g N_VGND_c_193_n 0.0109383f $X=0.955 $Y=0.745 $X2=0 $Y2=0
cc_64 B N_VGND_c_193_n 0.00117419f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A_M1003_g N_A_84_443#_c_99_n 0.00855706f $X=1.735 $Y=0.745 $X2=0 $Y2=0
cc_66 N_A_M1003_g N_A_84_443#_c_101_n 0.002022f $X=1.735 $Y=0.745 $X2=0 $Y2=0
cc_67 A N_A_84_443#_c_101_n 0.0395874f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A_c_73_n N_A_84_443#_c_101_n 0.0103306f $X=1.695 $Y=1.28 $X2=0 $Y2=0
cc_69 N_A_M1002_g N_A_84_443#_c_108_n 0.0317329f $X=1.665 $Y=2.425 $X2=0 $Y2=0
cc_70 A N_A_84_443#_c_108_n 0.0234404f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A_c_73_n N_A_84_443#_c_108_n 0.00313508f $X=1.695 $Y=1.28 $X2=0 $Y2=0
cc_72 N_A_M1003_g N_A_84_443#_c_102_n 0.00601582f $X=1.735 $Y=0.745 $X2=1.68
+ $Y2=0
cc_73 N_A_c_73_n N_A_84_443#_c_102_n 0.00354748f $X=1.695 $Y=1.28 $X2=1.68 $Y2=0
cc_74 N_A_M1002_g N_A_84_443#_c_135_n 7.03057e-19 $X=1.665 $Y=2.425 $X2=1.68
+ $Y2=0.058
cc_75 N_A_c_73_n N_A_84_443#_c_135_n 5.15092e-19 $X=1.695 $Y=1.28 $X2=1.68
+ $Y2=0.058
cc_76 N_A_M1002_g N_A_84_443#_M1004_g 0.0167588f $X=1.665 $Y=2.425 $X2=0 $Y2=0
cc_77 N_A_M1003_g N_A_84_443#_M1004_g 0.0308706f $X=1.735 $Y=0.745 $X2=0 $Y2=0
cc_78 A N_A_84_443#_M1004_g 0.00216669f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A_M1002_g N_VPWR_c_157_n 0.0579411f $X=1.665 $Y=2.425 $X2=0 $Y2=0
cc_80 N_A_M1003_g N_VGND_c_189_n 8.5578e-19 $X=1.735 $Y=0.745 $X2=0.24 $Y2=0
cc_81 N_A_M1003_g N_VGND_c_191_n 0.0151551f $X=1.735 $Y=0.745 $X2=0 $Y2=0
cc_82 A N_VGND_c_191_n 0.0119199f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A_M1003_g N_VGND_c_193_n 0.0228083f $X=1.735 $Y=0.745 $X2=0 $Y2=0
cc_84 A N_VGND_c_193_n 0.0103412f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A_84_443#_c_105_n N_VPWR_c_157_n 0.0183139f $X=0.565 $Y=2.425 $X2=0
+ $Y2=0
cc_86 N_A_84_443#_c_106_n N_VPWR_c_157_n 0.0253546f $X=1.18 $Y=1.99 $X2=0 $Y2=0
cc_87 N_A_84_443#_c_108_n N_VPWR_c_157_n 0.0759989f $X=2.445 $Y=1.99 $X2=0 $Y2=0
cc_88 N_A_84_443#_c_109_n N_VPWR_c_157_n 0.0122566f $X=1.265 $Y=1.99 $X2=0 $Y2=0
cc_89 N_A_84_443#_c_135_n N_VPWR_c_157_n 0.0252329f $X=2.61 $Y=1.89 $X2=0 $Y2=0
cc_90 N_A_84_443#_M1004_g N_VPWR_c_157_n 0.0755587f $X=2.675 $Y=0.91 $X2=0 $Y2=0
cc_91 N_A_84_443#_M1004_g N_VPWR_c_160_n 0.00915578f $X=2.675 $Y=0.91 $X2=3.12
+ $Y2=0
cc_92 N_A_84_443#_c_135_n N_X_c_176_n 0.0235826f $X=2.61 $Y=1.89 $X2=0 $Y2=0
cc_93 N_A_84_443#_M1004_g N_X_c_176_n 0.043741f $X=2.675 $Y=0.91 $X2=0 $Y2=0
cc_94 N_A_84_443#_c_99_n N_VGND_c_189_n 0.0360269f $X=1.345 $Y=0.745 $X2=0.24
+ $Y2=0
cc_95 N_A_84_443#_c_99_n N_VGND_c_191_n 0.00806507f $X=1.345 $Y=0.745 $X2=0
+ $Y2=0
cc_96 N_A_84_443#_c_108_n N_VGND_c_191_n 0.0143436f $X=2.445 $Y=1.99 $X2=0 $Y2=0
cc_97 N_A_84_443#_c_135_n N_VGND_c_191_n 0.00736155f $X=2.61 $Y=1.89 $X2=0 $Y2=0
cc_98 N_A_84_443#_M1004_g N_VGND_c_191_n 0.044738f $X=2.675 $Y=0.91 $X2=0 $Y2=0
cc_99 N_A_84_443#_c_99_n N_VGND_c_193_n 0.0299668f $X=1.345 $Y=0.745 $X2=0 $Y2=0
cc_100 N_A_84_443#_M1004_g N_VGND_c_193_n 0.0196534f $X=2.675 $Y=0.91 $X2=0
+ $Y2=0
cc_101 A_241_443# N_VPWR_c_157_n 0.00108862f $X=1.205 $Y=2.215 $X2=2.285
+ $Y2=2.34
cc_102 N_VPWR_c_160_n N_X_M1000_d 0.00221032f $X=2.715 $Y=3.59 $X2=0 $Y2=0
cc_103 N_VPWR_c_157_n N_X_c_176_n 0.0630924f $X=2.285 $Y=2.34 $X2=1.68 $Y2=4.07
cc_104 N_VPWR_c_160_n N_X_c_176_n 0.035852f $X=2.715 $Y=3.59 $X2=1.68 $Y2=4.07
cc_105 N_X_c_176_n N_VGND_c_191_n 0.0203006f $X=3.065 $Y=0.66 $X2=0 $Y2=0
cc_106 N_X_M1004_d N_VGND_c_193_n 0.00221032f $X=2.925 $Y=0.535 $X2=0 $Y2=0
cc_107 N_X_c_176_n N_VGND_c_193_n 0.0276948f $X=3.065 $Y=0.66 $X2=0 $Y2=0
