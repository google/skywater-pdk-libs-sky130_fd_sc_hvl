* File: sky130_fd_sc_hvl__sdfrbp_1.spice
* Created: Fri Aug 28 09:39:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__sdfrbp_1.pex.spice"
.subckt sky130_fd_sc_hvl__sdfrbp_1  VNB VPB SCE D SCD CLK RESET_B VPWR Q_N Q
+ VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1029 N_A_222_131#_M1029_d N_SCE_M1029_g N_VGND_M1029_s N_VNB_M1029_b NHV L=0.5
+ W=0.42 AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1040 noxref_26 N_D_M1040_g N_noxref_25_M1040_s N_VNB_M1029_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=13.566 NRS=0 M=1 R=0.84 SA=250000
+ SB=250004 A=0.21 P=1.84 MULT=1
MM1041 N_A_339_655#_M1041_d N_A_222_131#_M1041_g noxref_26 N_VNB_M1029_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250001 SB=250003 A=0.21 P=1.84 MULT=1
MM1031 noxref_27 N_SCE_M1031_g N_A_339_655#_M1041_d N_VNB_M1029_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1035 N_noxref_25_M1035_d N_SCD_M1035_g noxref_27 N_VNB_M1029_b NHV L=0.5
+ W=0.42 AD=0.090725 AS=0.0441 PD=0.895 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1007 N_VGND_M1007_d N_RESET_B_M1007_g N_noxref_25_M1035_d N_VNB_M1029_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.090725 PD=0.7 PS=0.895 NRD=0 NRS=28.4886 M=1
+ R=0.84 SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1026 N_A_1290_126#_M1026_d N_CLK_M1026_g N_VGND_M1007_d N_VNB_M1029_b NHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250003 SB=250000 A=0.21 P=1.84 MULT=1
MM1000 N_A_1569_126#_M1000_d N_A_1290_126#_M1000_g N_VGND_M1000_s N_VNB_M1029_b
+ NHV L=0.5 W=0.42 AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1027 N_A_1816_659#_M1027_d N_A_1290_126#_M1027_g N_A_339_655#_M1027_s
+ N_VNB_M1029_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250006 A=0.21 P=1.84 MULT=1
MM1004 A_1999_126# N_A_1569_126#_M1004_g N_A_1816_659#_M1027_d N_VNB_M1029_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250001 SB=250006 A=0.21 P=1.84 MULT=1
MM1005 A_2141_126# N_A_2014_537#_M1005_g A_1999_126# N_VNB_M1029_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=13.566 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1008 N_VGND_M1008_d N_RESET_B_M1008_g A_2141_126# N_VNB_M1029_b NHV L=0.5
+ W=0.42 AD=0.0971026 AS=0.0441 PD=0.84359 PS=0.63 NRD=24.4188 NRS=13.566 M=1
+ R=0.84 SA=250002 SB=250004 A=0.21 P=1.84 MULT=1
MM1039 N_A_2014_537#_M1039_d N_A_1816_659#_M1039_g N_VGND_M1008_d N_VNB_M1029_b
+ NHV L=0.5 W=0.75 AD=0.105 AS=0.173397 PD=1.03 PS=1.50641 NRD=0 NRS=9.1086 M=1
+ R=1.5 SA=250002 SB=250003 A=0.375 P=2.5 MULT=1
MM1028 N_A_2624_107#_M1028_d N_A_1569_126#_M1028_g N_A_2014_537#_M1039_d
+ N_VNB_M1029_b NHV L=0.5 W=0.75 AD=0.157019 AS=0.105 PD=1.44231 PS=1.03 NRD=0
+ NRS=0 M=1 R=1.5 SA=250003 SB=250002 A=0.375 P=2.5 MULT=1
MM1020 A_2799_107# N_A_1290_126#_M1020_g N_A_2624_107#_M1028_d N_VNB_M1029_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0879308 PD=0.63 PS=0.807692 NRD=13.566 NRS=25.7754
+ M=1 R=0.84 SA=250004 SB=250002 A=0.21 P=1.84 MULT=1
MM1030 N_VGND_M1030_d N_A_2841_81#_M1030_g A_2799_107# N_VNB_M1029_b NHV L=0.5
+ W=0.42 AD=0.05985 AS=0.0441 PD=0.705 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250005 SB=250002 A=0.21 P=1.84 MULT=1
MM1014 A_3098_107# N_RESET_B_M1014_g N_VGND_M1030_d N_VNB_M1029_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.05985 PD=0.63 PS=0.705 NRD=13.566 NRS=1.3566 M=1 R=0.84
+ SA=250006 SB=250001 A=0.21 P=1.84 MULT=1
MM1015 N_A_2841_81#_M1015_d N_A_2624_107#_M1015_g A_3098_107# N_VNB_M1029_b NHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250006 SB=250000 A=0.21 P=1.84 MULT=1
MM1023 N_Q_N_M1023_d N_A_2624_107#_M1023_g N_VGND_M1023_s N_VNB_M1029_b NHV
+ L=0.5 W=0.75 AD=0.19875 AS=0.19875 PD=2.03 PS=2.03 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1009 N_VGND_M1009_d N_A_2624_107#_M1009_g N_A_3613_443#_M1009_s N_VNB_M1029_b
+ NHV L=0.5 W=0.42 AD=0.0879308 AS=0.1113 PD=0.807692 PS=1.37 NRD=25.7754 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1010 N_Q_M1010_d N_A_3613_443#_M1010_g N_VGND_M1009_d N_VNB_M1029_b NHV L=0.5
+ W=0.75 AD=0.19875 AS=0.157019 PD=2.03 PS=1.44231 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1018 N_A_222_131#_M1018_d N_SCE_M1018_g N_VPWR_M1018_s N_VPB_M1018_b PHV L=0.5
+ W=0.42 AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1001 A_496_655# N_D_M1001_g N_A_339_655#_M1001_s N_VPB_M1018_b PHV L=0.5
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250000 SB=250004 A=0.21 P=1.84 MULT=1
MM1016 N_VPWR_M1016_d N_SCE_M1016_g A_496_655# N_VPB_M1018_b PHV L=0.5 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84 SA=250001
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1033 A_794_655# N_SCD_M1033_g N_VPWR_M1016_d N_VPB_M1018_b PHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84 SA=250002
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1006 N_A_339_655#_M1006_d N_A_222_131#_M1006_g A_794_655# N_VPB_M1018_b PHV
+ L=0.5 W=0.42 AD=0.0672 AS=0.0441 PD=0.74 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1012 N_VPWR_M1012_d N_RESET_B_M1012_g N_A_339_655#_M1006_d N_VPB_M1018_b PHV
+ L=0.5 W=0.42 AD=0.101608 AS=0.0672 PD=0.861538 PS=0.74 NRD=77.2977 NRS=18.1832
+ M=1 R=0.84 SA=250003 SB=250001 A=0.21 P=1.84 MULT=1
MM1002 N_A_1290_126#_M1002_d N_CLK_M1002_g N_VPWR_M1012_d N_VPB_M1018_b PHV
+ L=0.5 W=0.75 AD=0.21375 AS=0.181442 PD=2.07 PS=1.53846 NRD=0 NRS=0 M=1 R=1.5
+ SA=250002 SB=250000 A=0.375 P=2.5 MULT=1
MM1019 N_A_1569_126#_M1019_d N_A_1290_126#_M1019_g N_VPWR_M1019_s N_VPB_M1018_b
+ PHV L=0.5 W=0.75 AD=0.19875 AS=0.21375 PD=2.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1017 N_A_1816_659#_M1017_d N_A_1569_126#_M1017_g N_A_339_655#_M1017_s
+ N_VPB_M1018_b PHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1037 A_1972_659# N_A_1290_126#_M1037_g N_A_1816_659#_M1017_d N_VPB_M1018_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250001 SB=250002 A=0.21 P=1.84 MULT=1
MM1038 N_VPWR_M1038_d N_A_2014_537#_M1038_g A_1972_659# N_VPB_M1018_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1013 N_A_1816_659#_M1013_d N_RESET_B_M1013_g N_VPWR_M1038_d N_VPB_M1018_b PHV
+ L=0.5 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1003 N_A_2014_537#_M1003_d N_A_1816_659#_M1003_g N_VPWR_M1003_s N_VPB_M1018_b
+ PHV L=0.5 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=2 SA=250000
+ SB=250003 A=0.5 P=3 MULT=1
MM1024 N_A_2624_107#_M1024_d N_A_1290_126#_M1024_g N_A_2014_537#_M1003_d
+ N_VPB_M1018_b PHV L=0.5 W=1 AD=0.233239 AS=0.14 PD=1.96479 PS=1.28 NRD=0 NRS=0
+ M=1 R=2 SA=250001 SB=250002 A=0.5 P=3 MULT=1
MM1011 A_2871_543# N_A_1569_126#_M1011_g N_A_2624_107#_M1024_d N_VPB_M1018_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0979606 PD=0.63 PS=0.825211 NRD=22.729 NRS=52.2958
+ M=1 R=0.84 SA=250002 SB=250003 A=0.21 P=1.84 MULT=1
MM1025 N_VPWR_M1025_d N_A_2841_81#_M1025_g A_2871_543# N_VPB_M1018_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1034 N_A_2841_81#_M1034_d N_RESET_B_M1034_g N_VPWR_M1025_d N_VPB_M1018_b PHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=0.84
+ SA=250003 SB=250002 A=0.21 P=1.84 MULT=1
MM1021 N_VPWR_M1021_d N_A_2624_107#_M1021_g N_A_2841_81#_M1034_d N_VPB_M1018_b
+ PHV L=0.5 W=0.42 AD=0.0970594 AS=0.0588 PD=0.820312 PS=0.7 NRD=44.3311 NRS=0
+ M=1 R=0.84 SA=250004 SB=250001 A=0.21 P=1.84 MULT=1
MM1032 N_Q_N_M1032_d N_A_2624_107#_M1032_g N_VPWR_M1021_d N_VPB_M1018_b PHV
+ L=0.5 W=1.5 AD=0.3975 AS=0.346641 PD=3.53 PS=2.92969 NRD=0 NRS=0 M=1 R=3
+ SA=250001 SB=250000 A=0.75 P=4 MULT=1
MM1036 N_VPWR_M1036_d N_A_2624_107#_M1036_g N_A_3613_443#_M1036_s N_VPB_M1018_b
+ PHV L=0.5 W=0.75 AD=0.17 AS=0.19875 PD=1.26333 PS=2.03 NRD=29.2803 NRS=0 M=1
+ R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1022 N_Q_M1022_d N_A_3613_443#_M1022_g N_VPWR_M1036_d N_VPB_M1018_b PHV L=0.5
+ W=1.5 AD=0.4275 AS=0.34 PD=3.57 PS=2.52667 NRD=0 NRS=0 M=1 R=3 SA=250000
+ SB=250000 A=0.75 P=4 MULT=1
DX42_noxref N_VNB_M1029_b N_VPB_M1018_b NWDIODE A=54.4108 P=47.17
*
.include "sky130_fd_sc_hvl__sdfrbp_1.pxi.spice"
*
.ends
*
*
