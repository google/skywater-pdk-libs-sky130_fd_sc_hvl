* File: sky130_fd_sc_hvl__lsbufhv2lv_simple_1.pex.spice
* Created: Wed Sep  2 09:07:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%VNB 9 11 12 17 43
r25 12 29 0.00083912 $w=8.64e-06 $l=5.8e-08 $layer=MET1_cond $X=4.32 $Y=8.082
+ $X2=4.32 $Y2=8.14
r26 11 43 1.44676e-05 $w=8.64e-06 $l=1e-09 $layer=MET1_cond $X=4.32 $Y=0.057
+ $X2=4.32 $Y2=0.058
r27 11 17 0.000824653 $w=8.64e-06 $l=5.7e-08 $layer=MET1_cond $X=4.32 $Y=0.057
+ $X2=4.32 $Y2=0
r28 9 29 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=8.4 $Y=8.14
+ $X2=8.4 $Y2=8.14
r29 9 29 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=0.24 $Y=8.14
+ $X2=0.24 $Y2=8.14
r30 9 17 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r31 9 17 1.03333 $w=1.7e-07 $l=1.53e-06 $layer=mcon $count=9 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%VPB 7 8 11 14 20 21
r19 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=4.07 $X2=8.4
+ $Y2=4.07
r20 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=4.07
+ $X2=0.24 $Y2=4.07
r21 11 21 2.61775 $w=2.3e-07 $l=4.08e-06 $layer=MET1_cond $X=4.32 $Y=4.07
+ $X2=8.4 $Y2=4.07
r22 11 15 2.61775 $w=2.3e-07 $l=4.08e-06 $layer=MET1_cond $X=4.32 $Y=4.07
+ $X2=0.24 $Y2=4.07
r23 8 20 91 $w=1.7e-07 $l=6.86185e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=7.755 $Y=3.985 $X2=8.4 $Y2=4.07
r24 7 14 182 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_NTAP_notbjt $count=1 $X=0
+ $Y=3.985 $X2=0.24 $Y2=4.07
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%LVPWR 1 7 11 13 16 19
r35 22 25 9.26691 $w=5.53e-07 $l=4.3e-07 $layer=LI1_cond $X=3.897 $Y=3.16
+ $X2=3.897 $Y2=3.59
r36 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.075 $Y=3.16
+ $X2=4.075 $Y2=3.16
r37 19 22 17.6718 $w=5.53e-07 $l=8.2e-07 $layer=LI1_cond $X=3.897 $Y=2.34
+ $X2=3.897 $Y2=3.16
r38 16 23 0.122109 $w=2.85e-07 $l=2.45e-07 $layer=MET1_cond $X=4.32 $Y=3.162
+ $X2=4.075 $Y2=3.162
r39 13 25 7.8661 $w=5.53e-07 $l=3.65e-07 $layer=LI1_cond $X=3.897 $Y=3.955
+ $X2=3.897 $Y2=3.59
r40 13 15 3.4317 $w=5.55e-07 $l=3.88652e-07 $layer=LI1_cond $X=3.897 $Y=3.955
+ $X2=3.652 $Y2=4.24
r41 9 15 3.38637 $w=5.7e-07 $l=5.23e-07 $layer=LI1_cond $X=4.175 $Y=4.24
+ $X2=3.652 $Y2=4.24
r42 9 11 15.0034 $w=5.68e-07 $l=7.15e-07 $layer=LI1_cond $X=4.175 $Y=4.24
+ $X2=4.89 $Y2=4.24
r43 7 15 36.4 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=5
+ $X=3.13 $Y=3.985 $X2=3.335 $Y2=4.07
r44 7 11 36.4 $w=1.7e-07 $l=1.802e-06 $layer=licon1_NTAP_notbjt $count=5 $X=3.13
+ $Y=3.985 $X2=4.89 $Y2=4.07
r45 1 25 300 $w=1.7e-07 $l=1.4433e-06 $layer=licon1_PDIFF $count=2 $X=3.915
+ $Y=2.215 $X2=4.055 $Y2=3.59
r46 1 19 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=3.915
+ $Y=2.215 $X2=4.055 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%A_662_81# 1 2 9 12 16 17 19 20
+ 23 27 29 31
r47 25 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=1.285
+ $X2=4.99 $Y2=1.2
r48 25 27 48.6331 $w=2.48e-07 $l=1.055e-06 $layer=LI1_cond $X=4.99 $Y=1.285
+ $X2=4.99 $Y2=2.34
r49 21 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=1.115
+ $X2=4.99 $Y2=1.2
r50 21 23 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=4.99 $Y=1.115
+ $X2=4.99 $Y2=0.745
r51 19 29 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.865 $Y=1.2
+ $X2=4.99 $Y2=1.2
r52 19 20 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=4.865 $Y=1.2
+ $X2=3.895 $Y2=1.2
r53 17 32 29.6268 $w=6.05e-07 $l=3.15e-07 $layer=POLY_cond $X=3.612 $Y=1.58
+ $X2=3.612 $Y2=1.895
r54 17 31 18.1303 $w=6.05e-07 $l=1.85e-07 $layer=POLY_cond $X=3.612 $Y=1.58
+ $X2=3.612 $Y2=1.395
r55 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.58 $X2=3.73 $Y2=1.58
r56 14 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.73 $Y=1.285
+ $X2=3.895 $Y2=1.2
r57 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.73 $Y=1.285
+ $X2=3.73 $Y2=1.58
r58 12 32 114.496 $w=5e-07 $l=1.07e-06 $layer=POLY_cond $X=3.665 $Y=2.965
+ $X2=3.665 $Y2=1.895
r59 9 31 46.754 $w=5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.56 $Y=0.91 $X2=3.56
+ $Y2=1.395
r60 2 27 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.81
+ $Y=2.215 $X2=4.95 $Y2=2.34
r61 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.81
+ $Y=0.535 $X2=4.95 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%A 1 2 3 4 5 12 16 18
r23 15 18 111.286 $w=5e-07 $l=1.04e-06 $layer=POLY_cond $X=4.56 $Y=1.55 $X2=4.56
+ $Y2=2.59
r24 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.52
+ $Y=1.55 $X2=4.52 $Y2=1.55
r25 12 15 86.1397 $w=5e-07 $l=8.05e-07 $layer=POLY_cond $X=4.56 $Y=0.745
+ $X2=4.56 $Y2=1.55
r26 4 5 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=2.775 $X2=4.52
+ $Y2=3.145
r27 3 4 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=2.405 $X2=4.52
+ $Y2=2.775
r28 2 3 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=2.035 $X2=4.52
+ $Y2=2.405
r29 1 2 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.52 $Y=1.665 $X2=4.52
+ $Y2=2.035
r30 1 16 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.52 $Y=1.665
+ $X2=4.52 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%X 1 2 7 8 9 10 11 12 13 24 36
+ 46
r19 46 47 6.24827 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.217 $Y=2.34
+ $X2=3.217 $Y2=2.175
r20 34 36 0.207181 $w=4.43e-07 $l=8e-09 $layer=LI1_cond $X=3.217 $Y=2.397
+ $X2=3.217 $Y2=2.405
r21 13 43 11.5244 $w=4.43e-07 $l=4.45e-07 $layer=LI1_cond $X=3.217 $Y=3.145
+ $X2=3.217 $Y2=3.59
r22 12 13 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.217 $Y=2.775
+ $X2=3.217 $Y2=3.145
r23 11 34 1.01001 $w=4.43e-07 $l=3.9e-08 $layer=LI1_cond $X=3.217 $Y=2.358
+ $X2=3.217 $Y2=2.397
r24 11 46 0.466157 $w=4.43e-07 $l=1.8e-08 $layer=LI1_cond $X=3.217 $Y=2.358
+ $X2=3.217 $Y2=2.34
r25 11 12 8.598 $w=4.43e-07 $l=3.32e-07 $layer=LI1_cond $X=3.217 $Y=2.443
+ $X2=3.217 $Y2=2.775
r26 11 36 0.984109 $w=4.43e-07 $l=3.8e-08 $layer=LI1_cond $X=3.217 $Y=2.443
+ $X2=3.217 $Y2=2.405
r27 10 47 6.20546 $w=2.58e-07 $l=1.4e-07 $layer=LI1_cond $X=3.125 $Y=2.035
+ $X2=3.125 $Y2=2.175
r28 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.125 $Y=1.665
+ $X2=3.125 $Y2=2.035
r29 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.125 $Y=1.295
+ $X2=3.125 $Y2=1.665
r30 7 8 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.125 $Y=0.925
+ $X2=3.125 $Y2=1.295
r31 7 24 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=3.125 $Y=0.925
+ $X2=3.125 $Y2=0.68
r32 2 46 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.215 $X2=3.275 $Y2=2.34
r33 2 43 300 $w=1.7e-07 $l=1.44568e-06 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=2.215 $X2=3.275 $Y2=3.59
r34 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=3.045
+ $Y=0.535 $X2=3.17 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HVL__LSBUFHV2LV_SIMPLE_1%VGND 1 4 5 9 13
r23 9 15 2.684 $w=1.248e-06 $l=2.75e-07 $layer=LI1_cond $X=4.06 $Y=0.48 $X2=4.06
+ $Y2=0.755
r24 9 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.6 $Y=0.48 $X2=4.6
+ $Y2=0.48
r25 9 10 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.52 $Y=0.48
+ $X2=3.52 $Y2=0.48
r26 4 13 0.107494 $w=3.7e-07 $l=2.8e-07 $layer=MET1_cond $X=4.32 $Y=0.44 $X2=4.6
+ $Y2=0.44
r27 4 10 0.307124 $w=3.7e-07 $l=8e-07 $layer=MET1_cond $X=4.32 $Y=0.44 $X2=3.52
+ $Y2=0.44
r28 1 15 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=3.81
+ $Y=0.535 $X2=3.95 $Y2=0.755
.ends

