* File: sky130_fd_sc_hvl__sdfsbp_1.spice
* Created: Wed Sep  2 09:10:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hvl__sdfsbp_1.pex.spice"
.subckt sky130_fd_sc_hvl__sdfsbp_1  VNB VPB SCE D SCD CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_SCE_M1014_g N_A_30_569#_M1014_s N_VNB_M1014_b NHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250004 A=0.21 P=1.84 MULT=1
MM1029 A_348_107# N_D_M1029_g N_VGND_M1014_d N_VNB_M1014_b NHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84 SA=250001
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1028 N_A_485_569#_M1028_d N_A_30_569#_M1028_g A_348_107# N_VNB_M1014_b NHV
+ L=0.5 W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1016 A_646_107# N_SCE_M1016_g N_A_485_569#_M1028_d N_VNB_M1014_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1017 N_VGND_M1017_d N_SCD_M1017_g A_646_107# N_VNB_M1014_b NHV L=0.5 W=0.42
+ AD=0.09345 AS=0.0441 PD=0.865 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250003
+ SB=250001 A=0.21 P=1.84 MULT=1
MM1001 N_A_972_569#_M1001_d N_CLK_M1001_g N_VGND_M1017_d N_VNB_M1014_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.09345 PD=1.37 PS=0.865 NRD=0 NRS=44.7792 M=1 R=0.84
+ SA=250004 SB=250000 A=0.21 P=1.84 MULT=1
MM1022 N_A_1243_116#_M1022_d N_A_972_569#_M1022_g N_VGND_M1022_s N_VNB_M1014_b
+ NHV L=0.5 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=0.84
+ SA=250000 SB=250000 A=0.21 P=1.84 MULT=1
MM1007 N_A_1513_120#_M1007_d N_A_972_569#_M1007_g N_A_485_569#_M1007_s
+ N_VNB_M1014_b NHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250002 A=0.21 P=1.84 MULT=1
MM1023 A_1669_120# N_A_1243_116#_M1023_g N_A_1513_120#_M1007_d N_VNB_M1014_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250001 SB=250001 A=0.21 P=1.84 MULT=1
MM1040 N_VGND_M1040_d N_A_1711_94#_M1040_g A_1669_120# N_VNB_M1014_b NHV L=0.5
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84
+ SA=250002 SB=250000 A=0.21 P=1.84 MULT=1
MM1033 A_2077_107# N_A_1513_120#_M1033_g N_A_1711_94#_M1033_s N_VNB_M1014_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=13.566 NRS=0 M=1 R=0.84
+ SA=250000 SB=250003 A=0.21 P=1.84 MULT=1
MM1038 N_VGND_M1038_d N_SET_B_M1038_g A_2077_107# N_VNB_M1014_b NHV L=0.5 W=0.42
+ AD=0.0879308 AS=0.0441 PD=0.807692 PS=0.63 NRD=25.7754 NRS=13.566 M=1 R=0.84
+ SA=250001 SB=250002 A=0.21 P=1.84 MULT=1
MM1024 A_2394_107# N_A_1513_120#_M1024_g N_VGND_M1038_d N_VNB_M1014_b NHV L=0.5
+ W=0.75 AD=0.07875 AS=0.157019 PD=0.96 PS=1.44231 NRD=7.5924 NRS=0 M=1 R=1.5
+ SA=250001 SB=250002 A=0.375 P=2.5 MULT=1
MM1041 N_A_2501_543#_M1041_d N_A_1243_116#_M1041_g A_2394_107# N_VNB_M1014_b NHV
+ L=0.5 W=0.75 AD=0.166635 AS=0.07875 PD=1.46795 PS=0.96 NRD=0 NRS=7.5924 M=1
+ R=1.5 SA=250002 SB=250001 A=0.375 P=2.5 MULT=1
MM1008 A_2715_173# N_A_972_569#_M1008_g N_A_2501_543#_M1041_d N_VNB_M1014_b NHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0933154 PD=0.63 PS=0.822051 NRD=13.566 NRS=31.2132
+ M=1 R=0.84 SA=250002 SB=250001 A=0.21 P=1.84 MULT=1
MM1009 A_2857_173# N_A_2729_463#_M1009_g A_2715_173# N_VNB_M1014_b NHV L=0.5
+ W=0.42 AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=13.566 NRS=13.566 M=1 R=0.84
+ SA=250003 SB=250001 A=0.21 P=1.84 MULT=1
MM1010 N_VGND_M1010_d N_SET_B_M1010_g A_2857_173# N_VNB_M1014_b NHV L=0.5 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=13.566 M=1 R=0.84 SA=250003
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1027 N_VGND_M1027_d N_A_2501_543#_M1027_g N_A_2729_463#_M1027_s N_VNB_M1014_b
+ NHV L=0.5 W=0.42 AD=0.0933154 AS=0.1197 PD=0.822051 PS=1.41 NRD=31.2132 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1026 N_Q_N_M1026_d N_A_2501_543#_M1026_g N_VGND_M1027_d N_VNB_M1014_b NHV
+ L=0.5 W=0.75 AD=0.21375 AS=0.166635 PD=2.07 PS=1.46795 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1034 N_VGND_M1034_d N_A_2501_543#_M1034_g N_A_3609_173#_M1034_s N_VNB_M1014_b
+ NHV L=0.5 W=0.42 AD=0.0933154 AS=0.1197 PD=0.822051 PS=1.41 NRD=31.2132 NRS=0
+ M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1003 N_Q_M1003_d N_A_3609_173#_M1003_g N_VGND_M1034_d N_VNB_M1014_b NHV L=0.5
+ W=0.75 AD=0.21375 AS=0.166635 PD=2.07 PS=1.46795 NRD=0 NRS=0 M=1 R=1.5
+ SA=250001 SB=250000 A=0.375 P=2.5 MULT=1
MM1000 N_VPWR_M1000_d N_SCE_M1000_g N_A_30_569#_M1000_s N_VPB_M1000_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250004 A=0.21 P=1.84 MULT=1
MM1012 A_343_569# N_SCE_M1012_g N_VPWR_M1000_d N_VPB_M1000_b PHV L=0.5 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84 SA=250001
+ SB=250003 A=0.21 P=1.84 MULT=1
MM1015 N_A_485_569#_M1015_d N_D_M1015_g A_343_569# N_VPB_M1000_b PHV L=0.5
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1005 A_641_569# N_A_30_569#_M1005_g N_A_485_569#_M1015_d N_VPB_M1000_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250002 SB=250002 A=0.21 P=1.84 MULT=1
MM1006 N_VPWR_M1006_d N_SCD_M1006_g A_641_569# N_VPB_M1000_b PHV L=0.5 W=0.42
+ AD=0.100854 AS=0.0441 PD=0.857949 PS=0.63 NRD=75.0248 NRS=22.729 M=1 R=0.84
+ SA=250003 SB=250001 A=0.21 P=1.84 MULT=1
MM1025 N_A_972_569#_M1025_d N_CLK_M1025_g N_VPWR_M1006_d N_VPB_M1000_b PHV L=0.5
+ W=0.75 AD=0.21375 AS=0.180096 PD=2.07 PS=1.53205 NRD=0 NRS=0 M=1 R=1.5
+ SA=250002 SB=250000 A=0.375 P=2.5 MULT=1
MM1011 N_A_1243_116#_M1011_d N_A_972_569#_M1011_g N_VPWR_M1011_s N_VPB_M1000_b
+ PHV L=0.5 W=0.75 AD=0.19875 AS=0.21375 PD=2.03 PS=2.07 NRD=0 NRS=0 M=1 R=1.5
+ SA=250000 SB=250000 A=0.375 P=2.5 MULT=1
MM1004 N_A_1513_120#_M1004_d N_A_1243_116#_M1004_g N_A_485_569#_M1004_s
+ N_VPB_M1000_b PHV L=0.5 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0
+ M=1 R=0.84 SA=250000 SB=250007 A=0.21 P=1.84 MULT=1
MM1030 A_1710_556# N_A_972_569#_M1030_g N_A_1513_120#_M1004_d N_VPB_M1000_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=22.729 NRS=0 M=1 R=0.84
+ SA=250001 SB=250006 A=0.21 P=1.84 MULT=1
MM1035 N_VPWR_M1035_d N_A_1711_94#_M1035_g A_1710_556# N_VPB_M1000_b PHV L=0.5
+ W=0.42 AD=0.0756 AS=0.0441 PD=0.78 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1013 N_A_1711_94#_M1013_d N_A_1513_120#_M1013_g N_VPWR_M1035_d N_VPB_M1000_b
+ PHV L=0.5 W=0.42 AD=0.0588 AS=0.0756 PD=0.7 PS=0.78 NRD=0 NRS=36.3664 M=1
+ R=0.84 SA=250002 SB=250005 A=0.21 P=1.84 MULT=1
MM1018 N_VPWR_M1018_d N_SET_B_M1018_g N_A_1711_94#_M1013_d N_VPB_M1000_b PHV
+ L=0.5 W=0.42 AD=0.0979606 AS=0.0588 PD=0.825211 PS=0.7 NRD=81.0413 NRS=0 M=1
+ R=0.84 SA=250003 SB=250004 A=0.21 P=1.84 MULT=1
MM1021 A_2359_543# N_A_1513_120#_M1021_g N_VPWR_M1018_d N_VPB_M1000_b PHV L=0.5
+ W=1 AD=0.105 AS=0.233239 PD=1.21 PS=1.96479 NRD=9.5309 NRS=0 M=1 R=2 SA=250002
+ SB=250002 A=0.5 P=3 MULT=1
MM1037 N_A_2501_543#_M1037_d N_A_972_569#_M1037_g A_2359_543# N_VPB_M1000_b PHV
+ L=0.5 W=1 AD=0.257887 AS=0.105 PD=2.01408 PS=1.21 NRD=6.6659 NRS=9.5309 M=1
+ R=2 SA=250002 SB=250001 A=0.5 P=3 MULT=1
MM1020 A_2687_543# N_A_1243_116#_M1020_g N_A_2501_543#_M1037_d N_VPB_M1000_b PHV
+ L=0.5 W=0.42 AD=0.0441 AS=0.108313 PD=0.63 PS=0.845915 NRD=22.729 NRS=52.2958
+ M=1 R=0.84 SA=250005 SB=250002 A=0.21 P=1.84 MULT=1
MM1039 N_VPWR_M1039_d N_A_2729_463#_M1039_g A_2687_543# N_VPB_M1000_b PHV L=0.5
+ W=0.42 AD=0.0735 AS=0.0441 PD=0.77 PS=0.63 NRD=0 NRS=22.729 M=1 R=0.84
+ SA=250006 SB=250001 A=0.21 P=1.84 MULT=1
MM1031 N_A_2501_543#_M1031_d N_SET_B_M1031_g N_VPWR_M1039_d N_VPB_M1000_b PHV
+ L=0.5 W=0.42 AD=0.1197 AS=0.0735 PD=1.41 PS=0.77 NRD=0 NRS=31.8206 M=1 R=0.84
+ SA=250007 SB=250000 A=0.21 P=1.84 MULT=1
MM1002 N_VPWR_M1002_d N_A_2501_543#_M1002_g N_A_2729_463#_M1002_s N_VPB_M1000_b
+ PHV L=0.5 W=0.42 AD=0.0970594 AS=0.168 PD=0.820312 PS=1.64 NRD=43.1851
+ NRS=52.2958 M=1 R=0.84 SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1036 N_Q_N_M1036_d N_A_2501_543#_M1036_g N_VPWR_M1002_d N_VPB_M1000_b PHV
+ L=0.5 W=1.5 AD=0.3975 AS=0.346641 PD=3.53 PS=2.92969 NRD=0 NRS=0 M=1 R=3
+ SA=250000 SB=250000 A=0.75 P=4 MULT=1
MM1032 N_VPWR_M1032_d N_A_2501_543#_M1032_g N_A_3609_173#_M1032_s N_VPB_M1000_b
+ PHV L=0.5 W=0.75 AD=0.1575 AS=0.21375 PD=1.19571 PS=2.07 NRD=29.2803 NRS=0 M=1
+ R=1.5 SA=250000 SB=250001 A=0.375 P=2.5 MULT=1
MM1019 N_Q_M1019_d N_A_3609_173#_M1019_g N_VPWR_M1032_d N_VPB_M1000_b PHV L=0.5
+ W=1 AD=0.285 AS=0.21 PD=2.57 PS=1.59429 NRD=0 NRS=0 M=1 R=2 SA=250001
+ SB=250000 A=0.5 P=3 MULT=1
DX42_noxref N_VNB_M1014_b N_VPB_M1000_b NWDIODE A=54.132 P=46.84
*
.include "sky130_fd_sc_hvl__sdfsbp_1.pxi.spice"
*
.ends
*
*
